module LDSTUnit(
  input  [4:0]  io_dinst_rd_bits,
  input  [4:0]  io_dinst_rs1,
  input  [4:0]  io_dinst_rs2,
  input  [25:0] io_dinst_imm,
  input         io_dinst_shift_val_valid,
  input  [5:0]  io_dinst_shift_val_bits,
  input  [4:0]  io_dinst_itype,
  input  [3:0]  io_dinst_op,
  input  [63:0] io_rVal1,
  input  [63:0] io_rVal2,
  output        io_minst_valid,
  output [1:0]  io_minst_bits_size,
  output        io_minst_bits_isPair,
  output        io_minst_bits_isLoad,
  output [63:0] io_minst_bits_memReq_0_addr,
  output [4:0]  io_minst_bits_memReq_0_reg,
  output [63:0] io_minst_bits_memReq_1_addr,
  output [4:0]  io_minst_bits_memReq_1_reg,
  output [63:0] io_minst_bits_rd_res,
  output        io_minst_bits_rd_valid,
  output [4:0]  io_minst_bits_rd_bits,
  output        io_minst_bits_unalignedExcpSP
);
  wire [63:0] extendReg_io_value; // @[LoadStore.scala 90:25]
  wire [2:0] extendReg_io_option; // @[LoadStore.scala 90:25]
  wire [1:0] extendReg_io_shift; // @[LoadStore.scala 90:25]
  wire [63:0] extendReg_io_res; // @[LoadStore.scala 90:25]
  wire [1:0] size; // @[LoadStore.scala 76:34]
  wire [6:0] _T_4; // @[LoadStore.scala 79:41]
  wire [63:0] offstSignExt7; // @[LoadStore.scala 79:56]
  wire [8:0] _T_7; // @[LoadStore.scala 80:41]
  wire [63:0] offstSignExt9; // @[LoadStore.scala 80:56]
  wire  _T_9; // @[LoadStore.scala 95:23]
  wire [14:0] _GEN_25; // @[LoadStore.scala 98:33]
  wire [14:0] _T_11; // @[LoadStore.scala 98:33]
  wire  _T_12; // @[LoadStore.scala 99:29]
  wire  _T_13; // @[LoadStore.scala 103:29]
  wire [66:0] _GEN_26; // @[LoadStore.scala 106:28]
  wire [66:0] _T_14; // @[LoadStore.scala 106:28]
  wire  _T_15; // @[LoadStore.scala 107:29]
  wire  _T_17; // @[LoadStore.scala 111:29]
  wire  _T_19; // @[LoadStore.scala 115:29]
  wire  _T_20; // @[LoadStore.scala 119:29]
  wire  _T_21; // @[LoadStore.scala 123:29]
  wire [63:0] _GEN_2; // @[LoadStore.scala 123:44]
  wire  _GEN_3; // @[LoadStore.scala 119:42]
  wire [63:0] _GEN_5; // @[LoadStore.scala 119:42]
  wire  _GEN_6; // @[LoadStore.scala 115:44]
  wire [63:0] _GEN_8; // @[LoadStore.scala 115:44]
  wire  _GEN_9; // @[LoadStore.scala 111:45]
  wire  _GEN_10; // @[LoadStore.scala 111:45]
  wire [66:0] _GEN_11; // @[LoadStore.scala 111:45]
  wire  _GEN_12; // @[LoadStore.scala 107:43]
  wire  _GEN_13; // @[LoadStore.scala 107:43]
  wire [66:0] _GEN_14; // @[LoadStore.scala 107:43]
  wire  _GEN_15; // @[LoadStore.scala 103:45]
  wire  _GEN_16; // @[LoadStore.scala 103:45]
  wire [66:0] _GEN_17; // @[LoadStore.scala 103:45]
  wire  _GEN_18; // @[LoadStore.scala 99:43]
  wire  _GEN_19; // @[LoadStore.scala 99:43]
  wire [66:0] _GEN_20; // @[LoadStore.scala 99:43]
  wire  postindex; // @[LoadStore.scala 95:37]
  wire [66:0] _GEN_23; // @[LoadStore.scala 95:37]
  wire  _T_22; // @[LoadStore.scala 133:21]
  wire [63:0] offst; // @[LoadStore.scala 98:11 LoadStore.scala 102:11 LoadStore.scala 106:11 LoadStore.scala 110:11 LoadStore.scala 114:11 LoadStore.scala 118:11 LoadStore.scala 122:11 LoadStore.scala 126:11]
  wire [63:0] _T_24; // @[LoadStore.scala 146:44]
  wire [63:0] ldst_address; // @[LoadStore.scala 147:19]
  wire  _T_31; // @[Mux.scala 80:60]
  wire  _T_33; // @[Mux.scala 80:60]
  wire  _T_34; // @[Mux.scala 80:57]
  wire  _T_35; // @[Mux.scala 80:60]
  wire  _T_36; // @[Mux.scala 80:57]
  wire  _T_37; // @[Mux.scala 80:60]
  wire  _T_38; // @[Mux.scala 80:57]
  wire  _T_39; // @[Mux.scala 80:60]
  wire  _T_40; // @[Mux.scala 80:57]
  wire  _T_41; // @[Mux.scala 80:60]
  wire  _T_42; // @[Mux.scala 80:57]
  wire  _T_43; // @[Mux.scala 80:60]
  wire  _T_44; // @[Mux.scala 80:57]
  wire  _T_45; // @[Mux.scala 80:60]
  wire [3:0] dbytes; // @[LoadStore.scala 195:20]
  wire  _T_49; // @[LoadStore.scala 197:34]
  wire [63:0] _GEN_29; // @[LoadStore.scala 200:48]
  wire  _T_58; // @[LoadStore.scala 215:77]
  ExtendReg extendReg ( // @[LoadStore.scala 90:25]
    .io_value(extendReg_io_value),
    .io_option(extendReg_io_option),
    .io_shift(extendReg_io_shift),
    .io_res(extendReg_io_res)
  );
  assign size = io_dinst_op[1:0]; // @[LoadStore.scala 76:34]
  assign _T_4 = io_dinst_imm[6:0]; // @[LoadStore.scala 79:41]
  assign offstSignExt7 = {{57{_T_4[6]}},_T_4}; // @[LoadStore.scala 79:56]
  assign _T_7 = io_dinst_imm[8:0]; // @[LoadStore.scala 80:41]
  assign offstSignExt9 = {{55{_T_7[8]}},_T_7}; // @[LoadStore.scala 80:56]
  assign _T_9 = io_dinst_itype == 5'h14; // @[LoadStore.scala 95:23]
  assign _GEN_25 = {{3'd0}, io_dinst_imm[11:0]}; // @[LoadStore.scala 98:33]
  assign _T_11 = _GEN_25 << size; // @[LoadStore.scala 98:33]
  assign _T_12 = io_dinst_itype == 5'h10; // @[LoadStore.scala 99:29]
  assign _T_13 = io_dinst_itype == 5'h15; // @[LoadStore.scala 103:29]
  assign _GEN_26 = {{3'd0}, offstSignExt7}; // @[LoadStore.scala 106:28]
  assign _T_14 = _GEN_26 << size; // @[LoadStore.scala 106:28]
  assign _T_15 = io_dinst_itype == 5'h16; // @[LoadStore.scala 107:29]
  assign _T_17 = io_dinst_itype == 5'h17; // @[LoadStore.scala 111:29]
  assign _T_19 = io_dinst_itype == 5'h11; // @[LoadStore.scala 115:29]
  assign _T_20 = io_dinst_itype == 5'h12; // @[LoadStore.scala 119:29]
  assign _T_21 = io_dinst_itype == 5'h13; // @[LoadStore.scala 123:29]
  assign _GEN_2 = _T_21 ? offstSignExt9 : {{38'd0}, io_dinst_imm}; // @[LoadStore.scala 123:44]
  assign _GEN_3 = _T_20 ? 1'h0 : _T_21; // @[LoadStore.scala 119:42]
  assign _GEN_5 = _T_20 ? extendReg_io_res : _GEN_2; // @[LoadStore.scala 119:42]
  assign _GEN_6 = _T_19 | _GEN_3; // @[LoadStore.scala 115:44]
  assign _GEN_8 = _T_19 ? offstSignExt9 : _GEN_5; // @[LoadStore.scala 115:44]
  assign _GEN_9 = _T_17 | _GEN_6; // @[LoadStore.scala 111:45]
  assign _GEN_10 = _T_17 ? 1'h0 : _T_19; // @[LoadStore.scala 111:45]
  assign _GEN_11 = _T_17 ? _T_14 : {{3'd0}, _GEN_8}; // @[LoadStore.scala 111:45]
  assign _GEN_12 = _T_15 ? 1'h0 : _GEN_9; // @[LoadStore.scala 107:43]
  assign _GEN_13 = _T_15 ? 1'h0 : _GEN_10; // @[LoadStore.scala 107:43]
  assign _GEN_14 = _T_15 ? _T_14 : _GEN_11; // @[LoadStore.scala 107:43]
  assign _GEN_15 = _T_13 | _GEN_12; // @[LoadStore.scala 103:45]
  assign _GEN_16 = _T_13 | _GEN_13; // @[LoadStore.scala 103:45]
  assign _GEN_17 = _T_13 ? _T_14 : _GEN_14; // @[LoadStore.scala 103:45]
  assign _GEN_18 = _T_12 ? 1'h0 : _GEN_15; // @[LoadStore.scala 99:43]
  assign _GEN_19 = _T_12 ? 1'h0 : _GEN_16; // @[LoadStore.scala 99:43]
  assign _GEN_20 = _T_12 ? {{3'd0}, offstSignExt9} : _GEN_17; // @[LoadStore.scala 99:43]
  assign postindex = _T_9 ? 1'h0 : _GEN_19; // @[LoadStore.scala 95:37]
  assign _GEN_23 = _T_9 ? {{52'd0}, _T_11} : _GEN_20; // @[LoadStore.scala 95:37]
  assign _T_22 = io_dinst_rs1 == 5'h1f; // @[LoadStore.scala 133:21]
  assign offst = _GEN_23[63:0]; // @[LoadStore.scala 98:11 LoadStore.scala 102:11 LoadStore.scala 106:11 LoadStore.scala 110:11 LoadStore.scala 114:11 LoadStore.scala 118:11 LoadStore.scala 122:11 LoadStore.scala 126:11]
  assign _T_24 = io_rVal1 + offst; // @[LoadStore.scala 146:44]
  assign ldst_address = postindex ? io_rVal1 : _T_24; // @[LoadStore.scala 147:19]
  assign _T_31 = 5'h17 == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_33 = 5'h16 == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_34 = _T_33 | _T_31; // @[Mux.scala 80:57]
  assign _T_35 = 5'h15 == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_36 = _T_35 | _T_34; // @[Mux.scala 80:57]
  assign _T_37 = 5'h10 == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_38 = _T_37 | _T_36; // @[Mux.scala 80:57]
  assign _T_39 = 5'h13 == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_40 = _T_39 | _T_38; // @[Mux.scala 80:57]
  assign _T_41 = 5'h12 == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_42 = _T_41 | _T_40; // @[Mux.scala 80:57]
  assign _T_43 = 5'h11 == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_44 = _T_43 | _T_42; // @[Mux.scala 80:57]
  assign _T_45 = 5'h14 == io_dinst_itype; // @[Mux.scala 80:60]
  assign dbytes = 4'h1 << size; // @[LoadStore.scala 195:20]
  assign _T_49 = _T_17 | _T_15; // @[LoadStore.scala 197:34]
  assign _GEN_29 = {{60'd0}, dbytes}; // @[LoadStore.scala 200:48]
  assign _T_58 = _T_24[1:0] != 2'h0; // @[LoadStore.scala 215:77]
  assign io_minst_valid = _T_45 | _T_44; // @[LoadStore.scala 180:18]
  assign io_minst_bits_size = io_dinst_op[1:0]; // @[LoadStore.scala 176:22]
  assign io_minst_bits_isPair = _T_49 | _T_13; // @[LoadStore.scala 196:24]
  assign io_minst_bits_isLoad = io_dinst_op[2]; // @[LoadStore.scala 179:24]
  assign io_minst_bits_memReq_0_addr = postindex ? io_rVal1 : _T_24; // @[LoadStore.scala 191:32]
  assign io_minst_bits_memReq_0_reg = io_dinst_rd_bits; // @[LoadStore.scala 193:31]
  assign io_minst_bits_memReq_1_addr = ldst_address + _GEN_29; // @[LoadStore.scala 200:32]
  assign io_minst_bits_memReq_1_reg = io_dinst_rs2; // @[LoadStore.scala 202:31]
  assign io_minst_bits_rd_res = io_rVal1 + offst; // @[LoadStore.scala 216:24]
  assign io_minst_bits_rd_valid = _T_9 ? 1'h0 : _GEN_18; // @[LoadStore.scala 218:26]
  assign io_minst_bits_rd_bits = io_dinst_rs1; // @[LoadStore.scala 217:25]
  assign io_minst_bits_unalignedExcpSP = _T_22 & _T_58; // @[LoadStore.scala 215:33]
  assign extendReg_io_value = io_rVal2; // @[LoadStore.scala 91:22]
  assign extendReg_io_option = io_dinst_shift_val_bits[2:0]; // @[LoadStore.scala 92:23]
  assign extendReg_io_shift = io_dinst_shift_val_valid ? size : 2'h0; // @[LoadStore.scala 93:22]
endmodule
