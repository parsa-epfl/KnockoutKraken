module BranchUnit( // @[:@2674.2]
  input  [25:0] io_dinst_imm_bits, // @[:@2677.4]
  input  [3:0]  io_dinst_cond_bits, // @[:@2677.4]
  input  [2:0]  io_dinst_itype, // @[:@2677.4]
  input  [2:0]  io_dinst_op, // @[:@2677.4]
  input         io_dinst_tag, // @[:@2677.4]
  input  [3:0]  io_nzcv, // @[:@2677.4]
  output        io_binst_valid, // @[:@2677.4]
  output [63:0] io_binst_bits_offset, // @[:@2677.4]
  output        io_binst_bits_tag // @[:@2677.4]
);
  wire [3:0] cond_io_cond; // @[branch.scala 61:20:@2686.4]
  wire [3:0] cond_io_nzcv; // @[branch.scala 61:20:@2686.4]
  wire  cond_io_res; // @[branch.scala 61:20:@2686.4]
  wire [25:0] _T_99; // @[branch.scala 57:37:@2682.4]
  wire [63:0] signExtended; // @[branch.scala 56:26:@2681.4 branch.scala 57:16:@2683.4]
  wire  _T_101; // @[branch.scala 64:24:@2691.4]
  wire  _T_102; // @[branch.scala 64:54:@2692.4]
  wire  _T_103; // @[branch.scala 64:36:@2693.4]
  wire  _T_104; // @[branch.scala 65:22:@2695.6]
  wire  _T_105; // @[branch.scala 67:28:@2700.8]
  wire  _GEN_1; // @[branch.scala 65:36:@2696.6]
  CondUnit cond ( // @[branch.scala 61:20:@2686.4]
    .io_cond(cond_io_cond),
    .io_nzcv(cond_io_nzcv),
    .io_res(cond_io_res)
  );
  assign _T_99 = $signed(io_dinst_imm_bits); // @[branch.scala 57:37:@2682.4]
  assign signExtended = {{38{_T_99[25]}},_T_99}; // @[branch.scala 56:26:@2681.4 branch.scala 57:16:@2683.4]
  assign _T_101 = io_dinst_itype == 3'h2; // @[branch.scala 64:24:@2691.4]
  assign _T_102 = io_dinst_itype == 3'h3; // @[branch.scala 64:54:@2692.4]
  assign _T_103 = _T_101 | _T_102; // @[branch.scala 64:36:@2693.4]
  assign _T_104 = io_dinst_op == 3'h1; // @[branch.scala 65:22:@2695.6]
  assign _T_105 = io_dinst_op == 3'h0; // @[branch.scala 67:28:@2700.8]
  assign _GEN_1 = _T_104 ? cond_io_res : _T_105; // @[branch.scala 65:36:@2696.6]
  assign io_binst_valid = _T_103 ? _GEN_1 : 1'h0; // @[branch.scala 52:18:@2679.4 branch.scala 66:22:@2697.8 branch.scala 68:22:@2702.10]
  assign io_binst_bits_offset = $unsigned(signExtended); // @[branch.scala 58:24:@2685.4]
  assign io_binst_bits_tag = io_dinst_tag; // @[branch.scala 53:21:@2680.4]
  assign cond_io_cond = io_dinst_cond_bits; // @[branch.scala 62:16:@2689.4]
  assign cond_io_nzcv = io_nzcv; // @[branch.scala 63:16:@2690.4]
endmodule
