module BasicALU( // @[:@2440.2]
  input  [63:0] io_a, // @[:@2443.4]
  input  [63:0] io_b, // @[:@2443.4]
  input  [2:0]  io_opcode, // @[:@2443.4]
  output [63:0] io_res, // @[:@2443.4]
  output [3:0]  io_nzcv // @[:@2443.4]
);
  wire [63:0] _T_16; // @[execute.scala 30:34:@2445.4]
  wire [63:0] _T_17; // @[execute.scala 31:36:@2446.4]
  wire [63:0] _T_18; // @[execute.scala 31:34:@2447.4]
  wire [63:0] _T_19; // @[execute.scala 32:34:@2448.4]
  wire [63:0] _T_21; // @[execute.scala 33:34:@2450.4]
  wire [63:0] _T_22; // @[execute.scala 34:34:@2451.4]
  wire [63:0] _T_24; // @[execute.scala 35:34:@2453.4]
  wire [64:0] _T_25; // @[execute.scala 36:34:@2454.4]
  wire [63:0] _T_26; // @[execute.scala 36:34:@2455.4]
  wire [64:0] _T_27; // @[execute.scala 37:34:@2456.4]
  wire [64:0] _T_28; // @[execute.scala 37:34:@2457.4]
  wire [63:0] _T_29; // @[execute.scala 37:34:@2458.4]
  wire  _T_30; // @[Mux.scala 46:19:@2459.4]
  wire [63:0] _T_31; // @[Mux.scala 46:16:@2460.4]
  wire  _T_32; // @[Mux.scala 46:19:@2461.4]
  wire [63:0] _T_33; // @[Mux.scala 46:16:@2462.4]
  wire  _T_34; // @[Mux.scala 46:19:@2463.4]
  wire [63:0] _T_35; // @[Mux.scala 46:16:@2464.4]
  wire  _T_36; // @[Mux.scala 46:19:@2465.4]
  wire [63:0] _T_37; // @[Mux.scala 46:16:@2466.4]
  wire  _T_38; // @[Mux.scala 46:19:@2467.4]
  wire [63:0] _T_39; // @[Mux.scala 46:16:@2468.4]
  wire  _T_40; // @[Mux.scala 46:19:@2469.4]
  wire [63:0] _T_41; // @[Mux.scala 46:16:@2470.4]
  wire  _T_42; // @[Mux.scala 46:19:@2471.4]
  wire [63:0] _T_43; // @[Mux.scala 46:16:@2472.4]
  wire  _T_44; // @[Mux.scala 46:19:@2473.4]
  wire [63:0] res; // @[Mux.scala 46:16:@2474.4]
  wire [63:0] _T_58; // @[execute.scala 44:18:@2480.4]
  wire  nzcv_0; // @[execute.scala 44:25:@2481.4]
  wire  nzcv_1; // @[execute.scala 45:18:@2483.4]
  wire  nzcv_2; // @[execute.scala 47:28:@2486.4]
  wire [63:0] _T_67; // @[execute.scala 49:23:@2489.4]
  wire [63:0] _T_68; // @[execute.scala 49:37:@2490.4]
  wire [64:0] _T_69; // @[execute.scala 49:30:@2491.4]
  wire [63:0] _T_70; // @[execute.scala 49:30:@2492.4]
  wire [63:0] sign_sum; // @[execute.scala 49:30:@2493.4]
  wire  _T_73; // @[execute.scala 50:27:@2495.4]
  wire  _T_76; // @[execute.scala 50:47:@2497.4]
  wire  isPos; // @[execute.scala 50:33:@2498.4]
  wire  _T_79; // @[execute.scala 51:27:@2500.4]
  wire  _T_82; // @[execute.scala 51:47:@2502.4]
  wire  isNeg; // @[execute.scala 51:33:@2503.4]
  wire  _T_84; // @[execute.scala 53:27:@2505.6]
  wire  _T_86; // @[execute.scala 53:16:@2506.6]
  wire  _T_88; // @[execute.scala 55:27:@2511.8]
  wire  _T_90; // @[execute.scala 55:16:@2512.8]
  wire  _GEN_0; // @[execute.scala 54:21:@2510.6]
  wire  nzcv_3; // @[execute.scala 52:15:@2504.4]
  wire [1:0] _T_92; // @[execute.scala 60:19:@2518.4]
  wire [1:0] _T_93; // @[execute.scala 60:19:@2519.4]
  assign _T_16 = io_a & io_b; // @[execute.scala 30:34:@2445.4]
  assign _T_17 = ~ io_b; // @[execute.scala 31:36:@2446.4]
  assign _T_18 = io_a & _T_17; // @[execute.scala 31:34:@2447.4]
  assign _T_19 = io_a | io_b; // @[execute.scala 32:34:@2448.4]
  assign _T_21 = io_a | _T_17; // @[execute.scala 33:34:@2450.4]
  assign _T_22 = io_a ^ io_b; // @[execute.scala 34:34:@2451.4]
  assign _T_24 = io_a ^ _T_17; // @[execute.scala 35:34:@2453.4]
  assign _T_25 = io_a + io_b; // @[execute.scala 36:34:@2454.4]
  assign _T_26 = io_a + io_b; // @[execute.scala 36:34:@2455.4]
  assign _T_27 = io_a - io_b; // @[execute.scala 37:34:@2456.4]
  assign _T_28 = $unsigned(_T_27); // @[execute.scala 37:34:@2457.4]
  assign _T_29 = _T_28[63:0]; // @[execute.scala 37:34:@2458.4]
  assign _T_30 = 3'h7 == io_opcode; // @[Mux.scala 46:19:@2459.4]
  assign _T_31 = _T_30 ? _T_29 : 64'h0; // @[Mux.scala 46:16:@2460.4]
  assign _T_32 = 3'h6 == io_opcode; // @[Mux.scala 46:19:@2461.4]
  assign _T_33 = _T_32 ? _T_26 : _T_31; // @[Mux.scala 46:16:@2462.4]
  assign _T_34 = 3'h5 == io_opcode; // @[Mux.scala 46:19:@2463.4]
  assign _T_35 = _T_34 ? _T_24 : _T_33; // @[Mux.scala 46:16:@2464.4]
  assign _T_36 = 3'h4 == io_opcode; // @[Mux.scala 46:19:@2465.4]
  assign _T_37 = _T_36 ? _T_22 : _T_35; // @[Mux.scala 46:16:@2466.4]
  assign _T_38 = 3'h3 == io_opcode; // @[Mux.scala 46:19:@2467.4]
  assign _T_39 = _T_38 ? _T_21 : _T_37; // @[Mux.scala 46:16:@2468.4]
  assign _T_40 = 3'h2 == io_opcode; // @[Mux.scala 46:19:@2469.4]
  assign _T_41 = _T_40 ? _T_19 : _T_39; // @[Mux.scala 46:16:@2470.4]
  assign _T_42 = 3'h1 == io_opcode; // @[Mux.scala 46:19:@2471.4]
  assign _T_43 = _T_42 ? _T_18 : _T_41; // @[Mux.scala 46:16:@2472.4]
  assign _T_44 = 3'h0 == io_opcode; // @[Mux.scala 46:19:@2473.4]
  assign res = _T_44 ? _T_16 : _T_43; // @[Mux.scala 46:16:@2474.4]
  assign _T_58 = $signed(res); // @[execute.scala 44:18:@2480.4]
  assign nzcv_0 = $signed(_T_58) < $signed(64'sh0); // @[execute.scala 44:25:@2481.4]
  assign nzcv_1 = res == 64'h0; // @[execute.scala 45:18:@2483.4]
  assign nzcv_2 = _T_25[64]; // @[execute.scala 47:28:@2486.4]
  assign _T_67 = $signed(io_a); // @[execute.scala 49:23:@2489.4]
  assign _T_68 = $signed(io_b); // @[execute.scala 49:37:@2490.4]
  assign _T_69 = $signed(_T_67) + $signed(_T_68); // @[execute.scala 49:30:@2491.4]
  assign _T_70 = $signed(_T_67) + $signed(_T_68); // @[execute.scala 49:30:@2492.4]
  assign sign_sum = $signed(_T_70); // @[execute.scala 49:30:@2493.4]
  assign _T_73 = $signed(_T_67) > $signed(64'sh0); // @[execute.scala 50:27:@2495.4]
  assign _T_76 = $signed(_T_68) > $signed(64'sh0); // @[execute.scala 50:47:@2497.4]
  assign isPos = _T_73 & _T_76; // @[execute.scala 50:33:@2498.4]
  assign _T_79 = $signed(_T_67) < $signed(64'sh0); // @[execute.scala 51:27:@2500.4]
  assign _T_82 = $signed(_T_68) < $signed(64'sh0); // @[execute.scala 51:47:@2502.4]
  assign isNeg = _T_79 & _T_82; // @[execute.scala 51:33:@2503.4]
  assign _T_84 = $signed(sign_sum) > $signed(64'sh0); // @[execute.scala 53:27:@2505.6]
  assign _T_86 = _T_84 == 1'h0; // @[execute.scala 53:16:@2506.6]
  assign _T_88 = $signed(sign_sum) < $signed(64'sh0); // @[execute.scala 55:27:@2511.8]
  assign _T_90 = _T_88 == 1'h0; // @[execute.scala 55:16:@2512.8]
  assign _GEN_0 = isNeg ? _T_90 : 1'h0; // @[execute.scala 54:21:@2510.6]
  assign nzcv_3 = isPos ? _T_86 : _GEN_0; // @[execute.scala 52:15:@2504.4]
  assign _T_92 = {nzcv_1,nzcv_0}; // @[execute.scala 60:19:@2518.4]
  assign _T_93 = {nzcv_3,nzcv_2}; // @[execute.scala 60:19:@2519.4]
  assign io_res = _T_44 ? _T_16 : _T_43; // @[execute.scala 62:10:@2522.4]
  assign io_nzcv = {_T_93,_T_92}; // @[execute.scala 60:11:@2521.4]
endmodule
