module DecodeBitMasks(
  input         io_immn,
  input  [5:0]  io_imms,
  input  [5:0]  io_immr,
  output [63:0] io_wmask,
  output [63:0] io_tmask,
  input         io_is32bit
);
  wire [5:0] _T; // @[Execute.scala 289:54]
  wire [6:0] toBeEncoded; // @[Cat.scala 29:58]
  wire [1:0] _T_10; // @[Mux.scala 47:69]
  wire [1:0] _T_11; // @[Mux.scala 47:69]
  wire [2:0] _T_12; // @[Mux.scala 47:69]
  wire [2:0] _T_13; // @[Mux.scala 47:69]
  wire [2:0] len; // @[Mux.scala 47:69]
  wire [6:0] _T_15;
  wire [63:0] _GEN_1; // @[Execute.scala 291:39]
  wire [63:0] _GEN_2; // @[Execute.scala 291:39]
  wire [63:0] _GEN_3; // @[Execute.scala 291:39]
  wire [63:0] _GEN_4; // @[Execute.scala 291:39]
  wire [63:0] _GEN_5; // @[Execute.scala 291:39]
  wire [63:0] _GEN_6; // @[Execute.scala 291:39]
  wire [63:0] _GEN_7; // @[Execute.scala 291:39]
  wire [63:0] _GEN_8; // @[Execute.scala 291:39]
  wire [63:0] _GEN_9; // @[Execute.scala 291:39]
  wire [63:0] _GEN_10; // @[Execute.scala 291:39]
  wire [63:0] _GEN_11; // @[Execute.scala 291:39]
  wire [63:0] _GEN_12; // @[Execute.scala 291:39]
  wire [63:0] _GEN_13; // @[Execute.scala 291:39]
  wire [63:0] _GEN_14; // @[Execute.scala 291:39]
  wire [63:0] _GEN_15; // @[Execute.scala 291:39]
  wire [63:0] _GEN_16; // @[Execute.scala 291:39]
  wire [63:0] _GEN_17; // @[Execute.scala 291:39]
  wire [63:0] _GEN_18; // @[Execute.scala 291:39]
  wire [63:0] _GEN_19; // @[Execute.scala 291:39]
  wire [63:0] _GEN_20; // @[Execute.scala 291:39]
  wire [63:0] _GEN_21; // @[Execute.scala 291:39]
  wire [63:0] _GEN_22; // @[Execute.scala 291:39]
  wire [63:0] _GEN_23; // @[Execute.scala 291:39]
  wire [63:0] _GEN_24; // @[Execute.scala 291:39]
  wire [63:0] _GEN_25; // @[Execute.scala 291:39]
  wire [63:0] _GEN_26; // @[Execute.scala 291:39]
  wire [63:0] _GEN_27; // @[Execute.scala 291:39]
  wire [63:0] _GEN_28; // @[Execute.scala 291:39]
  wire [63:0] _GEN_29; // @[Execute.scala 291:39]
  wire [63:0] _GEN_30; // @[Execute.scala 291:39]
  wire [63:0] _GEN_31; // @[Execute.scala 291:39]
  wire [63:0] _GEN_32; // @[Execute.scala 291:39]
  wire [63:0] _GEN_33; // @[Execute.scala 291:39]
  wire [63:0] _GEN_34; // @[Execute.scala 291:39]
  wire [63:0] _GEN_35; // @[Execute.scala 291:39]
  wire [63:0] _GEN_36; // @[Execute.scala 291:39]
  wire [63:0] _GEN_37; // @[Execute.scala 291:39]
  wire [63:0] _GEN_38; // @[Execute.scala 291:39]
  wire [63:0] _GEN_39; // @[Execute.scala 291:39]
  wire [63:0] _GEN_40; // @[Execute.scala 291:39]
  wire [63:0] _GEN_41; // @[Execute.scala 291:39]
  wire [63:0] _GEN_42; // @[Execute.scala 291:39]
  wire [63:0] _GEN_43; // @[Execute.scala 291:39]
  wire [63:0] _GEN_44; // @[Execute.scala 291:39]
  wire [63:0] _GEN_45; // @[Execute.scala 291:39]
  wire [63:0] _GEN_46; // @[Execute.scala 291:39]
  wire [63:0] _GEN_47; // @[Execute.scala 291:39]
  wire [63:0] _GEN_48; // @[Execute.scala 291:39]
  wire [63:0] _GEN_49; // @[Execute.scala 291:39]
  wire [63:0] _GEN_50; // @[Execute.scala 291:39]
  wire [63:0] _GEN_51; // @[Execute.scala 291:39]
  wire [63:0] _GEN_52; // @[Execute.scala 291:39]
  wire [63:0] _GEN_53; // @[Execute.scala 291:39]
  wire [63:0] _GEN_54; // @[Execute.scala 291:39]
  wire [63:0] _GEN_55; // @[Execute.scala 291:39]
  wire [63:0] _GEN_56; // @[Execute.scala 291:39]
  wire [63:0] _GEN_57; // @[Execute.scala 291:39]
  wire [63:0] _GEN_58; // @[Execute.scala 291:39]
  wire [63:0] _GEN_59; // @[Execute.scala 291:39]
  wire [63:0] _GEN_60; // @[Execute.scala 291:39]
  wire [63:0] _GEN_61; // @[Execute.scala 291:39]
  wire [63:0] _GEN_62; // @[Execute.scala 291:39]
  wire [63:0] _GEN_63; // @[Execute.scala 291:39]
  wire [63:0] _GEN_64; // @[Execute.scala 291:39]
  wire [5:0] levels; // @[Execute.scala 291:39]
  wire [5:0] s; // @[Execute.scala 293:28]
  wire [5:0] r; // @[Execute.scala 294:28]
  wire [6:0] diff; // @[Execute.scala 295:25]
  wire [6:0] _GEN_10436; // @[Execute.scala 297:25]
  wire [6:0] d; // @[Execute.scala 297:25]
  wire [6:0] onesS; // @[Execute.scala 298:26]
  wire [7:0] onesD; // @[Execute.scala 299:26]
  wire [63:0] _GEN_66; // @[Execute.scala 301:9]
  wire [63:0] _GEN_67; // @[Execute.scala 301:9]
  wire [63:0] _GEN_68; // @[Execute.scala 301:9]
  wire [63:0] _GEN_69; // @[Execute.scala 301:9]
  wire [63:0] _GEN_70; // @[Execute.scala 301:9]
  wire [63:0] _GEN_71; // @[Execute.scala 301:9]
  wire [63:0] _GEN_72; // @[Execute.scala 301:9]
  wire [63:0] _GEN_73; // @[Execute.scala 301:9]
  wire [63:0] _GEN_74; // @[Execute.scala 301:9]
  wire [63:0] _GEN_75; // @[Execute.scala 301:9]
  wire [63:0] _GEN_76; // @[Execute.scala 301:9]
  wire [63:0] _GEN_77; // @[Execute.scala 301:9]
  wire [63:0] _GEN_78; // @[Execute.scala 301:9]
  wire [63:0] _GEN_79; // @[Execute.scala 301:9]
  wire [63:0] _GEN_80; // @[Execute.scala 301:9]
  wire [63:0] _GEN_81; // @[Execute.scala 301:9]
  wire [63:0] _GEN_82; // @[Execute.scala 301:9]
  wire [63:0] _GEN_83; // @[Execute.scala 301:9]
  wire [63:0] _GEN_84; // @[Execute.scala 301:9]
  wire [63:0] _GEN_85; // @[Execute.scala 301:9]
  wire [63:0] _GEN_86; // @[Execute.scala 301:9]
  wire [63:0] _GEN_87; // @[Execute.scala 301:9]
  wire [63:0] _GEN_88; // @[Execute.scala 301:9]
  wire [63:0] _GEN_89; // @[Execute.scala 301:9]
  wire [63:0] _GEN_90; // @[Execute.scala 301:9]
  wire [63:0] _GEN_91; // @[Execute.scala 301:9]
  wire [63:0] _GEN_92; // @[Execute.scala 301:9]
  wire [63:0] _GEN_93; // @[Execute.scala 301:9]
  wire [63:0] _GEN_94; // @[Execute.scala 301:9]
  wire [63:0] _GEN_95; // @[Execute.scala 301:9]
  wire [63:0] _GEN_96; // @[Execute.scala 301:9]
  wire [63:0] _GEN_97; // @[Execute.scala 301:9]
  wire [63:0] _GEN_98; // @[Execute.scala 301:9]
  wire [63:0] _GEN_99; // @[Execute.scala 301:9]
  wire [63:0] _GEN_100; // @[Execute.scala 301:9]
  wire [63:0] _GEN_101; // @[Execute.scala 301:9]
  wire [63:0] _GEN_102; // @[Execute.scala 301:9]
  wire [63:0] _GEN_103; // @[Execute.scala 301:9]
  wire [63:0] _GEN_104; // @[Execute.scala 301:9]
  wire [63:0] _GEN_105; // @[Execute.scala 301:9]
  wire [63:0] _GEN_106; // @[Execute.scala 301:9]
  wire [63:0] _GEN_107; // @[Execute.scala 301:9]
  wire [63:0] _GEN_108; // @[Execute.scala 301:9]
  wire [63:0] _GEN_109; // @[Execute.scala 301:9]
  wire [63:0] _GEN_110; // @[Execute.scala 301:9]
  wire [63:0] _GEN_111; // @[Execute.scala 301:9]
  wire [63:0] _GEN_112; // @[Execute.scala 301:9]
  wire [63:0] _GEN_113; // @[Execute.scala 301:9]
  wire [63:0] _GEN_114; // @[Execute.scala 301:9]
  wire [63:0] _GEN_115; // @[Execute.scala 301:9]
  wire [63:0] _GEN_116; // @[Execute.scala 301:9]
  wire [63:0] _GEN_117; // @[Execute.scala 301:9]
  wire [63:0] _GEN_118; // @[Execute.scala 301:9]
  wire [63:0] _GEN_119; // @[Execute.scala 301:9]
  wire [63:0] _GEN_120; // @[Execute.scala 301:9]
  wire [63:0] _GEN_121; // @[Execute.scala 301:9]
  wire [63:0] _GEN_122; // @[Execute.scala 301:9]
  wire [63:0] _GEN_123; // @[Execute.scala 301:9]
  wire [63:0] _GEN_124; // @[Execute.scala 301:9]
  wire [63:0] _GEN_125; // @[Execute.scala 301:9]
  wire [63:0] _GEN_126; // @[Execute.scala 301:9]
  wire [63:0] _GEN_127; // @[Execute.scala 301:9]
  wire [63:0] _GEN_128; // @[Execute.scala 301:9]
  wire [63:0] welem; // @[Execute.scala 301:9]
  wire [6:0] _GEN_10437; // @[Execute.scala 117:37]
  wire [6:0] _T_94; // @[Execute.scala 117:37]
  wire  _GEN_131; // @[Execute.scala 117:10]
  wire  _GEN_132; // @[Execute.scala 117:10]
  wire  _GEN_133; // @[Execute.scala 117:10]
  wire  _GEN_134; // @[Execute.scala 117:10]
  wire  _GEN_135; // @[Execute.scala 117:10]
  wire  _GEN_136; // @[Execute.scala 117:10]
  wire  _GEN_137; // @[Execute.scala 117:10]
  wire  _GEN_138; // @[Execute.scala 117:10]
  wire  _GEN_139; // @[Execute.scala 117:10]
  wire  _GEN_140; // @[Execute.scala 117:10]
  wire  _GEN_141; // @[Execute.scala 117:10]
  wire  _GEN_142; // @[Execute.scala 117:10]
  wire  _GEN_143; // @[Execute.scala 117:10]
  wire  _GEN_144; // @[Execute.scala 117:10]
  wire  _GEN_145; // @[Execute.scala 117:10]
  wire  _GEN_146; // @[Execute.scala 117:10]
  wire  _GEN_147; // @[Execute.scala 117:10]
  wire  _GEN_148; // @[Execute.scala 117:10]
  wire  _GEN_149; // @[Execute.scala 117:10]
  wire  _GEN_150; // @[Execute.scala 117:10]
  wire  _GEN_151; // @[Execute.scala 117:10]
  wire  _GEN_152; // @[Execute.scala 117:10]
  wire  _GEN_153; // @[Execute.scala 117:10]
  wire  _GEN_154; // @[Execute.scala 117:10]
  wire  _GEN_155; // @[Execute.scala 117:10]
  wire  _GEN_156; // @[Execute.scala 117:10]
  wire  _GEN_157; // @[Execute.scala 117:10]
  wire  _GEN_158; // @[Execute.scala 117:10]
  wire  _GEN_159; // @[Execute.scala 117:10]
  wire  _GEN_160; // @[Execute.scala 117:10]
  wire  _GEN_161; // @[Execute.scala 117:10]
  wire  _GEN_162; // @[Execute.scala 117:10]
  wire  _GEN_163; // @[Execute.scala 117:10]
  wire  _GEN_164; // @[Execute.scala 117:10]
  wire  _GEN_165; // @[Execute.scala 117:10]
  wire  _GEN_166; // @[Execute.scala 117:10]
  wire  _GEN_167; // @[Execute.scala 117:10]
  wire  _GEN_168; // @[Execute.scala 117:10]
  wire  _GEN_169; // @[Execute.scala 117:10]
  wire  _GEN_170; // @[Execute.scala 117:10]
  wire  _GEN_171; // @[Execute.scala 117:10]
  wire  _GEN_172; // @[Execute.scala 117:10]
  wire  _GEN_173; // @[Execute.scala 117:10]
  wire  _GEN_174; // @[Execute.scala 117:10]
  wire  _GEN_175; // @[Execute.scala 117:10]
  wire  _GEN_176; // @[Execute.scala 117:10]
  wire  _GEN_177; // @[Execute.scala 117:10]
  wire  _GEN_178; // @[Execute.scala 117:10]
  wire  _GEN_179; // @[Execute.scala 117:10]
  wire  _GEN_180; // @[Execute.scala 117:10]
  wire  _GEN_181; // @[Execute.scala 117:10]
  wire  _GEN_182; // @[Execute.scala 117:10]
  wire  _GEN_183; // @[Execute.scala 117:10]
  wire  _GEN_184; // @[Execute.scala 117:10]
  wire  _GEN_185; // @[Execute.scala 117:10]
  wire  _GEN_186; // @[Execute.scala 117:10]
  wire  _GEN_187; // @[Execute.scala 117:10]
  wire  _GEN_188; // @[Execute.scala 117:10]
  wire  _GEN_189; // @[Execute.scala 117:10]
  wire  _GEN_190; // @[Execute.scala 117:10]
  wire  _GEN_191; // @[Execute.scala 117:10]
  wire  _GEN_192; // @[Execute.scala 117:10]
  wire  _GEN_193; // @[Execute.scala 117:10]
  wire  _T_102; // @[Execute.scala 117:15]
  wire [5:0] _T_104; // @[Execute.scala 117:37]
  wire [5:0] _T_108; // @[Execute.scala 117:60]
  wire  _GEN_259; // @[Execute.scala 117:10]
  wire  _GEN_260; // @[Execute.scala 117:10]
  wire  _GEN_261; // @[Execute.scala 117:10]
  wire  _GEN_262; // @[Execute.scala 117:10]
  wire  _GEN_263; // @[Execute.scala 117:10]
  wire  _GEN_264; // @[Execute.scala 117:10]
  wire  _GEN_265; // @[Execute.scala 117:10]
  wire  _GEN_266; // @[Execute.scala 117:10]
  wire  _GEN_267; // @[Execute.scala 117:10]
  wire  _GEN_268; // @[Execute.scala 117:10]
  wire  _GEN_269; // @[Execute.scala 117:10]
  wire  _GEN_270; // @[Execute.scala 117:10]
  wire  _GEN_271; // @[Execute.scala 117:10]
  wire  _GEN_272; // @[Execute.scala 117:10]
  wire  _GEN_273; // @[Execute.scala 117:10]
  wire  _GEN_274; // @[Execute.scala 117:10]
  wire  _GEN_275; // @[Execute.scala 117:10]
  wire  _GEN_276; // @[Execute.scala 117:10]
  wire  _GEN_277; // @[Execute.scala 117:10]
  wire  _GEN_278; // @[Execute.scala 117:10]
  wire  _GEN_279; // @[Execute.scala 117:10]
  wire  _GEN_280; // @[Execute.scala 117:10]
  wire  _GEN_281; // @[Execute.scala 117:10]
  wire  _GEN_282; // @[Execute.scala 117:10]
  wire  _GEN_283; // @[Execute.scala 117:10]
  wire  _GEN_284; // @[Execute.scala 117:10]
  wire  _GEN_285; // @[Execute.scala 117:10]
  wire  _GEN_286; // @[Execute.scala 117:10]
  wire  _GEN_287; // @[Execute.scala 117:10]
  wire  _GEN_288; // @[Execute.scala 117:10]
  wire  _GEN_289; // @[Execute.scala 117:10]
  wire  _GEN_290; // @[Execute.scala 117:10]
  wire  _GEN_291; // @[Execute.scala 117:10]
  wire  _GEN_292; // @[Execute.scala 117:10]
  wire  _GEN_293; // @[Execute.scala 117:10]
  wire  _GEN_294; // @[Execute.scala 117:10]
  wire  _GEN_295; // @[Execute.scala 117:10]
  wire  _GEN_296; // @[Execute.scala 117:10]
  wire  _GEN_297; // @[Execute.scala 117:10]
  wire  _GEN_298; // @[Execute.scala 117:10]
  wire  _GEN_299; // @[Execute.scala 117:10]
  wire  _GEN_300; // @[Execute.scala 117:10]
  wire  _GEN_301; // @[Execute.scala 117:10]
  wire  _GEN_302; // @[Execute.scala 117:10]
  wire  _GEN_303; // @[Execute.scala 117:10]
  wire  _GEN_304; // @[Execute.scala 117:10]
  wire  _GEN_305; // @[Execute.scala 117:10]
  wire  _GEN_306; // @[Execute.scala 117:10]
  wire  _GEN_307; // @[Execute.scala 117:10]
  wire  _GEN_308; // @[Execute.scala 117:10]
  wire  _GEN_309; // @[Execute.scala 117:10]
  wire  _GEN_310; // @[Execute.scala 117:10]
  wire  _GEN_311; // @[Execute.scala 117:10]
  wire  _GEN_312; // @[Execute.scala 117:10]
  wire  _GEN_313; // @[Execute.scala 117:10]
  wire  _GEN_314; // @[Execute.scala 117:10]
  wire  _GEN_315; // @[Execute.scala 117:10]
  wire  _GEN_316; // @[Execute.scala 117:10]
  wire  _GEN_317; // @[Execute.scala 117:10]
  wire  _GEN_318; // @[Execute.scala 117:10]
  wire  _GEN_319; // @[Execute.scala 117:10]
  wire  _GEN_320; // @[Execute.scala 117:10]
  wire  _GEN_321; // @[Execute.scala 117:10]
  wire  _GEN_323; // @[Execute.scala 117:10]
  wire  _GEN_324; // @[Execute.scala 117:10]
  wire  _GEN_325; // @[Execute.scala 117:10]
  wire  _GEN_326; // @[Execute.scala 117:10]
  wire  _GEN_327; // @[Execute.scala 117:10]
  wire  _GEN_328; // @[Execute.scala 117:10]
  wire  _GEN_329; // @[Execute.scala 117:10]
  wire  _GEN_330; // @[Execute.scala 117:10]
  wire  _GEN_331; // @[Execute.scala 117:10]
  wire  _GEN_332; // @[Execute.scala 117:10]
  wire  _GEN_333; // @[Execute.scala 117:10]
  wire  _GEN_334; // @[Execute.scala 117:10]
  wire  _GEN_335; // @[Execute.scala 117:10]
  wire  _GEN_336; // @[Execute.scala 117:10]
  wire  _GEN_337; // @[Execute.scala 117:10]
  wire  _GEN_338; // @[Execute.scala 117:10]
  wire  _GEN_339; // @[Execute.scala 117:10]
  wire  _GEN_340; // @[Execute.scala 117:10]
  wire  _GEN_341; // @[Execute.scala 117:10]
  wire  _GEN_342; // @[Execute.scala 117:10]
  wire  _GEN_343; // @[Execute.scala 117:10]
  wire  _GEN_344; // @[Execute.scala 117:10]
  wire  _GEN_345; // @[Execute.scala 117:10]
  wire  _GEN_346; // @[Execute.scala 117:10]
  wire  _GEN_347; // @[Execute.scala 117:10]
  wire  _GEN_348; // @[Execute.scala 117:10]
  wire  _GEN_349; // @[Execute.scala 117:10]
  wire  _GEN_350; // @[Execute.scala 117:10]
  wire  _GEN_351; // @[Execute.scala 117:10]
  wire  _GEN_352; // @[Execute.scala 117:10]
  wire  _GEN_353; // @[Execute.scala 117:10]
  wire  _GEN_354; // @[Execute.scala 117:10]
  wire  _GEN_355; // @[Execute.scala 117:10]
  wire  _GEN_356; // @[Execute.scala 117:10]
  wire  _GEN_357; // @[Execute.scala 117:10]
  wire  _GEN_358; // @[Execute.scala 117:10]
  wire  _GEN_359; // @[Execute.scala 117:10]
  wire  _GEN_360; // @[Execute.scala 117:10]
  wire  _GEN_361; // @[Execute.scala 117:10]
  wire  _GEN_362; // @[Execute.scala 117:10]
  wire  _GEN_363; // @[Execute.scala 117:10]
  wire  _GEN_364; // @[Execute.scala 117:10]
  wire  _GEN_365; // @[Execute.scala 117:10]
  wire  _GEN_366; // @[Execute.scala 117:10]
  wire  _GEN_367; // @[Execute.scala 117:10]
  wire  _GEN_368; // @[Execute.scala 117:10]
  wire  _GEN_369; // @[Execute.scala 117:10]
  wire  _GEN_370; // @[Execute.scala 117:10]
  wire  _GEN_371; // @[Execute.scala 117:10]
  wire  _GEN_372; // @[Execute.scala 117:10]
  wire  _GEN_373; // @[Execute.scala 117:10]
  wire  _GEN_374; // @[Execute.scala 117:10]
  wire  _GEN_375; // @[Execute.scala 117:10]
  wire  _GEN_376; // @[Execute.scala 117:10]
  wire  _GEN_377; // @[Execute.scala 117:10]
  wire  _GEN_378; // @[Execute.scala 117:10]
  wire  _GEN_379; // @[Execute.scala 117:10]
  wire  _GEN_380; // @[Execute.scala 117:10]
  wire  _GEN_381; // @[Execute.scala 117:10]
  wire  _GEN_382; // @[Execute.scala 117:10]
  wire  _GEN_383; // @[Execute.scala 117:10]
  wire  _GEN_384; // @[Execute.scala 117:10]
  wire  _GEN_385; // @[Execute.scala 117:10]
  wire  _T_111; // @[Execute.scala 117:10]
  wire  _T_112; // @[Execute.scala 117:15]
  wire [5:0] _T_114; // @[Execute.scala 117:37]
  wire [5:0] _T_118; // @[Execute.scala 117:60]
  wire  _GEN_387; // @[Execute.scala 117:10]
  wire  _GEN_388; // @[Execute.scala 117:10]
  wire  _GEN_389; // @[Execute.scala 117:10]
  wire  _GEN_390; // @[Execute.scala 117:10]
  wire  _GEN_391; // @[Execute.scala 117:10]
  wire  _GEN_392; // @[Execute.scala 117:10]
  wire  _GEN_393; // @[Execute.scala 117:10]
  wire  _GEN_394; // @[Execute.scala 117:10]
  wire  _GEN_395; // @[Execute.scala 117:10]
  wire  _GEN_396; // @[Execute.scala 117:10]
  wire  _GEN_397; // @[Execute.scala 117:10]
  wire  _GEN_398; // @[Execute.scala 117:10]
  wire  _GEN_399; // @[Execute.scala 117:10]
  wire  _GEN_400; // @[Execute.scala 117:10]
  wire  _GEN_401; // @[Execute.scala 117:10]
  wire  _GEN_402; // @[Execute.scala 117:10]
  wire  _GEN_403; // @[Execute.scala 117:10]
  wire  _GEN_404; // @[Execute.scala 117:10]
  wire  _GEN_405; // @[Execute.scala 117:10]
  wire  _GEN_406; // @[Execute.scala 117:10]
  wire  _GEN_407; // @[Execute.scala 117:10]
  wire  _GEN_408; // @[Execute.scala 117:10]
  wire  _GEN_409; // @[Execute.scala 117:10]
  wire  _GEN_410; // @[Execute.scala 117:10]
  wire  _GEN_411; // @[Execute.scala 117:10]
  wire  _GEN_412; // @[Execute.scala 117:10]
  wire  _GEN_413; // @[Execute.scala 117:10]
  wire  _GEN_414; // @[Execute.scala 117:10]
  wire  _GEN_415; // @[Execute.scala 117:10]
  wire  _GEN_416; // @[Execute.scala 117:10]
  wire  _GEN_417; // @[Execute.scala 117:10]
  wire  _GEN_418; // @[Execute.scala 117:10]
  wire  _GEN_419; // @[Execute.scala 117:10]
  wire  _GEN_420; // @[Execute.scala 117:10]
  wire  _GEN_421; // @[Execute.scala 117:10]
  wire  _GEN_422; // @[Execute.scala 117:10]
  wire  _GEN_423; // @[Execute.scala 117:10]
  wire  _GEN_424; // @[Execute.scala 117:10]
  wire  _GEN_425; // @[Execute.scala 117:10]
  wire  _GEN_426; // @[Execute.scala 117:10]
  wire  _GEN_427; // @[Execute.scala 117:10]
  wire  _GEN_428; // @[Execute.scala 117:10]
  wire  _GEN_429; // @[Execute.scala 117:10]
  wire  _GEN_430; // @[Execute.scala 117:10]
  wire  _GEN_431; // @[Execute.scala 117:10]
  wire  _GEN_432; // @[Execute.scala 117:10]
  wire  _GEN_433; // @[Execute.scala 117:10]
  wire  _GEN_434; // @[Execute.scala 117:10]
  wire  _GEN_435; // @[Execute.scala 117:10]
  wire  _GEN_436; // @[Execute.scala 117:10]
  wire  _GEN_437; // @[Execute.scala 117:10]
  wire  _GEN_438; // @[Execute.scala 117:10]
  wire  _GEN_439; // @[Execute.scala 117:10]
  wire  _GEN_440; // @[Execute.scala 117:10]
  wire  _GEN_441; // @[Execute.scala 117:10]
  wire  _GEN_442; // @[Execute.scala 117:10]
  wire  _GEN_443; // @[Execute.scala 117:10]
  wire  _GEN_444; // @[Execute.scala 117:10]
  wire  _GEN_445; // @[Execute.scala 117:10]
  wire  _GEN_446; // @[Execute.scala 117:10]
  wire  _GEN_447; // @[Execute.scala 117:10]
  wire  _GEN_448; // @[Execute.scala 117:10]
  wire  _GEN_449; // @[Execute.scala 117:10]
  wire  _GEN_451; // @[Execute.scala 117:10]
  wire  _GEN_452; // @[Execute.scala 117:10]
  wire  _GEN_453; // @[Execute.scala 117:10]
  wire  _GEN_454; // @[Execute.scala 117:10]
  wire  _GEN_455; // @[Execute.scala 117:10]
  wire  _GEN_456; // @[Execute.scala 117:10]
  wire  _GEN_457; // @[Execute.scala 117:10]
  wire  _GEN_458; // @[Execute.scala 117:10]
  wire  _GEN_459; // @[Execute.scala 117:10]
  wire  _GEN_460; // @[Execute.scala 117:10]
  wire  _GEN_461; // @[Execute.scala 117:10]
  wire  _GEN_462; // @[Execute.scala 117:10]
  wire  _GEN_463; // @[Execute.scala 117:10]
  wire  _GEN_464; // @[Execute.scala 117:10]
  wire  _GEN_465; // @[Execute.scala 117:10]
  wire  _GEN_466; // @[Execute.scala 117:10]
  wire  _GEN_467; // @[Execute.scala 117:10]
  wire  _GEN_468; // @[Execute.scala 117:10]
  wire  _GEN_469; // @[Execute.scala 117:10]
  wire  _GEN_470; // @[Execute.scala 117:10]
  wire  _GEN_471; // @[Execute.scala 117:10]
  wire  _GEN_472; // @[Execute.scala 117:10]
  wire  _GEN_473; // @[Execute.scala 117:10]
  wire  _GEN_474; // @[Execute.scala 117:10]
  wire  _GEN_475; // @[Execute.scala 117:10]
  wire  _GEN_476; // @[Execute.scala 117:10]
  wire  _GEN_477; // @[Execute.scala 117:10]
  wire  _GEN_478; // @[Execute.scala 117:10]
  wire  _GEN_479; // @[Execute.scala 117:10]
  wire  _GEN_480; // @[Execute.scala 117:10]
  wire  _GEN_481; // @[Execute.scala 117:10]
  wire  _GEN_482; // @[Execute.scala 117:10]
  wire  _GEN_483; // @[Execute.scala 117:10]
  wire  _GEN_484; // @[Execute.scala 117:10]
  wire  _GEN_485; // @[Execute.scala 117:10]
  wire  _GEN_486; // @[Execute.scala 117:10]
  wire  _GEN_487; // @[Execute.scala 117:10]
  wire  _GEN_488; // @[Execute.scala 117:10]
  wire  _GEN_489; // @[Execute.scala 117:10]
  wire  _GEN_490; // @[Execute.scala 117:10]
  wire  _GEN_491; // @[Execute.scala 117:10]
  wire  _GEN_492; // @[Execute.scala 117:10]
  wire  _GEN_493; // @[Execute.scala 117:10]
  wire  _GEN_494; // @[Execute.scala 117:10]
  wire  _GEN_495; // @[Execute.scala 117:10]
  wire  _GEN_496; // @[Execute.scala 117:10]
  wire  _GEN_497; // @[Execute.scala 117:10]
  wire  _GEN_498; // @[Execute.scala 117:10]
  wire  _GEN_499; // @[Execute.scala 117:10]
  wire  _GEN_500; // @[Execute.scala 117:10]
  wire  _GEN_501; // @[Execute.scala 117:10]
  wire  _GEN_502; // @[Execute.scala 117:10]
  wire  _GEN_503; // @[Execute.scala 117:10]
  wire  _GEN_504; // @[Execute.scala 117:10]
  wire  _GEN_505; // @[Execute.scala 117:10]
  wire  _GEN_506; // @[Execute.scala 117:10]
  wire  _GEN_507; // @[Execute.scala 117:10]
  wire  _GEN_508; // @[Execute.scala 117:10]
  wire  _GEN_509; // @[Execute.scala 117:10]
  wire  _GEN_510; // @[Execute.scala 117:10]
  wire  _GEN_511; // @[Execute.scala 117:10]
  wire  _GEN_512; // @[Execute.scala 117:10]
  wire  _GEN_513; // @[Execute.scala 117:10]
  wire  _T_121; // @[Execute.scala 117:10]
  wire  _T_122; // @[Execute.scala 117:15]
  wire [5:0] _T_124; // @[Execute.scala 117:37]
  wire [5:0] _T_128; // @[Execute.scala 117:60]
  wire  _GEN_515; // @[Execute.scala 117:10]
  wire  _GEN_516; // @[Execute.scala 117:10]
  wire  _GEN_517; // @[Execute.scala 117:10]
  wire  _GEN_518; // @[Execute.scala 117:10]
  wire  _GEN_519; // @[Execute.scala 117:10]
  wire  _GEN_520; // @[Execute.scala 117:10]
  wire  _GEN_521; // @[Execute.scala 117:10]
  wire  _GEN_522; // @[Execute.scala 117:10]
  wire  _GEN_523; // @[Execute.scala 117:10]
  wire  _GEN_524; // @[Execute.scala 117:10]
  wire  _GEN_525; // @[Execute.scala 117:10]
  wire  _GEN_526; // @[Execute.scala 117:10]
  wire  _GEN_527; // @[Execute.scala 117:10]
  wire  _GEN_528; // @[Execute.scala 117:10]
  wire  _GEN_529; // @[Execute.scala 117:10]
  wire  _GEN_530; // @[Execute.scala 117:10]
  wire  _GEN_531; // @[Execute.scala 117:10]
  wire  _GEN_532; // @[Execute.scala 117:10]
  wire  _GEN_533; // @[Execute.scala 117:10]
  wire  _GEN_534; // @[Execute.scala 117:10]
  wire  _GEN_535; // @[Execute.scala 117:10]
  wire  _GEN_536; // @[Execute.scala 117:10]
  wire  _GEN_537; // @[Execute.scala 117:10]
  wire  _GEN_538; // @[Execute.scala 117:10]
  wire  _GEN_539; // @[Execute.scala 117:10]
  wire  _GEN_540; // @[Execute.scala 117:10]
  wire  _GEN_541; // @[Execute.scala 117:10]
  wire  _GEN_542; // @[Execute.scala 117:10]
  wire  _GEN_543; // @[Execute.scala 117:10]
  wire  _GEN_544; // @[Execute.scala 117:10]
  wire  _GEN_545; // @[Execute.scala 117:10]
  wire  _GEN_546; // @[Execute.scala 117:10]
  wire  _GEN_547; // @[Execute.scala 117:10]
  wire  _GEN_548; // @[Execute.scala 117:10]
  wire  _GEN_549; // @[Execute.scala 117:10]
  wire  _GEN_550; // @[Execute.scala 117:10]
  wire  _GEN_551; // @[Execute.scala 117:10]
  wire  _GEN_552; // @[Execute.scala 117:10]
  wire  _GEN_553; // @[Execute.scala 117:10]
  wire  _GEN_554; // @[Execute.scala 117:10]
  wire  _GEN_555; // @[Execute.scala 117:10]
  wire  _GEN_556; // @[Execute.scala 117:10]
  wire  _GEN_557; // @[Execute.scala 117:10]
  wire  _GEN_558; // @[Execute.scala 117:10]
  wire  _GEN_559; // @[Execute.scala 117:10]
  wire  _GEN_560; // @[Execute.scala 117:10]
  wire  _GEN_561; // @[Execute.scala 117:10]
  wire  _GEN_562; // @[Execute.scala 117:10]
  wire  _GEN_563; // @[Execute.scala 117:10]
  wire  _GEN_564; // @[Execute.scala 117:10]
  wire  _GEN_565; // @[Execute.scala 117:10]
  wire  _GEN_566; // @[Execute.scala 117:10]
  wire  _GEN_567; // @[Execute.scala 117:10]
  wire  _GEN_568; // @[Execute.scala 117:10]
  wire  _GEN_569; // @[Execute.scala 117:10]
  wire  _GEN_570; // @[Execute.scala 117:10]
  wire  _GEN_571; // @[Execute.scala 117:10]
  wire  _GEN_572; // @[Execute.scala 117:10]
  wire  _GEN_573; // @[Execute.scala 117:10]
  wire  _GEN_574; // @[Execute.scala 117:10]
  wire  _GEN_575; // @[Execute.scala 117:10]
  wire  _GEN_576; // @[Execute.scala 117:10]
  wire  _GEN_577; // @[Execute.scala 117:10]
  wire  _GEN_579; // @[Execute.scala 117:10]
  wire  _GEN_580; // @[Execute.scala 117:10]
  wire  _GEN_581; // @[Execute.scala 117:10]
  wire  _GEN_582; // @[Execute.scala 117:10]
  wire  _GEN_583; // @[Execute.scala 117:10]
  wire  _GEN_584; // @[Execute.scala 117:10]
  wire  _GEN_585; // @[Execute.scala 117:10]
  wire  _GEN_586; // @[Execute.scala 117:10]
  wire  _GEN_587; // @[Execute.scala 117:10]
  wire  _GEN_588; // @[Execute.scala 117:10]
  wire  _GEN_589; // @[Execute.scala 117:10]
  wire  _GEN_590; // @[Execute.scala 117:10]
  wire  _GEN_591; // @[Execute.scala 117:10]
  wire  _GEN_592; // @[Execute.scala 117:10]
  wire  _GEN_593; // @[Execute.scala 117:10]
  wire  _GEN_594; // @[Execute.scala 117:10]
  wire  _GEN_595; // @[Execute.scala 117:10]
  wire  _GEN_596; // @[Execute.scala 117:10]
  wire  _GEN_597; // @[Execute.scala 117:10]
  wire  _GEN_598; // @[Execute.scala 117:10]
  wire  _GEN_599; // @[Execute.scala 117:10]
  wire  _GEN_600; // @[Execute.scala 117:10]
  wire  _GEN_601; // @[Execute.scala 117:10]
  wire  _GEN_602; // @[Execute.scala 117:10]
  wire  _GEN_603; // @[Execute.scala 117:10]
  wire  _GEN_604; // @[Execute.scala 117:10]
  wire  _GEN_605; // @[Execute.scala 117:10]
  wire  _GEN_606; // @[Execute.scala 117:10]
  wire  _GEN_607; // @[Execute.scala 117:10]
  wire  _GEN_608; // @[Execute.scala 117:10]
  wire  _GEN_609; // @[Execute.scala 117:10]
  wire  _GEN_610; // @[Execute.scala 117:10]
  wire  _GEN_611; // @[Execute.scala 117:10]
  wire  _GEN_612; // @[Execute.scala 117:10]
  wire  _GEN_613; // @[Execute.scala 117:10]
  wire  _GEN_614; // @[Execute.scala 117:10]
  wire  _GEN_615; // @[Execute.scala 117:10]
  wire  _GEN_616; // @[Execute.scala 117:10]
  wire  _GEN_617; // @[Execute.scala 117:10]
  wire  _GEN_618; // @[Execute.scala 117:10]
  wire  _GEN_619; // @[Execute.scala 117:10]
  wire  _GEN_620; // @[Execute.scala 117:10]
  wire  _GEN_621; // @[Execute.scala 117:10]
  wire  _GEN_622; // @[Execute.scala 117:10]
  wire  _GEN_623; // @[Execute.scala 117:10]
  wire  _GEN_624; // @[Execute.scala 117:10]
  wire  _GEN_625; // @[Execute.scala 117:10]
  wire  _GEN_626; // @[Execute.scala 117:10]
  wire  _GEN_627; // @[Execute.scala 117:10]
  wire  _GEN_628; // @[Execute.scala 117:10]
  wire  _GEN_629; // @[Execute.scala 117:10]
  wire  _GEN_630; // @[Execute.scala 117:10]
  wire  _GEN_631; // @[Execute.scala 117:10]
  wire  _GEN_632; // @[Execute.scala 117:10]
  wire  _GEN_633; // @[Execute.scala 117:10]
  wire  _GEN_634; // @[Execute.scala 117:10]
  wire  _GEN_635; // @[Execute.scala 117:10]
  wire  _GEN_636; // @[Execute.scala 117:10]
  wire  _GEN_637; // @[Execute.scala 117:10]
  wire  _GEN_638; // @[Execute.scala 117:10]
  wire  _GEN_639; // @[Execute.scala 117:10]
  wire  _GEN_640; // @[Execute.scala 117:10]
  wire  _GEN_641; // @[Execute.scala 117:10]
  wire  _T_131; // @[Execute.scala 117:10]
  wire  _T_132; // @[Execute.scala 117:15]
  wire [5:0] _T_134; // @[Execute.scala 117:37]
  wire [5:0] _T_138; // @[Execute.scala 117:60]
  wire  _GEN_643; // @[Execute.scala 117:10]
  wire  _GEN_644; // @[Execute.scala 117:10]
  wire  _GEN_645; // @[Execute.scala 117:10]
  wire  _GEN_646; // @[Execute.scala 117:10]
  wire  _GEN_647; // @[Execute.scala 117:10]
  wire  _GEN_648; // @[Execute.scala 117:10]
  wire  _GEN_649; // @[Execute.scala 117:10]
  wire  _GEN_650; // @[Execute.scala 117:10]
  wire  _GEN_651; // @[Execute.scala 117:10]
  wire  _GEN_652; // @[Execute.scala 117:10]
  wire  _GEN_653; // @[Execute.scala 117:10]
  wire  _GEN_654; // @[Execute.scala 117:10]
  wire  _GEN_655; // @[Execute.scala 117:10]
  wire  _GEN_656; // @[Execute.scala 117:10]
  wire  _GEN_657; // @[Execute.scala 117:10]
  wire  _GEN_658; // @[Execute.scala 117:10]
  wire  _GEN_659; // @[Execute.scala 117:10]
  wire  _GEN_660; // @[Execute.scala 117:10]
  wire  _GEN_661; // @[Execute.scala 117:10]
  wire  _GEN_662; // @[Execute.scala 117:10]
  wire  _GEN_663; // @[Execute.scala 117:10]
  wire  _GEN_664; // @[Execute.scala 117:10]
  wire  _GEN_665; // @[Execute.scala 117:10]
  wire  _GEN_666; // @[Execute.scala 117:10]
  wire  _GEN_667; // @[Execute.scala 117:10]
  wire  _GEN_668; // @[Execute.scala 117:10]
  wire  _GEN_669; // @[Execute.scala 117:10]
  wire  _GEN_670; // @[Execute.scala 117:10]
  wire  _GEN_671; // @[Execute.scala 117:10]
  wire  _GEN_672; // @[Execute.scala 117:10]
  wire  _GEN_673; // @[Execute.scala 117:10]
  wire  _GEN_674; // @[Execute.scala 117:10]
  wire  _GEN_675; // @[Execute.scala 117:10]
  wire  _GEN_676; // @[Execute.scala 117:10]
  wire  _GEN_677; // @[Execute.scala 117:10]
  wire  _GEN_678; // @[Execute.scala 117:10]
  wire  _GEN_679; // @[Execute.scala 117:10]
  wire  _GEN_680; // @[Execute.scala 117:10]
  wire  _GEN_681; // @[Execute.scala 117:10]
  wire  _GEN_682; // @[Execute.scala 117:10]
  wire  _GEN_683; // @[Execute.scala 117:10]
  wire  _GEN_684; // @[Execute.scala 117:10]
  wire  _GEN_685; // @[Execute.scala 117:10]
  wire  _GEN_686; // @[Execute.scala 117:10]
  wire  _GEN_687; // @[Execute.scala 117:10]
  wire  _GEN_688; // @[Execute.scala 117:10]
  wire  _GEN_689; // @[Execute.scala 117:10]
  wire  _GEN_690; // @[Execute.scala 117:10]
  wire  _GEN_691; // @[Execute.scala 117:10]
  wire  _GEN_692; // @[Execute.scala 117:10]
  wire  _GEN_693; // @[Execute.scala 117:10]
  wire  _GEN_694; // @[Execute.scala 117:10]
  wire  _GEN_695; // @[Execute.scala 117:10]
  wire  _GEN_696; // @[Execute.scala 117:10]
  wire  _GEN_697; // @[Execute.scala 117:10]
  wire  _GEN_698; // @[Execute.scala 117:10]
  wire  _GEN_699; // @[Execute.scala 117:10]
  wire  _GEN_700; // @[Execute.scala 117:10]
  wire  _GEN_701; // @[Execute.scala 117:10]
  wire  _GEN_702; // @[Execute.scala 117:10]
  wire  _GEN_703; // @[Execute.scala 117:10]
  wire  _GEN_704; // @[Execute.scala 117:10]
  wire  _GEN_705; // @[Execute.scala 117:10]
  wire  _GEN_707; // @[Execute.scala 117:10]
  wire  _GEN_708; // @[Execute.scala 117:10]
  wire  _GEN_709; // @[Execute.scala 117:10]
  wire  _GEN_710; // @[Execute.scala 117:10]
  wire  _GEN_711; // @[Execute.scala 117:10]
  wire  _GEN_712; // @[Execute.scala 117:10]
  wire  _GEN_713; // @[Execute.scala 117:10]
  wire  _GEN_714; // @[Execute.scala 117:10]
  wire  _GEN_715; // @[Execute.scala 117:10]
  wire  _GEN_716; // @[Execute.scala 117:10]
  wire  _GEN_717; // @[Execute.scala 117:10]
  wire  _GEN_718; // @[Execute.scala 117:10]
  wire  _GEN_719; // @[Execute.scala 117:10]
  wire  _GEN_720; // @[Execute.scala 117:10]
  wire  _GEN_721; // @[Execute.scala 117:10]
  wire  _GEN_722; // @[Execute.scala 117:10]
  wire  _GEN_723; // @[Execute.scala 117:10]
  wire  _GEN_724; // @[Execute.scala 117:10]
  wire  _GEN_725; // @[Execute.scala 117:10]
  wire  _GEN_726; // @[Execute.scala 117:10]
  wire  _GEN_727; // @[Execute.scala 117:10]
  wire  _GEN_728; // @[Execute.scala 117:10]
  wire  _GEN_729; // @[Execute.scala 117:10]
  wire  _GEN_730; // @[Execute.scala 117:10]
  wire  _GEN_731; // @[Execute.scala 117:10]
  wire  _GEN_732; // @[Execute.scala 117:10]
  wire  _GEN_733; // @[Execute.scala 117:10]
  wire  _GEN_734; // @[Execute.scala 117:10]
  wire  _GEN_735; // @[Execute.scala 117:10]
  wire  _GEN_736; // @[Execute.scala 117:10]
  wire  _GEN_737; // @[Execute.scala 117:10]
  wire  _GEN_738; // @[Execute.scala 117:10]
  wire  _GEN_739; // @[Execute.scala 117:10]
  wire  _GEN_740; // @[Execute.scala 117:10]
  wire  _GEN_741; // @[Execute.scala 117:10]
  wire  _GEN_742; // @[Execute.scala 117:10]
  wire  _GEN_743; // @[Execute.scala 117:10]
  wire  _GEN_744; // @[Execute.scala 117:10]
  wire  _GEN_745; // @[Execute.scala 117:10]
  wire  _GEN_746; // @[Execute.scala 117:10]
  wire  _GEN_747; // @[Execute.scala 117:10]
  wire  _GEN_748; // @[Execute.scala 117:10]
  wire  _GEN_749; // @[Execute.scala 117:10]
  wire  _GEN_750; // @[Execute.scala 117:10]
  wire  _GEN_751; // @[Execute.scala 117:10]
  wire  _GEN_752; // @[Execute.scala 117:10]
  wire  _GEN_753; // @[Execute.scala 117:10]
  wire  _GEN_754; // @[Execute.scala 117:10]
  wire  _GEN_755; // @[Execute.scala 117:10]
  wire  _GEN_756; // @[Execute.scala 117:10]
  wire  _GEN_757; // @[Execute.scala 117:10]
  wire  _GEN_758; // @[Execute.scala 117:10]
  wire  _GEN_759; // @[Execute.scala 117:10]
  wire  _GEN_760; // @[Execute.scala 117:10]
  wire  _GEN_761; // @[Execute.scala 117:10]
  wire  _GEN_762; // @[Execute.scala 117:10]
  wire  _GEN_763; // @[Execute.scala 117:10]
  wire  _GEN_764; // @[Execute.scala 117:10]
  wire  _GEN_765; // @[Execute.scala 117:10]
  wire  _GEN_766; // @[Execute.scala 117:10]
  wire  _GEN_767; // @[Execute.scala 117:10]
  wire  _GEN_768; // @[Execute.scala 117:10]
  wire  _GEN_769; // @[Execute.scala 117:10]
  wire  _T_141; // @[Execute.scala 117:10]
  wire  _T_142; // @[Execute.scala 117:15]
  wire [5:0] _T_144; // @[Execute.scala 117:37]
  wire [5:0] _T_148; // @[Execute.scala 117:60]
  wire  _GEN_771; // @[Execute.scala 117:10]
  wire  _GEN_772; // @[Execute.scala 117:10]
  wire  _GEN_773; // @[Execute.scala 117:10]
  wire  _GEN_774; // @[Execute.scala 117:10]
  wire  _GEN_775; // @[Execute.scala 117:10]
  wire  _GEN_776; // @[Execute.scala 117:10]
  wire  _GEN_777; // @[Execute.scala 117:10]
  wire  _GEN_778; // @[Execute.scala 117:10]
  wire  _GEN_779; // @[Execute.scala 117:10]
  wire  _GEN_780; // @[Execute.scala 117:10]
  wire  _GEN_781; // @[Execute.scala 117:10]
  wire  _GEN_782; // @[Execute.scala 117:10]
  wire  _GEN_783; // @[Execute.scala 117:10]
  wire  _GEN_784; // @[Execute.scala 117:10]
  wire  _GEN_785; // @[Execute.scala 117:10]
  wire  _GEN_786; // @[Execute.scala 117:10]
  wire  _GEN_787; // @[Execute.scala 117:10]
  wire  _GEN_788; // @[Execute.scala 117:10]
  wire  _GEN_789; // @[Execute.scala 117:10]
  wire  _GEN_790; // @[Execute.scala 117:10]
  wire  _GEN_791; // @[Execute.scala 117:10]
  wire  _GEN_792; // @[Execute.scala 117:10]
  wire  _GEN_793; // @[Execute.scala 117:10]
  wire  _GEN_794; // @[Execute.scala 117:10]
  wire  _GEN_795; // @[Execute.scala 117:10]
  wire  _GEN_796; // @[Execute.scala 117:10]
  wire  _GEN_797; // @[Execute.scala 117:10]
  wire  _GEN_798; // @[Execute.scala 117:10]
  wire  _GEN_799; // @[Execute.scala 117:10]
  wire  _GEN_800; // @[Execute.scala 117:10]
  wire  _GEN_801; // @[Execute.scala 117:10]
  wire  _GEN_802; // @[Execute.scala 117:10]
  wire  _GEN_803; // @[Execute.scala 117:10]
  wire  _GEN_804; // @[Execute.scala 117:10]
  wire  _GEN_805; // @[Execute.scala 117:10]
  wire  _GEN_806; // @[Execute.scala 117:10]
  wire  _GEN_807; // @[Execute.scala 117:10]
  wire  _GEN_808; // @[Execute.scala 117:10]
  wire  _GEN_809; // @[Execute.scala 117:10]
  wire  _GEN_810; // @[Execute.scala 117:10]
  wire  _GEN_811; // @[Execute.scala 117:10]
  wire  _GEN_812; // @[Execute.scala 117:10]
  wire  _GEN_813; // @[Execute.scala 117:10]
  wire  _GEN_814; // @[Execute.scala 117:10]
  wire  _GEN_815; // @[Execute.scala 117:10]
  wire  _GEN_816; // @[Execute.scala 117:10]
  wire  _GEN_817; // @[Execute.scala 117:10]
  wire  _GEN_818; // @[Execute.scala 117:10]
  wire  _GEN_819; // @[Execute.scala 117:10]
  wire  _GEN_820; // @[Execute.scala 117:10]
  wire  _GEN_821; // @[Execute.scala 117:10]
  wire  _GEN_822; // @[Execute.scala 117:10]
  wire  _GEN_823; // @[Execute.scala 117:10]
  wire  _GEN_824; // @[Execute.scala 117:10]
  wire  _GEN_825; // @[Execute.scala 117:10]
  wire  _GEN_826; // @[Execute.scala 117:10]
  wire  _GEN_827; // @[Execute.scala 117:10]
  wire  _GEN_828; // @[Execute.scala 117:10]
  wire  _GEN_829; // @[Execute.scala 117:10]
  wire  _GEN_830; // @[Execute.scala 117:10]
  wire  _GEN_831; // @[Execute.scala 117:10]
  wire  _GEN_832; // @[Execute.scala 117:10]
  wire  _GEN_833; // @[Execute.scala 117:10]
  wire  _GEN_835; // @[Execute.scala 117:10]
  wire  _GEN_836; // @[Execute.scala 117:10]
  wire  _GEN_837; // @[Execute.scala 117:10]
  wire  _GEN_838; // @[Execute.scala 117:10]
  wire  _GEN_839; // @[Execute.scala 117:10]
  wire  _GEN_840; // @[Execute.scala 117:10]
  wire  _GEN_841; // @[Execute.scala 117:10]
  wire  _GEN_842; // @[Execute.scala 117:10]
  wire  _GEN_843; // @[Execute.scala 117:10]
  wire  _GEN_844; // @[Execute.scala 117:10]
  wire  _GEN_845; // @[Execute.scala 117:10]
  wire  _GEN_846; // @[Execute.scala 117:10]
  wire  _GEN_847; // @[Execute.scala 117:10]
  wire  _GEN_848; // @[Execute.scala 117:10]
  wire  _GEN_849; // @[Execute.scala 117:10]
  wire  _GEN_850; // @[Execute.scala 117:10]
  wire  _GEN_851; // @[Execute.scala 117:10]
  wire  _GEN_852; // @[Execute.scala 117:10]
  wire  _GEN_853; // @[Execute.scala 117:10]
  wire  _GEN_854; // @[Execute.scala 117:10]
  wire  _GEN_855; // @[Execute.scala 117:10]
  wire  _GEN_856; // @[Execute.scala 117:10]
  wire  _GEN_857; // @[Execute.scala 117:10]
  wire  _GEN_858; // @[Execute.scala 117:10]
  wire  _GEN_859; // @[Execute.scala 117:10]
  wire  _GEN_860; // @[Execute.scala 117:10]
  wire  _GEN_861; // @[Execute.scala 117:10]
  wire  _GEN_862; // @[Execute.scala 117:10]
  wire  _GEN_863; // @[Execute.scala 117:10]
  wire  _GEN_864; // @[Execute.scala 117:10]
  wire  _GEN_865; // @[Execute.scala 117:10]
  wire  _GEN_866; // @[Execute.scala 117:10]
  wire  _GEN_867; // @[Execute.scala 117:10]
  wire  _GEN_868; // @[Execute.scala 117:10]
  wire  _GEN_869; // @[Execute.scala 117:10]
  wire  _GEN_870; // @[Execute.scala 117:10]
  wire  _GEN_871; // @[Execute.scala 117:10]
  wire  _GEN_872; // @[Execute.scala 117:10]
  wire  _GEN_873; // @[Execute.scala 117:10]
  wire  _GEN_874; // @[Execute.scala 117:10]
  wire  _GEN_875; // @[Execute.scala 117:10]
  wire  _GEN_876; // @[Execute.scala 117:10]
  wire  _GEN_877; // @[Execute.scala 117:10]
  wire  _GEN_878; // @[Execute.scala 117:10]
  wire  _GEN_879; // @[Execute.scala 117:10]
  wire  _GEN_880; // @[Execute.scala 117:10]
  wire  _GEN_881; // @[Execute.scala 117:10]
  wire  _GEN_882; // @[Execute.scala 117:10]
  wire  _GEN_883; // @[Execute.scala 117:10]
  wire  _GEN_884; // @[Execute.scala 117:10]
  wire  _GEN_885; // @[Execute.scala 117:10]
  wire  _GEN_886; // @[Execute.scala 117:10]
  wire  _GEN_887; // @[Execute.scala 117:10]
  wire  _GEN_888; // @[Execute.scala 117:10]
  wire  _GEN_889; // @[Execute.scala 117:10]
  wire  _GEN_890; // @[Execute.scala 117:10]
  wire  _GEN_891; // @[Execute.scala 117:10]
  wire  _GEN_892; // @[Execute.scala 117:10]
  wire  _GEN_893; // @[Execute.scala 117:10]
  wire  _GEN_894; // @[Execute.scala 117:10]
  wire  _GEN_895; // @[Execute.scala 117:10]
  wire  _GEN_896; // @[Execute.scala 117:10]
  wire  _GEN_897; // @[Execute.scala 117:10]
  wire  _T_151; // @[Execute.scala 117:10]
  wire  _T_152; // @[Execute.scala 117:15]
  wire [5:0] _T_154; // @[Execute.scala 117:37]
  wire [5:0] _T_158; // @[Execute.scala 117:60]
  wire  _GEN_899; // @[Execute.scala 117:10]
  wire  _GEN_900; // @[Execute.scala 117:10]
  wire  _GEN_901; // @[Execute.scala 117:10]
  wire  _GEN_902; // @[Execute.scala 117:10]
  wire  _GEN_903; // @[Execute.scala 117:10]
  wire  _GEN_904; // @[Execute.scala 117:10]
  wire  _GEN_905; // @[Execute.scala 117:10]
  wire  _GEN_906; // @[Execute.scala 117:10]
  wire  _GEN_907; // @[Execute.scala 117:10]
  wire  _GEN_908; // @[Execute.scala 117:10]
  wire  _GEN_909; // @[Execute.scala 117:10]
  wire  _GEN_910; // @[Execute.scala 117:10]
  wire  _GEN_911; // @[Execute.scala 117:10]
  wire  _GEN_912; // @[Execute.scala 117:10]
  wire  _GEN_913; // @[Execute.scala 117:10]
  wire  _GEN_914; // @[Execute.scala 117:10]
  wire  _GEN_915; // @[Execute.scala 117:10]
  wire  _GEN_916; // @[Execute.scala 117:10]
  wire  _GEN_917; // @[Execute.scala 117:10]
  wire  _GEN_918; // @[Execute.scala 117:10]
  wire  _GEN_919; // @[Execute.scala 117:10]
  wire  _GEN_920; // @[Execute.scala 117:10]
  wire  _GEN_921; // @[Execute.scala 117:10]
  wire  _GEN_922; // @[Execute.scala 117:10]
  wire  _GEN_923; // @[Execute.scala 117:10]
  wire  _GEN_924; // @[Execute.scala 117:10]
  wire  _GEN_925; // @[Execute.scala 117:10]
  wire  _GEN_926; // @[Execute.scala 117:10]
  wire  _GEN_927; // @[Execute.scala 117:10]
  wire  _GEN_928; // @[Execute.scala 117:10]
  wire  _GEN_929; // @[Execute.scala 117:10]
  wire  _GEN_930; // @[Execute.scala 117:10]
  wire  _GEN_931; // @[Execute.scala 117:10]
  wire  _GEN_932; // @[Execute.scala 117:10]
  wire  _GEN_933; // @[Execute.scala 117:10]
  wire  _GEN_934; // @[Execute.scala 117:10]
  wire  _GEN_935; // @[Execute.scala 117:10]
  wire  _GEN_936; // @[Execute.scala 117:10]
  wire  _GEN_937; // @[Execute.scala 117:10]
  wire  _GEN_938; // @[Execute.scala 117:10]
  wire  _GEN_939; // @[Execute.scala 117:10]
  wire  _GEN_940; // @[Execute.scala 117:10]
  wire  _GEN_941; // @[Execute.scala 117:10]
  wire  _GEN_942; // @[Execute.scala 117:10]
  wire  _GEN_943; // @[Execute.scala 117:10]
  wire  _GEN_944; // @[Execute.scala 117:10]
  wire  _GEN_945; // @[Execute.scala 117:10]
  wire  _GEN_946; // @[Execute.scala 117:10]
  wire  _GEN_947; // @[Execute.scala 117:10]
  wire  _GEN_948; // @[Execute.scala 117:10]
  wire  _GEN_949; // @[Execute.scala 117:10]
  wire  _GEN_950; // @[Execute.scala 117:10]
  wire  _GEN_951; // @[Execute.scala 117:10]
  wire  _GEN_952; // @[Execute.scala 117:10]
  wire  _GEN_953; // @[Execute.scala 117:10]
  wire  _GEN_954; // @[Execute.scala 117:10]
  wire  _GEN_955; // @[Execute.scala 117:10]
  wire  _GEN_956; // @[Execute.scala 117:10]
  wire  _GEN_957; // @[Execute.scala 117:10]
  wire  _GEN_958; // @[Execute.scala 117:10]
  wire  _GEN_959; // @[Execute.scala 117:10]
  wire  _GEN_960; // @[Execute.scala 117:10]
  wire  _GEN_961; // @[Execute.scala 117:10]
  wire  _GEN_963; // @[Execute.scala 117:10]
  wire  _GEN_964; // @[Execute.scala 117:10]
  wire  _GEN_965; // @[Execute.scala 117:10]
  wire  _GEN_966; // @[Execute.scala 117:10]
  wire  _GEN_967; // @[Execute.scala 117:10]
  wire  _GEN_968; // @[Execute.scala 117:10]
  wire  _GEN_969; // @[Execute.scala 117:10]
  wire  _GEN_970; // @[Execute.scala 117:10]
  wire  _GEN_971; // @[Execute.scala 117:10]
  wire  _GEN_972; // @[Execute.scala 117:10]
  wire  _GEN_973; // @[Execute.scala 117:10]
  wire  _GEN_974; // @[Execute.scala 117:10]
  wire  _GEN_975; // @[Execute.scala 117:10]
  wire  _GEN_976; // @[Execute.scala 117:10]
  wire  _GEN_977; // @[Execute.scala 117:10]
  wire  _GEN_978; // @[Execute.scala 117:10]
  wire  _GEN_979; // @[Execute.scala 117:10]
  wire  _GEN_980; // @[Execute.scala 117:10]
  wire  _GEN_981; // @[Execute.scala 117:10]
  wire  _GEN_982; // @[Execute.scala 117:10]
  wire  _GEN_983; // @[Execute.scala 117:10]
  wire  _GEN_984; // @[Execute.scala 117:10]
  wire  _GEN_985; // @[Execute.scala 117:10]
  wire  _GEN_986; // @[Execute.scala 117:10]
  wire  _GEN_987; // @[Execute.scala 117:10]
  wire  _GEN_988; // @[Execute.scala 117:10]
  wire  _GEN_989; // @[Execute.scala 117:10]
  wire  _GEN_990; // @[Execute.scala 117:10]
  wire  _GEN_991; // @[Execute.scala 117:10]
  wire  _GEN_992; // @[Execute.scala 117:10]
  wire  _GEN_993; // @[Execute.scala 117:10]
  wire  _GEN_994; // @[Execute.scala 117:10]
  wire  _GEN_995; // @[Execute.scala 117:10]
  wire  _GEN_996; // @[Execute.scala 117:10]
  wire  _GEN_997; // @[Execute.scala 117:10]
  wire  _GEN_998; // @[Execute.scala 117:10]
  wire  _GEN_999; // @[Execute.scala 117:10]
  wire  _GEN_1000; // @[Execute.scala 117:10]
  wire  _GEN_1001; // @[Execute.scala 117:10]
  wire  _GEN_1002; // @[Execute.scala 117:10]
  wire  _GEN_1003; // @[Execute.scala 117:10]
  wire  _GEN_1004; // @[Execute.scala 117:10]
  wire  _GEN_1005; // @[Execute.scala 117:10]
  wire  _GEN_1006; // @[Execute.scala 117:10]
  wire  _GEN_1007; // @[Execute.scala 117:10]
  wire  _GEN_1008; // @[Execute.scala 117:10]
  wire  _GEN_1009; // @[Execute.scala 117:10]
  wire  _GEN_1010; // @[Execute.scala 117:10]
  wire  _GEN_1011; // @[Execute.scala 117:10]
  wire  _GEN_1012; // @[Execute.scala 117:10]
  wire  _GEN_1013; // @[Execute.scala 117:10]
  wire  _GEN_1014; // @[Execute.scala 117:10]
  wire  _GEN_1015; // @[Execute.scala 117:10]
  wire  _GEN_1016; // @[Execute.scala 117:10]
  wire  _GEN_1017; // @[Execute.scala 117:10]
  wire  _GEN_1018; // @[Execute.scala 117:10]
  wire  _GEN_1019; // @[Execute.scala 117:10]
  wire  _GEN_1020; // @[Execute.scala 117:10]
  wire  _GEN_1021; // @[Execute.scala 117:10]
  wire  _GEN_1022; // @[Execute.scala 117:10]
  wire  _GEN_1023; // @[Execute.scala 117:10]
  wire  _GEN_1024; // @[Execute.scala 117:10]
  wire  _GEN_1025; // @[Execute.scala 117:10]
  wire  _T_161; // @[Execute.scala 117:10]
  wire  _T_162; // @[Execute.scala 117:15]
  wire [5:0] _T_164; // @[Execute.scala 117:37]
  wire [5:0] _T_168; // @[Execute.scala 117:60]
  wire  _GEN_1027; // @[Execute.scala 117:10]
  wire  _GEN_1028; // @[Execute.scala 117:10]
  wire  _GEN_1029; // @[Execute.scala 117:10]
  wire  _GEN_1030; // @[Execute.scala 117:10]
  wire  _GEN_1031; // @[Execute.scala 117:10]
  wire  _GEN_1032; // @[Execute.scala 117:10]
  wire  _GEN_1033; // @[Execute.scala 117:10]
  wire  _GEN_1034; // @[Execute.scala 117:10]
  wire  _GEN_1035; // @[Execute.scala 117:10]
  wire  _GEN_1036; // @[Execute.scala 117:10]
  wire  _GEN_1037; // @[Execute.scala 117:10]
  wire  _GEN_1038; // @[Execute.scala 117:10]
  wire  _GEN_1039; // @[Execute.scala 117:10]
  wire  _GEN_1040; // @[Execute.scala 117:10]
  wire  _GEN_1041; // @[Execute.scala 117:10]
  wire  _GEN_1042; // @[Execute.scala 117:10]
  wire  _GEN_1043; // @[Execute.scala 117:10]
  wire  _GEN_1044; // @[Execute.scala 117:10]
  wire  _GEN_1045; // @[Execute.scala 117:10]
  wire  _GEN_1046; // @[Execute.scala 117:10]
  wire  _GEN_1047; // @[Execute.scala 117:10]
  wire  _GEN_1048; // @[Execute.scala 117:10]
  wire  _GEN_1049; // @[Execute.scala 117:10]
  wire  _GEN_1050; // @[Execute.scala 117:10]
  wire  _GEN_1051; // @[Execute.scala 117:10]
  wire  _GEN_1052; // @[Execute.scala 117:10]
  wire  _GEN_1053; // @[Execute.scala 117:10]
  wire  _GEN_1054; // @[Execute.scala 117:10]
  wire  _GEN_1055; // @[Execute.scala 117:10]
  wire  _GEN_1056; // @[Execute.scala 117:10]
  wire  _GEN_1057; // @[Execute.scala 117:10]
  wire  _GEN_1058; // @[Execute.scala 117:10]
  wire  _GEN_1059; // @[Execute.scala 117:10]
  wire  _GEN_1060; // @[Execute.scala 117:10]
  wire  _GEN_1061; // @[Execute.scala 117:10]
  wire  _GEN_1062; // @[Execute.scala 117:10]
  wire  _GEN_1063; // @[Execute.scala 117:10]
  wire  _GEN_1064; // @[Execute.scala 117:10]
  wire  _GEN_1065; // @[Execute.scala 117:10]
  wire  _GEN_1066; // @[Execute.scala 117:10]
  wire  _GEN_1067; // @[Execute.scala 117:10]
  wire  _GEN_1068; // @[Execute.scala 117:10]
  wire  _GEN_1069; // @[Execute.scala 117:10]
  wire  _GEN_1070; // @[Execute.scala 117:10]
  wire  _GEN_1071; // @[Execute.scala 117:10]
  wire  _GEN_1072; // @[Execute.scala 117:10]
  wire  _GEN_1073; // @[Execute.scala 117:10]
  wire  _GEN_1074; // @[Execute.scala 117:10]
  wire  _GEN_1075; // @[Execute.scala 117:10]
  wire  _GEN_1076; // @[Execute.scala 117:10]
  wire  _GEN_1077; // @[Execute.scala 117:10]
  wire  _GEN_1078; // @[Execute.scala 117:10]
  wire  _GEN_1079; // @[Execute.scala 117:10]
  wire  _GEN_1080; // @[Execute.scala 117:10]
  wire  _GEN_1081; // @[Execute.scala 117:10]
  wire  _GEN_1082; // @[Execute.scala 117:10]
  wire  _GEN_1083; // @[Execute.scala 117:10]
  wire  _GEN_1084; // @[Execute.scala 117:10]
  wire  _GEN_1085; // @[Execute.scala 117:10]
  wire  _GEN_1086; // @[Execute.scala 117:10]
  wire  _GEN_1087; // @[Execute.scala 117:10]
  wire  _GEN_1088; // @[Execute.scala 117:10]
  wire  _GEN_1089; // @[Execute.scala 117:10]
  wire  _GEN_1091; // @[Execute.scala 117:10]
  wire  _GEN_1092; // @[Execute.scala 117:10]
  wire  _GEN_1093; // @[Execute.scala 117:10]
  wire  _GEN_1094; // @[Execute.scala 117:10]
  wire  _GEN_1095; // @[Execute.scala 117:10]
  wire  _GEN_1096; // @[Execute.scala 117:10]
  wire  _GEN_1097; // @[Execute.scala 117:10]
  wire  _GEN_1098; // @[Execute.scala 117:10]
  wire  _GEN_1099; // @[Execute.scala 117:10]
  wire  _GEN_1100; // @[Execute.scala 117:10]
  wire  _GEN_1101; // @[Execute.scala 117:10]
  wire  _GEN_1102; // @[Execute.scala 117:10]
  wire  _GEN_1103; // @[Execute.scala 117:10]
  wire  _GEN_1104; // @[Execute.scala 117:10]
  wire  _GEN_1105; // @[Execute.scala 117:10]
  wire  _GEN_1106; // @[Execute.scala 117:10]
  wire  _GEN_1107; // @[Execute.scala 117:10]
  wire  _GEN_1108; // @[Execute.scala 117:10]
  wire  _GEN_1109; // @[Execute.scala 117:10]
  wire  _GEN_1110; // @[Execute.scala 117:10]
  wire  _GEN_1111; // @[Execute.scala 117:10]
  wire  _GEN_1112; // @[Execute.scala 117:10]
  wire  _GEN_1113; // @[Execute.scala 117:10]
  wire  _GEN_1114; // @[Execute.scala 117:10]
  wire  _GEN_1115; // @[Execute.scala 117:10]
  wire  _GEN_1116; // @[Execute.scala 117:10]
  wire  _GEN_1117; // @[Execute.scala 117:10]
  wire  _GEN_1118; // @[Execute.scala 117:10]
  wire  _GEN_1119; // @[Execute.scala 117:10]
  wire  _GEN_1120; // @[Execute.scala 117:10]
  wire  _GEN_1121; // @[Execute.scala 117:10]
  wire  _GEN_1122; // @[Execute.scala 117:10]
  wire  _GEN_1123; // @[Execute.scala 117:10]
  wire  _GEN_1124; // @[Execute.scala 117:10]
  wire  _GEN_1125; // @[Execute.scala 117:10]
  wire  _GEN_1126; // @[Execute.scala 117:10]
  wire  _GEN_1127; // @[Execute.scala 117:10]
  wire  _GEN_1128; // @[Execute.scala 117:10]
  wire  _GEN_1129; // @[Execute.scala 117:10]
  wire  _GEN_1130; // @[Execute.scala 117:10]
  wire  _GEN_1131; // @[Execute.scala 117:10]
  wire  _GEN_1132; // @[Execute.scala 117:10]
  wire  _GEN_1133; // @[Execute.scala 117:10]
  wire  _GEN_1134; // @[Execute.scala 117:10]
  wire  _GEN_1135; // @[Execute.scala 117:10]
  wire  _GEN_1136; // @[Execute.scala 117:10]
  wire  _GEN_1137; // @[Execute.scala 117:10]
  wire  _GEN_1138; // @[Execute.scala 117:10]
  wire  _GEN_1139; // @[Execute.scala 117:10]
  wire  _GEN_1140; // @[Execute.scala 117:10]
  wire  _GEN_1141; // @[Execute.scala 117:10]
  wire  _GEN_1142; // @[Execute.scala 117:10]
  wire  _GEN_1143; // @[Execute.scala 117:10]
  wire  _GEN_1144; // @[Execute.scala 117:10]
  wire  _GEN_1145; // @[Execute.scala 117:10]
  wire  _GEN_1146; // @[Execute.scala 117:10]
  wire  _GEN_1147; // @[Execute.scala 117:10]
  wire  _GEN_1148; // @[Execute.scala 117:10]
  wire  _GEN_1149; // @[Execute.scala 117:10]
  wire  _GEN_1150; // @[Execute.scala 117:10]
  wire  _GEN_1151; // @[Execute.scala 117:10]
  wire  _GEN_1152; // @[Execute.scala 117:10]
  wire  _GEN_1153; // @[Execute.scala 117:10]
  wire  _T_171; // @[Execute.scala 117:10]
  wire  _T_172; // @[Execute.scala 117:15]
  wire [5:0] _T_174; // @[Execute.scala 117:37]
  wire [5:0] _T_178; // @[Execute.scala 117:60]
  wire  _GEN_1155; // @[Execute.scala 117:10]
  wire  _GEN_1156; // @[Execute.scala 117:10]
  wire  _GEN_1157; // @[Execute.scala 117:10]
  wire  _GEN_1158; // @[Execute.scala 117:10]
  wire  _GEN_1159; // @[Execute.scala 117:10]
  wire  _GEN_1160; // @[Execute.scala 117:10]
  wire  _GEN_1161; // @[Execute.scala 117:10]
  wire  _GEN_1162; // @[Execute.scala 117:10]
  wire  _GEN_1163; // @[Execute.scala 117:10]
  wire  _GEN_1164; // @[Execute.scala 117:10]
  wire  _GEN_1165; // @[Execute.scala 117:10]
  wire  _GEN_1166; // @[Execute.scala 117:10]
  wire  _GEN_1167; // @[Execute.scala 117:10]
  wire  _GEN_1168; // @[Execute.scala 117:10]
  wire  _GEN_1169; // @[Execute.scala 117:10]
  wire  _GEN_1170; // @[Execute.scala 117:10]
  wire  _GEN_1171; // @[Execute.scala 117:10]
  wire  _GEN_1172; // @[Execute.scala 117:10]
  wire  _GEN_1173; // @[Execute.scala 117:10]
  wire  _GEN_1174; // @[Execute.scala 117:10]
  wire  _GEN_1175; // @[Execute.scala 117:10]
  wire  _GEN_1176; // @[Execute.scala 117:10]
  wire  _GEN_1177; // @[Execute.scala 117:10]
  wire  _GEN_1178; // @[Execute.scala 117:10]
  wire  _GEN_1179; // @[Execute.scala 117:10]
  wire  _GEN_1180; // @[Execute.scala 117:10]
  wire  _GEN_1181; // @[Execute.scala 117:10]
  wire  _GEN_1182; // @[Execute.scala 117:10]
  wire  _GEN_1183; // @[Execute.scala 117:10]
  wire  _GEN_1184; // @[Execute.scala 117:10]
  wire  _GEN_1185; // @[Execute.scala 117:10]
  wire  _GEN_1186; // @[Execute.scala 117:10]
  wire  _GEN_1187; // @[Execute.scala 117:10]
  wire  _GEN_1188; // @[Execute.scala 117:10]
  wire  _GEN_1189; // @[Execute.scala 117:10]
  wire  _GEN_1190; // @[Execute.scala 117:10]
  wire  _GEN_1191; // @[Execute.scala 117:10]
  wire  _GEN_1192; // @[Execute.scala 117:10]
  wire  _GEN_1193; // @[Execute.scala 117:10]
  wire  _GEN_1194; // @[Execute.scala 117:10]
  wire  _GEN_1195; // @[Execute.scala 117:10]
  wire  _GEN_1196; // @[Execute.scala 117:10]
  wire  _GEN_1197; // @[Execute.scala 117:10]
  wire  _GEN_1198; // @[Execute.scala 117:10]
  wire  _GEN_1199; // @[Execute.scala 117:10]
  wire  _GEN_1200; // @[Execute.scala 117:10]
  wire  _GEN_1201; // @[Execute.scala 117:10]
  wire  _GEN_1202; // @[Execute.scala 117:10]
  wire  _GEN_1203; // @[Execute.scala 117:10]
  wire  _GEN_1204; // @[Execute.scala 117:10]
  wire  _GEN_1205; // @[Execute.scala 117:10]
  wire  _GEN_1206; // @[Execute.scala 117:10]
  wire  _GEN_1207; // @[Execute.scala 117:10]
  wire  _GEN_1208; // @[Execute.scala 117:10]
  wire  _GEN_1209; // @[Execute.scala 117:10]
  wire  _GEN_1210; // @[Execute.scala 117:10]
  wire  _GEN_1211; // @[Execute.scala 117:10]
  wire  _GEN_1212; // @[Execute.scala 117:10]
  wire  _GEN_1213; // @[Execute.scala 117:10]
  wire  _GEN_1214; // @[Execute.scala 117:10]
  wire  _GEN_1215; // @[Execute.scala 117:10]
  wire  _GEN_1216; // @[Execute.scala 117:10]
  wire  _GEN_1217; // @[Execute.scala 117:10]
  wire  _GEN_1219; // @[Execute.scala 117:10]
  wire  _GEN_1220; // @[Execute.scala 117:10]
  wire  _GEN_1221; // @[Execute.scala 117:10]
  wire  _GEN_1222; // @[Execute.scala 117:10]
  wire  _GEN_1223; // @[Execute.scala 117:10]
  wire  _GEN_1224; // @[Execute.scala 117:10]
  wire  _GEN_1225; // @[Execute.scala 117:10]
  wire  _GEN_1226; // @[Execute.scala 117:10]
  wire  _GEN_1227; // @[Execute.scala 117:10]
  wire  _GEN_1228; // @[Execute.scala 117:10]
  wire  _GEN_1229; // @[Execute.scala 117:10]
  wire  _GEN_1230; // @[Execute.scala 117:10]
  wire  _GEN_1231; // @[Execute.scala 117:10]
  wire  _GEN_1232; // @[Execute.scala 117:10]
  wire  _GEN_1233; // @[Execute.scala 117:10]
  wire  _GEN_1234; // @[Execute.scala 117:10]
  wire  _GEN_1235; // @[Execute.scala 117:10]
  wire  _GEN_1236; // @[Execute.scala 117:10]
  wire  _GEN_1237; // @[Execute.scala 117:10]
  wire  _GEN_1238; // @[Execute.scala 117:10]
  wire  _GEN_1239; // @[Execute.scala 117:10]
  wire  _GEN_1240; // @[Execute.scala 117:10]
  wire  _GEN_1241; // @[Execute.scala 117:10]
  wire  _GEN_1242; // @[Execute.scala 117:10]
  wire  _GEN_1243; // @[Execute.scala 117:10]
  wire  _GEN_1244; // @[Execute.scala 117:10]
  wire  _GEN_1245; // @[Execute.scala 117:10]
  wire  _GEN_1246; // @[Execute.scala 117:10]
  wire  _GEN_1247; // @[Execute.scala 117:10]
  wire  _GEN_1248; // @[Execute.scala 117:10]
  wire  _GEN_1249; // @[Execute.scala 117:10]
  wire  _GEN_1250; // @[Execute.scala 117:10]
  wire  _GEN_1251; // @[Execute.scala 117:10]
  wire  _GEN_1252; // @[Execute.scala 117:10]
  wire  _GEN_1253; // @[Execute.scala 117:10]
  wire  _GEN_1254; // @[Execute.scala 117:10]
  wire  _GEN_1255; // @[Execute.scala 117:10]
  wire  _GEN_1256; // @[Execute.scala 117:10]
  wire  _GEN_1257; // @[Execute.scala 117:10]
  wire  _GEN_1258; // @[Execute.scala 117:10]
  wire  _GEN_1259; // @[Execute.scala 117:10]
  wire  _GEN_1260; // @[Execute.scala 117:10]
  wire  _GEN_1261; // @[Execute.scala 117:10]
  wire  _GEN_1262; // @[Execute.scala 117:10]
  wire  _GEN_1263; // @[Execute.scala 117:10]
  wire  _GEN_1264; // @[Execute.scala 117:10]
  wire  _GEN_1265; // @[Execute.scala 117:10]
  wire  _GEN_1266; // @[Execute.scala 117:10]
  wire  _GEN_1267; // @[Execute.scala 117:10]
  wire  _GEN_1268; // @[Execute.scala 117:10]
  wire  _GEN_1269; // @[Execute.scala 117:10]
  wire  _GEN_1270; // @[Execute.scala 117:10]
  wire  _GEN_1271; // @[Execute.scala 117:10]
  wire  _GEN_1272; // @[Execute.scala 117:10]
  wire  _GEN_1273; // @[Execute.scala 117:10]
  wire  _GEN_1274; // @[Execute.scala 117:10]
  wire  _GEN_1275; // @[Execute.scala 117:10]
  wire  _GEN_1276; // @[Execute.scala 117:10]
  wire  _GEN_1277; // @[Execute.scala 117:10]
  wire  _GEN_1278; // @[Execute.scala 117:10]
  wire  _GEN_1279; // @[Execute.scala 117:10]
  wire  _GEN_1280; // @[Execute.scala 117:10]
  wire  _GEN_1281; // @[Execute.scala 117:10]
  wire  _T_181; // @[Execute.scala 117:10]
  wire  _T_182; // @[Execute.scala 117:15]
  wire [5:0] _T_184; // @[Execute.scala 117:37]
  wire [5:0] _T_188; // @[Execute.scala 117:60]
  wire  _GEN_1283; // @[Execute.scala 117:10]
  wire  _GEN_1284; // @[Execute.scala 117:10]
  wire  _GEN_1285; // @[Execute.scala 117:10]
  wire  _GEN_1286; // @[Execute.scala 117:10]
  wire  _GEN_1287; // @[Execute.scala 117:10]
  wire  _GEN_1288; // @[Execute.scala 117:10]
  wire  _GEN_1289; // @[Execute.scala 117:10]
  wire  _GEN_1290; // @[Execute.scala 117:10]
  wire  _GEN_1291; // @[Execute.scala 117:10]
  wire  _GEN_1292; // @[Execute.scala 117:10]
  wire  _GEN_1293; // @[Execute.scala 117:10]
  wire  _GEN_1294; // @[Execute.scala 117:10]
  wire  _GEN_1295; // @[Execute.scala 117:10]
  wire  _GEN_1296; // @[Execute.scala 117:10]
  wire  _GEN_1297; // @[Execute.scala 117:10]
  wire  _GEN_1298; // @[Execute.scala 117:10]
  wire  _GEN_1299; // @[Execute.scala 117:10]
  wire  _GEN_1300; // @[Execute.scala 117:10]
  wire  _GEN_1301; // @[Execute.scala 117:10]
  wire  _GEN_1302; // @[Execute.scala 117:10]
  wire  _GEN_1303; // @[Execute.scala 117:10]
  wire  _GEN_1304; // @[Execute.scala 117:10]
  wire  _GEN_1305; // @[Execute.scala 117:10]
  wire  _GEN_1306; // @[Execute.scala 117:10]
  wire  _GEN_1307; // @[Execute.scala 117:10]
  wire  _GEN_1308; // @[Execute.scala 117:10]
  wire  _GEN_1309; // @[Execute.scala 117:10]
  wire  _GEN_1310; // @[Execute.scala 117:10]
  wire  _GEN_1311; // @[Execute.scala 117:10]
  wire  _GEN_1312; // @[Execute.scala 117:10]
  wire  _GEN_1313; // @[Execute.scala 117:10]
  wire  _GEN_1314; // @[Execute.scala 117:10]
  wire  _GEN_1315; // @[Execute.scala 117:10]
  wire  _GEN_1316; // @[Execute.scala 117:10]
  wire  _GEN_1317; // @[Execute.scala 117:10]
  wire  _GEN_1318; // @[Execute.scala 117:10]
  wire  _GEN_1319; // @[Execute.scala 117:10]
  wire  _GEN_1320; // @[Execute.scala 117:10]
  wire  _GEN_1321; // @[Execute.scala 117:10]
  wire  _GEN_1322; // @[Execute.scala 117:10]
  wire  _GEN_1323; // @[Execute.scala 117:10]
  wire  _GEN_1324; // @[Execute.scala 117:10]
  wire  _GEN_1325; // @[Execute.scala 117:10]
  wire  _GEN_1326; // @[Execute.scala 117:10]
  wire  _GEN_1327; // @[Execute.scala 117:10]
  wire  _GEN_1328; // @[Execute.scala 117:10]
  wire  _GEN_1329; // @[Execute.scala 117:10]
  wire  _GEN_1330; // @[Execute.scala 117:10]
  wire  _GEN_1331; // @[Execute.scala 117:10]
  wire  _GEN_1332; // @[Execute.scala 117:10]
  wire  _GEN_1333; // @[Execute.scala 117:10]
  wire  _GEN_1334; // @[Execute.scala 117:10]
  wire  _GEN_1335; // @[Execute.scala 117:10]
  wire  _GEN_1336; // @[Execute.scala 117:10]
  wire  _GEN_1337; // @[Execute.scala 117:10]
  wire  _GEN_1338; // @[Execute.scala 117:10]
  wire  _GEN_1339; // @[Execute.scala 117:10]
  wire  _GEN_1340; // @[Execute.scala 117:10]
  wire  _GEN_1341; // @[Execute.scala 117:10]
  wire  _GEN_1342; // @[Execute.scala 117:10]
  wire  _GEN_1343; // @[Execute.scala 117:10]
  wire  _GEN_1344; // @[Execute.scala 117:10]
  wire  _GEN_1345; // @[Execute.scala 117:10]
  wire  _GEN_1347; // @[Execute.scala 117:10]
  wire  _GEN_1348; // @[Execute.scala 117:10]
  wire  _GEN_1349; // @[Execute.scala 117:10]
  wire  _GEN_1350; // @[Execute.scala 117:10]
  wire  _GEN_1351; // @[Execute.scala 117:10]
  wire  _GEN_1352; // @[Execute.scala 117:10]
  wire  _GEN_1353; // @[Execute.scala 117:10]
  wire  _GEN_1354; // @[Execute.scala 117:10]
  wire  _GEN_1355; // @[Execute.scala 117:10]
  wire  _GEN_1356; // @[Execute.scala 117:10]
  wire  _GEN_1357; // @[Execute.scala 117:10]
  wire  _GEN_1358; // @[Execute.scala 117:10]
  wire  _GEN_1359; // @[Execute.scala 117:10]
  wire  _GEN_1360; // @[Execute.scala 117:10]
  wire  _GEN_1361; // @[Execute.scala 117:10]
  wire  _GEN_1362; // @[Execute.scala 117:10]
  wire  _GEN_1363; // @[Execute.scala 117:10]
  wire  _GEN_1364; // @[Execute.scala 117:10]
  wire  _GEN_1365; // @[Execute.scala 117:10]
  wire  _GEN_1366; // @[Execute.scala 117:10]
  wire  _GEN_1367; // @[Execute.scala 117:10]
  wire  _GEN_1368; // @[Execute.scala 117:10]
  wire  _GEN_1369; // @[Execute.scala 117:10]
  wire  _GEN_1370; // @[Execute.scala 117:10]
  wire  _GEN_1371; // @[Execute.scala 117:10]
  wire  _GEN_1372; // @[Execute.scala 117:10]
  wire  _GEN_1373; // @[Execute.scala 117:10]
  wire  _GEN_1374; // @[Execute.scala 117:10]
  wire  _GEN_1375; // @[Execute.scala 117:10]
  wire  _GEN_1376; // @[Execute.scala 117:10]
  wire  _GEN_1377; // @[Execute.scala 117:10]
  wire  _GEN_1378; // @[Execute.scala 117:10]
  wire  _GEN_1379; // @[Execute.scala 117:10]
  wire  _GEN_1380; // @[Execute.scala 117:10]
  wire  _GEN_1381; // @[Execute.scala 117:10]
  wire  _GEN_1382; // @[Execute.scala 117:10]
  wire  _GEN_1383; // @[Execute.scala 117:10]
  wire  _GEN_1384; // @[Execute.scala 117:10]
  wire  _GEN_1385; // @[Execute.scala 117:10]
  wire  _GEN_1386; // @[Execute.scala 117:10]
  wire  _GEN_1387; // @[Execute.scala 117:10]
  wire  _GEN_1388; // @[Execute.scala 117:10]
  wire  _GEN_1389; // @[Execute.scala 117:10]
  wire  _GEN_1390; // @[Execute.scala 117:10]
  wire  _GEN_1391; // @[Execute.scala 117:10]
  wire  _GEN_1392; // @[Execute.scala 117:10]
  wire  _GEN_1393; // @[Execute.scala 117:10]
  wire  _GEN_1394; // @[Execute.scala 117:10]
  wire  _GEN_1395; // @[Execute.scala 117:10]
  wire  _GEN_1396; // @[Execute.scala 117:10]
  wire  _GEN_1397; // @[Execute.scala 117:10]
  wire  _GEN_1398; // @[Execute.scala 117:10]
  wire  _GEN_1399; // @[Execute.scala 117:10]
  wire  _GEN_1400; // @[Execute.scala 117:10]
  wire  _GEN_1401; // @[Execute.scala 117:10]
  wire  _GEN_1402; // @[Execute.scala 117:10]
  wire  _GEN_1403; // @[Execute.scala 117:10]
  wire  _GEN_1404; // @[Execute.scala 117:10]
  wire  _GEN_1405; // @[Execute.scala 117:10]
  wire  _GEN_1406; // @[Execute.scala 117:10]
  wire  _GEN_1407; // @[Execute.scala 117:10]
  wire  _GEN_1408; // @[Execute.scala 117:10]
  wire  _GEN_1409; // @[Execute.scala 117:10]
  wire  _T_191; // @[Execute.scala 117:10]
  wire  _T_192; // @[Execute.scala 117:15]
  wire [5:0] _T_194; // @[Execute.scala 117:37]
  wire [5:0] _T_198; // @[Execute.scala 117:60]
  wire  _GEN_1411; // @[Execute.scala 117:10]
  wire  _GEN_1412; // @[Execute.scala 117:10]
  wire  _GEN_1413; // @[Execute.scala 117:10]
  wire  _GEN_1414; // @[Execute.scala 117:10]
  wire  _GEN_1415; // @[Execute.scala 117:10]
  wire  _GEN_1416; // @[Execute.scala 117:10]
  wire  _GEN_1417; // @[Execute.scala 117:10]
  wire  _GEN_1418; // @[Execute.scala 117:10]
  wire  _GEN_1419; // @[Execute.scala 117:10]
  wire  _GEN_1420; // @[Execute.scala 117:10]
  wire  _GEN_1421; // @[Execute.scala 117:10]
  wire  _GEN_1422; // @[Execute.scala 117:10]
  wire  _GEN_1423; // @[Execute.scala 117:10]
  wire  _GEN_1424; // @[Execute.scala 117:10]
  wire  _GEN_1425; // @[Execute.scala 117:10]
  wire  _GEN_1426; // @[Execute.scala 117:10]
  wire  _GEN_1427; // @[Execute.scala 117:10]
  wire  _GEN_1428; // @[Execute.scala 117:10]
  wire  _GEN_1429; // @[Execute.scala 117:10]
  wire  _GEN_1430; // @[Execute.scala 117:10]
  wire  _GEN_1431; // @[Execute.scala 117:10]
  wire  _GEN_1432; // @[Execute.scala 117:10]
  wire  _GEN_1433; // @[Execute.scala 117:10]
  wire  _GEN_1434; // @[Execute.scala 117:10]
  wire  _GEN_1435; // @[Execute.scala 117:10]
  wire  _GEN_1436; // @[Execute.scala 117:10]
  wire  _GEN_1437; // @[Execute.scala 117:10]
  wire  _GEN_1438; // @[Execute.scala 117:10]
  wire  _GEN_1439; // @[Execute.scala 117:10]
  wire  _GEN_1440; // @[Execute.scala 117:10]
  wire  _GEN_1441; // @[Execute.scala 117:10]
  wire  _GEN_1442; // @[Execute.scala 117:10]
  wire  _GEN_1443; // @[Execute.scala 117:10]
  wire  _GEN_1444; // @[Execute.scala 117:10]
  wire  _GEN_1445; // @[Execute.scala 117:10]
  wire  _GEN_1446; // @[Execute.scala 117:10]
  wire  _GEN_1447; // @[Execute.scala 117:10]
  wire  _GEN_1448; // @[Execute.scala 117:10]
  wire  _GEN_1449; // @[Execute.scala 117:10]
  wire  _GEN_1450; // @[Execute.scala 117:10]
  wire  _GEN_1451; // @[Execute.scala 117:10]
  wire  _GEN_1452; // @[Execute.scala 117:10]
  wire  _GEN_1453; // @[Execute.scala 117:10]
  wire  _GEN_1454; // @[Execute.scala 117:10]
  wire  _GEN_1455; // @[Execute.scala 117:10]
  wire  _GEN_1456; // @[Execute.scala 117:10]
  wire  _GEN_1457; // @[Execute.scala 117:10]
  wire  _GEN_1458; // @[Execute.scala 117:10]
  wire  _GEN_1459; // @[Execute.scala 117:10]
  wire  _GEN_1460; // @[Execute.scala 117:10]
  wire  _GEN_1461; // @[Execute.scala 117:10]
  wire  _GEN_1462; // @[Execute.scala 117:10]
  wire  _GEN_1463; // @[Execute.scala 117:10]
  wire  _GEN_1464; // @[Execute.scala 117:10]
  wire  _GEN_1465; // @[Execute.scala 117:10]
  wire  _GEN_1466; // @[Execute.scala 117:10]
  wire  _GEN_1467; // @[Execute.scala 117:10]
  wire  _GEN_1468; // @[Execute.scala 117:10]
  wire  _GEN_1469; // @[Execute.scala 117:10]
  wire  _GEN_1470; // @[Execute.scala 117:10]
  wire  _GEN_1471; // @[Execute.scala 117:10]
  wire  _GEN_1472; // @[Execute.scala 117:10]
  wire  _GEN_1473; // @[Execute.scala 117:10]
  wire  _GEN_1475; // @[Execute.scala 117:10]
  wire  _GEN_1476; // @[Execute.scala 117:10]
  wire  _GEN_1477; // @[Execute.scala 117:10]
  wire  _GEN_1478; // @[Execute.scala 117:10]
  wire  _GEN_1479; // @[Execute.scala 117:10]
  wire  _GEN_1480; // @[Execute.scala 117:10]
  wire  _GEN_1481; // @[Execute.scala 117:10]
  wire  _GEN_1482; // @[Execute.scala 117:10]
  wire  _GEN_1483; // @[Execute.scala 117:10]
  wire  _GEN_1484; // @[Execute.scala 117:10]
  wire  _GEN_1485; // @[Execute.scala 117:10]
  wire  _GEN_1486; // @[Execute.scala 117:10]
  wire  _GEN_1487; // @[Execute.scala 117:10]
  wire  _GEN_1488; // @[Execute.scala 117:10]
  wire  _GEN_1489; // @[Execute.scala 117:10]
  wire  _GEN_1490; // @[Execute.scala 117:10]
  wire  _GEN_1491; // @[Execute.scala 117:10]
  wire  _GEN_1492; // @[Execute.scala 117:10]
  wire  _GEN_1493; // @[Execute.scala 117:10]
  wire  _GEN_1494; // @[Execute.scala 117:10]
  wire  _GEN_1495; // @[Execute.scala 117:10]
  wire  _GEN_1496; // @[Execute.scala 117:10]
  wire  _GEN_1497; // @[Execute.scala 117:10]
  wire  _GEN_1498; // @[Execute.scala 117:10]
  wire  _GEN_1499; // @[Execute.scala 117:10]
  wire  _GEN_1500; // @[Execute.scala 117:10]
  wire  _GEN_1501; // @[Execute.scala 117:10]
  wire  _GEN_1502; // @[Execute.scala 117:10]
  wire  _GEN_1503; // @[Execute.scala 117:10]
  wire  _GEN_1504; // @[Execute.scala 117:10]
  wire  _GEN_1505; // @[Execute.scala 117:10]
  wire  _GEN_1506; // @[Execute.scala 117:10]
  wire  _GEN_1507; // @[Execute.scala 117:10]
  wire  _GEN_1508; // @[Execute.scala 117:10]
  wire  _GEN_1509; // @[Execute.scala 117:10]
  wire  _GEN_1510; // @[Execute.scala 117:10]
  wire  _GEN_1511; // @[Execute.scala 117:10]
  wire  _GEN_1512; // @[Execute.scala 117:10]
  wire  _GEN_1513; // @[Execute.scala 117:10]
  wire  _GEN_1514; // @[Execute.scala 117:10]
  wire  _GEN_1515; // @[Execute.scala 117:10]
  wire  _GEN_1516; // @[Execute.scala 117:10]
  wire  _GEN_1517; // @[Execute.scala 117:10]
  wire  _GEN_1518; // @[Execute.scala 117:10]
  wire  _GEN_1519; // @[Execute.scala 117:10]
  wire  _GEN_1520; // @[Execute.scala 117:10]
  wire  _GEN_1521; // @[Execute.scala 117:10]
  wire  _GEN_1522; // @[Execute.scala 117:10]
  wire  _GEN_1523; // @[Execute.scala 117:10]
  wire  _GEN_1524; // @[Execute.scala 117:10]
  wire  _GEN_1525; // @[Execute.scala 117:10]
  wire  _GEN_1526; // @[Execute.scala 117:10]
  wire  _GEN_1527; // @[Execute.scala 117:10]
  wire  _GEN_1528; // @[Execute.scala 117:10]
  wire  _GEN_1529; // @[Execute.scala 117:10]
  wire  _GEN_1530; // @[Execute.scala 117:10]
  wire  _GEN_1531; // @[Execute.scala 117:10]
  wire  _GEN_1532; // @[Execute.scala 117:10]
  wire  _GEN_1533; // @[Execute.scala 117:10]
  wire  _GEN_1534; // @[Execute.scala 117:10]
  wire  _GEN_1535; // @[Execute.scala 117:10]
  wire  _GEN_1536; // @[Execute.scala 117:10]
  wire  _GEN_1537; // @[Execute.scala 117:10]
  wire  _T_201; // @[Execute.scala 117:10]
  wire  _T_202; // @[Execute.scala 117:15]
  wire [5:0] _T_204; // @[Execute.scala 117:37]
  wire [5:0] _T_208; // @[Execute.scala 117:60]
  wire  _GEN_1539; // @[Execute.scala 117:10]
  wire  _GEN_1540; // @[Execute.scala 117:10]
  wire  _GEN_1541; // @[Execute.scala 117:10]
  wire  _GEN_1542; // @[Execute.scala 117:10]
  wire  _GEN_1543; // @[Execute.scala 117:10]
  wire  _GEN_1544; // @[Execute.scala 117:10]
  wire  _GEN_1545; // @[Execute.scala 117:10]
  wire  _GEN_1546; // @[Execute.scala 117:10]
  wire  _GEN_1547; // @[Execute.scala 117:10]
  wire  _GEN_1548; // @[Execute.scala 117:10]
  wire  _GEN_1549; // @[Execute.scala 117:10]
  wire  _GEN_1550; // @[Execute.scala 117:10]
  wire  _GEN_1551; // @[Execute.scala 117:10]
  wire  _GEN_1552; // @[Execute.scala 117:10]
  wire  _GEN_1553; // @[Execute.scala 117:10]
  wire  _GEN_1554; // @[Execute.scala 117:10]
  wire  _GEN_1555; // @[Execute.scala 117:10]
  wire  _GEN_1556; // @[Execute.scala 117:10]
  wire  _GEN_1557; // @[Execute.scala 117:10]
  wire  _GEN_1558; // @[Execute.scala 117:10]
  wire  _GEN_1559; // @[Execute.scala 117:10]
  wire  _GEN_1560; // @[Execute.scala 117:10]
  wire  _GEN_1561; // @[Execute.scala 117:10]
  wire  _GEN_1562; // @[Execute.scala 117:10]
  wire  _GEN_1563; // @[Execute.scala 117:10]
  wire  _GEN_1564; // @[Execute.scala 117:10]
  wire  _GEN_1565; // @[Execute.scala 117:10]
  wire  _GEN_1566; // @[Execute.scala 117:10]
  wire  _GEN_1567; // @[Execute.scala 117:10]
  wire  _GEN_1568; // @[Execute.scala 117:10]
  wire  _GEN_1569; // @[Execute.scala 117:10]
  wire  _GEN_1570; // @[Execute.scala 117:10]
  wire  _GEN_1571; // @[Execute.scala 117:10]
  wire  _GEN_1572; // @[Execute.scala 117:10]
  wire  _GEN_1573; // @[Execute.scala 117:10]
  wire  _GEN_1574; // @[Execute.scala 117:10]
  wire  _GEN_1575; // @[Execute.scala 117:10]
  wire  _GEN_1576; // @[Execute.scala 117:10]
  wire  _GEN_1577; // @[Execute.scala 117:10]
  wire  _GEN_1578; // @[Execute.scala 117:10]
  wire  _GEN_1579; // @[Execute.scala 117:10]
  wire  _GEN_1580; // @[Execute.scala 117:10]
  wire  _GEN_1581; // @[Execute.scala 117:10]
  wire  _GEN_1582; // @[Execute.scala 117:10]
  wire  _GEN_1583; // @[Execute.scala 117:10]
  wire  _GEN_1584; // @[Execute.scala 117:10]
  wire  _GEN_1585; // @[Execute.scala 117:10]
  wire  _GEN_1586; // @[Execute.scala 117:10]
  wire  _GEN_1587; // @[Execute.scala 117:10]
  wire  _GEN_1588; // @[Execute.scala 117:10]
  wire  _GEN_1589; // @[Execute.scala 117:10]
  wire  _GEN_1590; // @[Execute.scala 117:10]
  wire  _GEN_1591; // @[Execute.scala 117:10]
  wire  _GEN_1592; // @[Execute.scala 117:10]
  wire  _GEN_1593; // @[Execute.scala 117:10]
  wire  _GEN_1594; // @[Execute.scala 117:10]
  wire  _GEN_1595; // @[Execute.scala 117:10]
  wire  _GEN_1596; // @[Execute.scala 117:10]
  wire  _GEN_1597; // @[Execute.scala 117:10]
  wire  _GEN_1598; // @[Execute.scala 117:10]
  wire  _GEN_1599; // @[Execute.scala 117:10]
  wire  _GEN_1600; // @[Execute.scala 117:10]
  wire  _GEN_1601; // @[Execute.scala 117:10]
  wire  _GEN_1603; // @[Execute.scala 117:10]
  wire  _GEN_1604; // @[Execute.scala 117:10]
  wire  _GEN_1605; // @[Execute.scala 117:10]
  wire  _GEN_1606; // @[Execute.scala 117:10]
  wire  _GEN_1607; // @[Execute.scala 117:10]
  wire  _GEN_1608; // @[Execute.scala 117:10]
  wire  _GEN_1609; // @[Execute.scala 117:10]
  wire  _GEN_1610; // @[Execute.scala 117:10]
  wire  _GEN_1611; // @[Execute.scala 117:10]
  wire  _GEN_1612; // @[Execute.scala 117:10]
  wire  _GEN_1613; // @[Execute.scala 117:10]
  wire  _GEN_1614; // @[Execute.scala 117:10]
  wire  _GEN_1615; // @[Execute.scala 117:10]
  wire  _GEN_1616; // @[Execute.scala 117:10]
  wire  _GEN_1617; // @[Execute.scala 117:10]
  wire  _GEN_1618; // @[Execute.scala 117:10]
  wire  _GEN_1619; // @[Execute.scala 117:10]
  wire  _GEN_1620; // @[Execute.scala 117:10]
  wire  _GEN_1621; // @[Execute.scala 117:10]
  wire  _GEN_1622; // @[Execute.scala 117:10]
  wire  _GEN_1623; // @[Execute.scala 117:10]
  wire  _GEN_1624; // @[Execute.scala 117:10]
  wire  _GEN_1625; // @[Execute.scala 117:10]
  wire  _GEN_1626; // @[Execute.scala 117:10]
  wire  _GEN_1627; // @[Execute.scala 117:10]
  wire  _GEN_1628; // @[Execute.scala 117:10]
  wire  _GEN_1629; // @[Execute.scala 117:10]
  wire  _GEN_1630; // @[Execute.scala 117:10]
  wire  _GEN_1631; // @[Execute.scala 117:10]
  wire  _GEN_1632; // @[Execute.scala 117:10]
  wire  _GEN_1633; // @[Execute.scala 117:10]
  wire  _GEN_1634; // @[Execute.scala 117:10]
  wire  _GEN_1635; // @[Execute.scala 117:10]
  wire  _GEN_1636; // @[Execute.scala 117:10]
  wire  _GEN_1637; // @[Execute.scala 117:10]
  wire  _GEN_1638; // @[Execute.scala 117:10]
  wire  _GEN_1639; // @[Execute.scala 117:10]
  wire  _GEN_1640; // @[Execute.scala 117:10]
  wire  _GEN_1641; // @[Execute.scala 117:10]
  wire  _GEN_1642; // @[Execute.scala 117:10]
  wire  _GEN_1643; // @[Execute.scala 117:10]
  wire  _GEN_1644; // @[Execute.scala 117:10]
  wire  _GEN_1645; // @[Execute.scala 117:10]
  wire  _GEN_1646; // @[Execute.scala 117:10]
  wire  _GEN_1647; // @[Execute.scala 117:10]
  wire  _GEN_1648; // @[Execute.scala 117:10]
  wire  _GEN_1649; // @[Execute.scala 117:10]
  wire  _GEN_1650; // @[Execute.scala 117:10]
  wire  _GEN_1651; // @[Execute.scala 117:10]
  wire  _GEN_1652; // @[Execute.scala 117:10]
  wire  _GEN_1653; // @[Execute.scala 117:10]
  wire  _GEN_1654; // @[Execute.scala 117:10]
  wire  _GEN_1655; // @[Execute.scala 117:10]
  wire  _GEN_1656; // @[Execute.scala 117:10]
  wire  _GEN_1657; // @[Execute.scala 117:10]
  wire  _GEN_1658; // @[Execute.scala 117:10]
  wire  _GEN_1659; // @[Execute.scala 117:10]
  wire  _GEN_1660; // @[Execute.scala 117:10]
  wire  _GEN_1661; // @[Execute.scala 117:10]
  wire  _GEN_1662; // @[Execute.scala 117:10]
  wire  _GEN_1663; // @[Execute.scala 117:10]
  wire  _GEN_1664; // @[Execute.scala 117:10]
  wire  _GEN_1665; // @[Execute.scala 117:10]
  wire  _T_211; // @[Execute.scala 117:10]
  wire  _T_212; // @[Execute.scala 117:15]
  wire [5:0] _T_214; // @[Execute.scala 117:37]
  wire [5:0] _T_218; // @[Execute.scala 117:60]
  wire  _GEN_1667; // @[Execute.scala 117:10]
  wire  _GEN_1668; // @[Execute.scala 117:10]
  wire  _GEN_1669; // @[Execute.scala 117:10]
  wire  _GEN_1670; // @[Execute.scala 117:10]
  wire  _GEN_1671; // @[Execute.scala 117:10]
  wire  _GEN_1672; // @[Execute.scala 117:10]
  wire  _GEN_1673; // @[Execute.scala 117:10]
  wire  _GEN_1674; // @[Execute.scala 117:10]
  wire  _GEN_1675; // @[Execute.scala 117:10]
  wire  _GEN_1676; // @[Execute.scala 117:10]
  wire  _GEN_1677; // @[Execute.scala 117:10]
  wire  _GEN_1678; // @[Execute.scala 117:10]
  wire  _GEN_1679; // @[Execute.scala 117:10]
  wire  _GEN_1680; // @[Execute.scala 117:10]
  wire  _GEN_1681; // @[Execute.scala 117:10]
  wire  _GEN_1682; // @[Execute.scala 117:10]
  wire  _GEN_1683; // @[Execute.scala 117:10]
  wire  _GEN_1684; // @[Execute.scala 117:10]
  wire  _GEN_1685; // @[Execute.scala 117:10]
  wire  _GEN_1686; // @[Execute.scala 117:10]
  wire  _GEN_1687; // @[Execute.scala 117:10]
  wire  _GEN_1688; // @[Execute.scala 117:10]
  wire  _GEN_1689; // @[Execute.scala 117:10]
  wire  _GEN_1690; // @[Execute.scala 117:10]
  wire  _GEN_1691; // @[Execute.scala 117:10]
  wire  _GEN_1692; // @[Execute.scala 117:10]
  wire  _GEN_1693; // @[Execute.scala 117:10]
  wire  _GEN_1694; // @[Execute.scala 117:10]
  wire  _GEN_1695; // @[Execute.scala 117:10]
  wire  _GEN_1696; // @[Execute.scala 117:10]
  wire  _GEN_1697; // @[Execute.scala 117:10]
  wire  _GEN_1698; // @[Execute.scala 117:10]
  wire  _GEN_1699; // @[Execute.scala 117:10]
  wire  _GEN_1700; // @[Execute.scala 117:10]
  wire  _GEN_1701; // @[Execute.scala 117:10]
  wire  _GEN_1702; // @[Execute.scala 117:10]
  wire  _GEN_1703; // @[Execute.scala 117:10]
  wire  _GEN_1704; // @[Execute.scala 117:10]
  wire  _GEN_1705; // @[Execute.scala 117:10]
  wire  _GEN_1706; // @[Execute.scala 117:10]
  wire  _GEN_1707; // @[Execute.scala 117:10]
  wire  _GEN_1708; // @[Execute.scala 117:10]
  wire  _GEN_1709; // @[Execute.scala 117:10]
  wire  _GEN_1710; // @[Execute.scala 117:10]
  wire  _GEN_1711; // @[Execute.scala 117:10]
  wire  _GEN_1712; // @[Execute.scala 117:10]
  wire  _GEN_1713; // @[Execute.scala 117:10]
  wire  _GEN_1714; // @[Execute.scala 117:10]
  wire  _GEN_1715; // @[Execute.scala 117:10]
  wire  _GEN_1716; // @[Execute.scala 117:10]
  wire  _GEN_1717; // @[Execute.scala 117:10]
  wire  _GEN_1718; // @[Execute.scala 117:10]
  wire  _GEN_1719; // @[Execute.scala 117:10]
  wire  _GEN_1720; // @[Execute.scala 117:10]
  wire  _GEN_1721; // @[Execute.scala 117:10]
  wire  _GEN_1722; // @[Execute.scala 117:10]
  wire  _GEN_1723; // @[Execute.scala 117:10]
  wire  _GEN_1724; // @[Execute.scala 117:10]
  wire  _GEN_1725; // @[Execute.scala 117:10]
  wire  _GEN_1726; // @[Execute.scala 117:10]
  wire  _GEN_1727; // @[Execute.scala 117:10]
  wire  _GEN_1728; // @[Execute.scala 117:10]
  wire  _GEN_1729; // @[Execute.scala 117:10]
  wire  _GEN_1731; // @[Execute.scala 117:10]
  wire  _GEN_1732; // @[Execute.scala 117:10]
  wire  _GEN_1733; // @[Execute.scala 117:10]
  wire  _GEN_1734; // @[Execute.scala 117:10]
  wire  _GEN_1735; // @[Execute.scala 117:10]
  wire  _GEN_1736; // @[Execute.scala 117:10]
  wire  _GEN_1737; // @[Execute.scala 117:10]
  wire  _GEN_1738; // @[Execute.scala 117:10]
  wire  _GEN_1739; // @[Execute.scala 117:10]
  wire  _GEN_1740; // @[Execute.scala 117:10]
  wire  _GEN_1741; // @[Execute.scala 117:10]
  wire  _GEN_1742; // @[Execute.scala 117:10]
  wire  _GEN_1743; // @[Execute.scala 117:10]
  wire  _GEN_1744; // @[Execute.scala 117:10]
  wire  _GEN_1745; // @[Execute.scala 117:10]
  wire  _GEN_1746; // @[Execute.scala 117:10]
  wire  _GEN_1747; // @[Execute.scala 117:10]
  wire  _GEN_1748; // @[Execute.scala 117:10]
  wire  _GEN_1749; // @[Execute.scala 117:10]
  wire  _GEN_1750; // @[Execute.scala 117:10]
  wire  _GEN_1751; // @[Execute.scala 117:10]
  wire  _GEN_1752; // @[Execute.scala 117:10]
  wire  _GEN_1753; // @[Execute.scala 117:10]
  wire  _GEN_1754; // @[Execute.scala 117:10]
  wire  _GEN_1755; // @[Execute.scala 117:10]
  wire  _GEN_1756; // @[Execute.scala 117:10]
  wire  _GEN_1757; // @[Execute.scala 117:10]
  wire  _GEN_1758; // @[Execute.scala 117:10]
  wire  _GEN_1759; // @[Execute.scala 117:10]
  wire  _GEN_1760; // @[Execute.scala 117:10]
  wire  _GEN_1761; // @[Execute.scala 117:10]
  wire  _GEN_1762; // @[Execute.scala 117:10]
  wire  _GEN_1763; // @[Execute.scala 117:10]
  wire  _GEN_1764; // @[Execute.scala 117:10]
  wire  _GEN_1765; // @[Execute.scala 117:10]
  wire  _GEN_1766; // @[Execute.scala 117:10]
  wire  _GEN_1767; // @[Execute.scala 117:10]
  wire  _GEN_1768; // @[Execute.scala 117:10]
  wire  _GEN_1769; // @[Execute.scala 117:10]
  wire  _GEN_1770; // @[Execute.scala 117:10]
  wire  _GEN_1771; // @[Execute.scala 117:10]
  wire  _GEN_1772; // @[Execute.scala 117:10]
  wire  _GEN_1773; // @[Execute.scala 117:10]
  wire  _GEN_1774; // @[Execute.scala 117:10]
  wire  _GEN_1775; // @[Execute.scala 117:10]
  wire  _GEN_1776; // @[Execute.scala 117:10]
  wire  _GEN_1777; // @[Execute.scala 117:10]
  wire  _GEN_1778; // @[Execute.scala 117:10]
  wire  _GEN_1779; // @[Execute.scala 117:10]
  wire  _GEN_1780; // @[Execute.scala 117:10]
  wire  _GEN_1781; // @[Execute.scala 117:10]
  wire  _GEN_1782; // @[Execute.scala 117:10]
  wire  _GEN_1783; // @[Execute.scala 117:10]
  wire  _GEN_1784; // @[Execute.scala 117:10]
  wire  _GEN_1785; // @[Execute.scala 117:10]
  wire  _GEN_1786; // @[Execute.scala 117:10]
  wire  _GEN_1787; // @[Execute.scala 117:10]
  wire  _GEN_1788; // @[Execute.scala 117:10]
  wire  _GEN_1789; // @[Execute.scala 117:10]
  wire  _GEN_1790; // @[Execute.scala 117:10]
  wire  _GEN_1791; // @[Execute.scala 117:10]
  wire  _GEN_1792; // @[Execute.scala 117:10]
  wire  _GEN_1793; // @[Execute.scala 117:10]
  wire  _T_221; // @[Execute.scala 117:10]
  wire  _T_222; // @[Execute.scala 117:15]
  wire [5:0] _T_224; // @[Execute.scala 117:37]
  wire [5:0] _T_228; // @[Execute.scala 117:60]
  wire  _GEN_1795; // @[Execute.scala 117:10]
  wire  _GEN_1796; // @[Execute.scala 117:10]
  wire  _GEN_1797; // @[Execute.scala 117:10]
  wire  _GEN_1798; // @[Execute.scala 117:10]
  wire  _GEN_1799; // @[Execute.scala 117:10]
  wire  _GEN_1800; // @[Execute.scala 117:10]
  wire  _GEN_1801; // @[Execute.scala 117:10]
  wire  _GEN_1802; // @[Execute.scala 117:10]
  wire  _GEN_1803; // @[Execute.scala 117:10]
  wire  _GEN_1804; // @[Execute.scala 117:10]
  wire  _GEN_1805; // @[Execute.scala 117:10]
  wire  _GEN_1806; // @[Execute.scala 117:10]
  wire  _GEN_1807; // @[Execute.scala 117:10]
  wire  _GEN_1808; // @[Execute.scala 117:10]
  wire  _GEN_1809; // @[Execute.scala 117:10]
  wire  _GEN_1810; // @[Execute.scala 117:10]
  wire  _GEN_1811; // @[Execute.scala 117:10]
  wire  _GEN_1812; // @[Execute.scala 117:10]
  wire  _GEN_1813; // @[Execute.scala 117:10]
  wire  _GEN_1814; // @[Execute.scala 117:10]
  wire  _GEN_1815; // @[Execute.scala 117:10]
  wire  _GEN_1816; // @[Execute.scala 117:10]
  wire  _GEN_1817; // @[Execute.scala 117:10]
  wire  _GEN_1818; // @[Execute.scala 117:10]
  wire  _GEN_1819; // @[Execute.scala 117:10]
  wire  _GEN_1820; // @[Execute.scala 117:10]
  wire  _GEN_1821; // @[Execute.scala 117:10]
  wire  _GEN_1822; // @[Execute.scala 117:10]
  wire  _GEN_1823; // @[Execute.scala 117:10]
  wire  _GEN_1824; // @[Execute.scala 117:10]
  wire  _GEN_1825; // @[Execute.scala 117:10]
  wire  _GEN_1826; // @[Execute.scala 117:10]
  wire  _GEN_1827; // @[Execute.scala 117:10]
  wire  _GEN_1828; // @[Execute.scala 117:10]
  wire  _GEN_1829; // @[Execute.scala 117:10]
  wire  _GEN_1830; // @[Execute.scala 117:10]
  wire  _GEN_1831; // @[Execute.scala 117:10]
  wire  _GEN_1832; // @[Execute.scala 117:10]
  wire  _GEN_1833; // @[Execute.scala 117:10]
  wire  _GEN_1834; // @[Execute.scala 117:10]
  wire  _GEN_1835; // @[Execute.scala 117:10]
  wire  _GEN_1836; // @[Execute.scala 117:10]
  wire  _GEN_1837; // @[Execute.scala 117:10]
  wire  _GEN_1838; // @[Execute.scala 117:10]
  wire  _GEN_1839; // @[Execute.scala 117:10]
  wire  _GEN_1840; // @[Execute.scala 117:10]
  wire  _GEN_1841; // @[Execute.scala 117:10]
  wire  _GEN_1842; // @[Execute.scala 117:10]
  wire  _GEN_1843; // @[Execute.scala 117:10]
  wire  _GEN_1844; // @[Execute.scala 117:10]
  wire  _GEN_1845; // @[Execute.scala 117:10]
  wire  _GEN_1846; // @[Execute.scala 117:10]
  wire  _GEN_1847; // @[Execute.scala 117:10]
  wire  _GEN_1848; // @[Execute.scala 117:10]
  wire  _GEN_1849; // @[Execute.scala 117:10]
  wire  _GEN_1850; // @[Execute.scala 117:10]
  wire  _GEN_1851; // @[Execute.scala 117:10]
  wire  _GEN_1852; // @[Execute.scala 117:10]
  wire  _GEN_1853; // @[Execute.scala 117:10]
  wire  _GEN_1854; // @[Execute.scala 117:10]
  wire  _GEN_1855; // @[Execute.scala 117:10]
  wire  _GEN_1856; // @[Execute.scala 117:10]
  wire  _GEN_1857; // @[Execute.scala 117:10]
  wire  _GEN_1859; // @[Execute.scala 117:10]
  wire  _GEN_1860; // @[Execute.scala 117:10]
  wire  _GEN_1861; // @[Execute.scala 117:10]
  wire  _GEN_1862; // @[Execute.scala 117:10]
  wire  _GEN_1863; // @[Execute.scala 117:10]
  wire  _GEN_1864; // @[Execute.scala 117:10]
  wire  _GEN_1865; // @[Execute.scala 117:10]
  wire  _GEN_1866; // @[Execute.scala 117:10]
  wire  _GEN_1867; // @[Execute.scala 117:10]
  wire  _GEN_1868; // @[Execute.scala 117:10]
  wire  _GEN_1869; // @[Execute.scala 117:10]
  wire  _GEN_1870; // @[Execute.scala 117:10]
  wire  _GEN_1871; // @[Execute.scala 117:10]
  wire  _GEN_1872; // @[Execute.scala 117:10]
  wire  _GEN_1873; // @[Execute.scala 117:10]
  wire  _GEN_1874; // @[Execute.scala 117:10]
  wire  _GEN_1875; // @[Execute.scala 117:10]
  wire  _GEN_1876; // @[Execute.scala 117:10]
  wire  _GEN_1877; // @[Execute.scala 117:10]
  wire  _GEN_1878; // @[Execute.scala 117:10]
  wire  _GEN_1879; // @[Execute.scala 117:10]
  wire  _GEN_1880; // @[Execute.scala 117:10]
  wire  _GEN_1881; // @[Execute.scala 117:10]
  wire  _GEN_1882; // @[Execute.scala 117:10]
  wire  _GEN_1883; // @[Execute.scala 117:10]
  wire  _GEN_1884; // @[Execute.scala 117:10]
  wire  _GEN_1885; // @[Execute.scala 117:10]
  wire  _GEN_1886; // @[Execute.scala 117:10]
  wire  _GEN_1887; // @[Execute.scala 117:10]
  wire  _GEN_1888; // @[Execute.scala 117:10]
  wire  _GEN_1889; // @[Execute.scala 117:10]
  wire  _GEN_1890; // @[Execute.scala 117:10]
  wire  _GEN_1891; // @[Execute.scala 117:10]
  wire  _GEN_1892; // @[Execute.scala 117:10]
  wire  _GEN_1893; // @[Execute.scala 117:10]
  wire  _GEN_1894; // @[Execute.scala 117:10]
  wire  _GEN_1895; // @[Execute.scala 117:10]
  wire  _GEN_1896; // @[Execute.scala 117:10]
  wire  _GEN_1897; // @[Execute.scala 117:10]
  wire  _GEN_1898; // @[Execute.scala 117:10]
  wire  _GEN_1899; // @[Execute.scala 117:10]
  wire  _GEN_1900; // @[Execute.scala 117:10]
  wire  _GEN_1901; // @[Execute.scala 117:10]
  wire  _GEN_1902; // @[Execute.scala 117:10]
  wire  _GEN_1903; // @[Execute.scala 117:10]
  wire  _GEN_1904; // @[Execute.scala 117:10]
  wire  _GEN_1905; // @[Execute.scala 117:10]
  wire  _GEN_1906; // @[Execute.scala 117:10]
  wire  _GEN_1907; // @[Execute.scala 117:10]
  wire  _GEN_1908; // @[Execute.scala 117:10]
  wire  _GEN_1909; // @[Execute.scala 117:10]
  wire  _GEN_1910; // @[Execute.scala 117:10]
  wire  _GEN_1911; // @[Execute.scala 117:10]
  wire  _GEN_1912; // @[Execute.scala 117:10]
  wire  _GEN_1913; // @[Execute.scala 117:10]
  wire  _GEN_1914; // @[Execute.scala 117:10]
  wire  _GEN_1915; // @[Execute.scala 117:10]
  wire  _GEN_1916; // @[Execute.scala 117:10]
  wire  _GEN_1917; // @[Execute.scala 117:10]
  wire  _GEN_1918; // @[Execute.scala 117:10]
  wire  _GEN_1919; // @[Execute.scala 117:10]
  wire  _GEN_1920; // @[Execute.scala 117:10]
  wire  _GEN_1921; // @[Execute.scala 117:10]
  wire  _T_231; // @[Execute.scala 117:10]
  wire  _T_232; // @[Execute.scala 117:15]
  wire [5:0] _T_234; // @[Execute.scala 117:37]
  wire [5:0] _T_238; // @[Execute.scala 117:60]
  wire  _GEN_1923; // @[Execute.scala 117:10]
  wire  _GEN_1924; // @[Execute.scala 117:10]
  wire  _GEN_1925; // @[Execute.scala 117:10]
  wire  _GEN_1926; // @[Execute.scala 117:10]
  wire  _GEN_1927; // @[Execute.scala 117:10]
  wire  _GEN_1928; // @[Execute.scala 117:10]
  wire  _GEN_1929; // @[Execute.scala 117:10]
  wire  _GEN_1930; // @[Execute.scala 117:10]
  wire  _GEN_1931; // @[Execute.scala 117:10]
  wire  _GEN_1932; // @[Execute.scala 117:10]
  wire  _GEN_1933; // @[Execute.scala 117:10]
  wire  _GEN_1934; // @[Execute.scala 117:10]
  wire  _GEN_1935; // @[Execute.scala 117:10]
  wire  _GEN_1936; // @[Execute.scala 117:10]
  wire  _GEN_1937; // @[Execute.scala 117:10]
  wire  _GEN_1938; // @[Execute.scala 117:10]
  wire  _GEN_1939; // @[Execute.scala 117:10]
  wire  _GEN_1940; // @[Execute.scala 117:10]
  wire  _GEN_1941; // @[Execute.scala 117:10]
  wire  _GEN_1942; // @[Execute.scala 117:10]
  wire  _GEN_1943; // @[Execute.scala 117:10]
  wire  _GEN_1944; // @[Execute.scala 117:10]
  wire  _GEN_1945; // @[Execute.scala 117:10]
  wire  _GEN_1946; // @[Execute.scala 117:10]
  wire  _GEN_1947; // @[Execute.scala 117:10]
  wire  _GEN_1948; // @[Execute.scala 117:10]
  wire  _GEN_1949; // @[Execute.scala 117:10]
  wire  _GEN_1950; // @[Execute.scala 117:10]
  wire  _GEN_1951; // @[Execute.scala 117:10]
  wire  _GEN_1952; // @[Execute.scala 117:10]
  wire  _GEN_1953; // @[Execute.scala 117:10]
  wire  _GEN_1954; // @[Execute.scala 117:10]
  wire  _GEN_1955; // @[Execute.scala 117:10]
  wire  _GEN_1956; // @[Execute.scala 117:10]
  wire  _GEN_1957; // @[Execute.scala 117:10]
  wire  _GEN_1958; // @[Execute.scala 117:10]
  wire  _GEN_1959; // @[Execute.scala 117:10]
  wire  _GEN_1960; // @[Execute.scala 117:10]
  wire  _GEN_1961; // @[Execute.scala 117:10]
  wire  _GEN_1962; // @[Execute.scala 117:10]
  wire  _GEN_1963; // @[Execute.scala 117:10]
  wire  _GEN_1964; // @[Execute.scala 117:10]
  wire  _GEN_1965; // @[Execute.scala 117:10]
  wire  _GEN_1966; // @[Execute.scala 117:10]
  wire  _GEN_1967; // @[Execute.scala 117:10]
  wire  _GEN_1968; // @[Execute.scala 117:10]
  wire  _GEN_1969; // @[Execute.scala 117:10]
  wire  _GEN_1970; // @[Execute.scala 117:10]
  wire  _GEN_1971; // @[Execute.scala 117:10]
  wire  _GEN_1972; // @[Execute.scala 117:10]
  wire  _GEN_1973; // @[Execute.scala 117:10]
  wire  _GEN_1974; // @[Execute.scala 117:10]
  wire  _GEN_1975; // @[Execute.scala 117:10]
  wire  _GEN_1976; // @[Execute.scala 117:10]
  wire  _GEN_1977; // @[Execute.scala 117:10]
  wire  _GEN_1978; // @[Execute.scala 117:10]
  wire  _GEN_1979; // @[Execute.scala 117:10]
  wire  _GEN_1980; // @[Execute.scala 117:10]
  wire  _GEN_1981; // @[Execute.scala 117:10]
  wire  _GEN_1982; // @[Execute.scala 117:10]
  wire  _GEN_1983; // @[Execute.scala 117:10]
  wire  _GEN_1984; // @[Execute.scala 117:10]
  wire  _GEN_1985; // @[Execute.scala 117:10]
  wire  _GEN_1987; // @[Execute.scala 117:10]
  wire  _GEN_1988; // @[Execute.scala 117:10]
  wire  _GEN_1989; // @[Execute.scala 117:10]
  wire  _GEN_1990; // @[Execute.scala 117:10]
  wire  _GEN_1991; // @[Execute.scala 117:10]
  wire  _GEN_1992; // @[Execute.scala 117:10]
  wire  _GEN_1993; // @[Execute.scala 117:10]
  wire  _GEN_1994; // @[Execute.scala 117:10]
  wire  _GEN_1995; // @[Execute.scala 117:10]
  wire  _GEN_1996; // @[Execute.scala 117:10]
  wire  _GEN_1997; // @[Execute.scala 117:10]
  wire  _GEN_1998; // @[Execute.scala 117:10]
  wire  _GEN_1999; // @[Execute.scala 117:10]
  wire  _GEN_2000; // @[Execute.scala 117:10]
  wire  _GEN_2001; // @[Execute.scala 117:10]
  wire  _GEN_2002; // @[Execute.scala 117:10]
  wire  _GEN_2003; // @[Execute.scala 117:10]
  wire  _GEN_2004; // @[Execute.scala 117:10]
  wire  _GEN_2005; // @[Execute.scala 117:10]
  wire  _GEN_2006; // @[Execute.scala 117:10]
  wire  _GEN_2007; // @[Execute.scala 117:10]
  wire  _GEN_2008; // @[Execute.scala 117:10]
  wire  _GEN_2009; // @[Execute.scala 117:10]
  wire  _GEN_2010; // @[Execute.scala 117:10]
  wire  _GEN_2011; // @[Execute.scala 117:10]
  wire  _GEN_2012; // @[Execute.scala 117:10]
  wire  _GEN_2013; // @[Execute.scala 117:10]
  wire  _GEN_2014; // @[Execute.scala 117:10]
  wire  _GEN_2015; // @[Execute.scala 117:10]
  wire  _GEN_2016; // @[Execute.scala 117:10]
  wire  _GEN_2017; // @[Execute.scala 117:10]
  wire  _GEN_2018; // @[Execute.scala 117:10]
  wire  _GEN_2019; // @[Execute.scala 117:10]
  wire  _GEN_2020; // @[Execute.scala 117:10]
  wire  _GEN_2021; // @[Execute.scala 117:10]
  wire  _GEN_2022; // @[Execute.scala 117:10]
  wire  _GEN_2023; // @[Execute.scala 117:10]
  wire  _GEN_2024; // @[Execute.scala 117:10]
  wire  _GEN_2025; // @[Execute.scala 117:10]
  wire  _GEN_2026; // @[Execute.scala 117:10]
  wire  _GEN_2027; // @[Execute.scala 117:10]
  wire  _GEN_2028; // @[Execute.scala 117:10]
  wire  _GEN_2029; // @[Execute.scala 117:10]
  wire  _GEN_2030; // @[Execute.scala 117:10]
  wire  _GEN_2031; // @[Execute.scala 117:10]
  wire  _GEN_2032; // @[Execute.scala 117:10]
  wire  _GEN_2033; // @[Execute.scala 117:10]
  wire  _GEN_2034; // @[Execute.scala 117:10]
  wire  _GEN_2035; // @[Execute.scala 117:10]
  wire  _GEN_2036; // @[Execute.scala 117:10]
  wire  _GEN_2037; // @[Execute.scala 117:10]
  wire  _GEN_2038; // @[Execute.scala 117:10]
  wire  _GEN_2039; // @[Execute.scala 117:10]
  wire  _GEN_2040; // @[Execute.scala 117:10]
  wire  _GEN_2041; // @[Execute.scala 117:10]
  wire  _GEN_2042; // @[Execute.scala 117:10]
  wire  _GEN_2043; // @[Execute.scala 117:10]
  wire  _GEN_2044; // @[Execute.scala 117:10]
  wire  _GEN_2045; // @[Execute.scala 117:10]
  wire  _GEN_2046; // @[Execute.scala 117:10]
  wire  _GEN_2047; // @[Execute.scala 117:10]
  wire  _GEN_2048; // @[Execute.scala 117:10]
  wire  _GEN_2049; // @[Execute.scala 117:10]
  wire  _T_241; // @[Execute.scala 117:10]
  wire  _T_242; // @[Execute.scala 117:15]
  wire [5:0] _T_244; // @[Execute.scala 117:37]
  wire [5:0] _T_248; // @[Execute.scala 117:60]
  wire  _GEN_2051; // @[Execute.scala 117:10]
  wire  _GEN_2052; // @[Execute.scala 117:10]
  wire  _GEN_2053; // @[Execute.scala 117:10]
  wire  _GEN_2054; // @[Execute.scala 117:10]
  wire  _GEN_2055; // @[Execute.scala 117:10]
  wire  _GEN_2056; // @[Execute.scala 117:10]
  wire  _GEN_2057; // @[Execute.scala 117:10]
  wire  _GEN_2058; // @[Execute.scala 117:10]
  wire  _GEN_2059; // @[Execute.scala 117:10]
  wire  _GEN_2060; // @[Execute.scala 117:10]
  wire  _GEN_2061; // @[Execute.scala 117:10]
  wire  _GEN_2062; // @[Execute.scala 117:10]
  wire  _GEN_2063; // @[Execute.scala 117:10]
  wire  _GEN_2064; // @[Execute.scala 117:10]
  wire  _GEN_2065; // @[Execute.scala 117:10]
  wire  _GEN_2066; // @[Execute.scala 117:10]
  wire  _GEN_2067; // @[Execute.scala 117:10]
  wire  _GEN_2068; // @[Execute.scala 117:10]
  wire  _GEN_2069; // @[Execute.scala 117:10]
  wire  _GEN_2070; // @[Execute.scala 117:10]
  wire  _GEN_2071; // @[Execute.scala 117:10]
  wire  _GEN_2072; // @[Execute.scala 117:10]
  wire  _GEN_2073; // @[Execute.scala 117:10]
  wire  _GEN_2074; // @[Execute.scala 117:10]
  wire  _GEN_2075; // @[Execute.scala 117:10]
  wire  _GEN_2076; // @[Execute.scala 117:10]
  wire  _GEN_2077; // @[Execute.scala 117:10]
  wire  _GEN_2078; // @[Execute.scala 117:10]
  wire  _GEN_2079; // @[Execute.scala 117:10]
  wire  _GEN_2080; // @[Execute.scala 117:10]
  wire  _GEN_2081; // @[Execute.scala 117:10]
  wire  _GEN_2082; // @[Execute.scala 117:10]
  wire  _GEN_2083; // @[Execute.scala 117:10]
  wire  _GEN_2084; // @[Execute.scala 117:10]
  wire  _GEN_2085; // @[Execute.scala 117:10]
  wire  _GEN_2086; // @[Execute.scala 117:10]
  wire  _GEN_2087; // @[Execute.scala 117:10]
  wire  _GEN_2088; // @[Execute.scala 117:10]
  wire  _GEN_2089; // @[Execute.scala 117:10]
  wire  _GEN_2090; // @[Execute.scala 117:10]
  wire  _GEN_2091; // @[Execute.scala 117:10]
  wire  _GEN_2092; // @[Execute.scala 117:10]
  wire  _GEN_2093; // @[Execute.scala 117:10]
  wire  _GEN_2094; // @[Execute.scala 117:10]
  wire  _GEN_2095; // @[Execute.scala 117:10]
  wire  _GEN_2096; // @[Execute.scala 117:10]
  wire  _GEN_2097; // @[Execute.scala 117:10]
  wire  _GEN_2098; // @[Execute.scala 117:10]
  wire  _GEN_2099; // @[Execute.scala 117:10]
  wire  _GEN_2100; // @[Execute.scala 117:10]
  wire  _GEN_2101; // @[Execute.scala 117:10]
  wire  _GEN_2102; // @[Execute.scala 117:10]
  wire  _GEN_2103; // @[Execute.scala 117:10]
  wire  _GEN_2104; // @[Execute.scala 117:10]
  wire  _GEN_2105; // @[Execute.scala 117:10]
  wire  _GEN_2106; // @[Execute.scala 117:10]
  wire  _GEN_2107; // @[Execute.scala 117:10]
  wire  _GEN_2108; // @[Execute.scala 117:10]
  wire  _GEN_2109; // @[Execute.scala 117:10]
  wire  _GEN_2110; // @[Execute.scala 117:10]
  wire  _GEN_2111; // @[Execute.scala 117:10]
  wire  _GEN_2112; // @[Execute.scala 117:10]
  wire  _GEN_2113; // @[Execute.scala 117:10]
  wire  _GEN_2115; // @[Execute.scala 117:10]
  wire  _GEN_2116; // @[Execute.scala 117:10]
  wire  _GEN_2117; // @[Execute.scala 117:10]
  wire  _GEN_2118; // @[Execute.scala 117:10]
  wire  _GEN_2119; // @[Execute.scala 117:10]
  wire  _GEN_2120; // @[Execute.scala 117:10]
  wire  _GEN_2121; // @[Execute.scala 117:10]
  wire  _GEN_2122; // @[Execute.scala 117:10]
  wire  _GEN_2123; // @[Execute.scala 117:10]
  wire  _GEN_2124; // @[Execute.scala 117:10]
  wire  _GEN_2125; // @[Execute.scala 117:10]
  wire  _GEN_2126; // @[Execute.scala 117:10]
  wire  _GEN_2127; // @[Execute.scala 117:10]
  wire  _GEN_2128; // @[Execute.scala 117:10]
  wire  _GEN_2129; // @[Execute.scala 117:10]
  wire  _GEN_2130; // @[Execute.scala 117:10]
  wire  _GEN_2131; // @[Execute.scala 117:10]
  wire  _GEN_2132; // @[Execute.scala 117:10]
  wire  _GEN_2133; // @[Execute.scala 117:10]
  wire  _GEN_2134; // @[Execute.scala 117:10]
  wire  _GEN_2135; // @[Execute.scala 117:10]
  wire  _GEN_2136; // @[Execute.scala 117:10]
  wire  _GEN_2137; // @[Execute.scala 117:10]
  wire  _GEN_2138; // @[Execute.scala 117:10]
  wire  _GEN_2139; // @[Execute.scala 117:10]
  wire  _GEN_2140; // @[Execute.scala 117:10]
  wire  _GEN_2141; // @[Execute.scala 117:10]
  wire  _GEN_2142; // @[Execute.scala 117:10]
  wire  _GEN_2143; // @[Execute.scala 117:10]
  wire  _GEN_2144; // @[Execute.scala 117:10]
  wire  _GEN_2145; // @[Execute.scala 117:10]
  wire  _GEN_2146; // @[Execute.scala 117:10]
  wire  _GEN_2147; // @[Execute.scala 117:10]
  wire  _GEN_2148; // @[Execute.scala 117:10]
  wire  _GEN_2149; // @[Execute.scala 117:10]
  wire  _GEN_2150; // @[Execute.scala 117:10]
  wire  _GEN_2151; // @[Execute.scala 117:10]
  wire  _GEN_2152; // @[Execute.scala 117:10]
  wire  _GEN_2153; // @[Execute.scala 117:10]
  wire  _GEN_2154; // @[Execute.scala 117:10]
  wire  _GEN_2155; // @[Execute.scala 117:10]
  wire  _GEN_2156; // @[Execute.scala 117:10]
  wire  _GEN_2157; // @[Execute.scala 117:10]
  wire  _GEN_2158; // @[Execute.scala 117:10]
  wire  _GEN_2159; // @[Execute.scala 117:10]
  wire  _GEN_2160; // @[Execute.scala 117:10]
  wire  _GEN_2161; // @[Execute.scala 117:10]
  wire  _GEN_2162; // @[Execute.scala 117:10]
  wire  _GEN_2163; // @[Execute.scala 117:10]
  wire  _GEN_2164; // @[Execute.scala 117:10]
  wire  _GEN_2165; // @[Execute.scala 117:10]
  wire  _GEN_2166; // @[Execute.scala 117:10]
  wire  _GEN_2167; // @[Execute.scala 117:10]
  wire  _GEN_2168; // @[Execute.scala 117:10]
  wire  _GEN_2169; // @[Execute.scala 117:10]
  wire  _GEN_2170; // @[Execute.scala 117:10]
  wire  _GEN_2171; // @[Execute.scala 117:10]
  wire  _GEN_2172; // @[Execute.scala 117:10]
  wire  _GEN_2173; // @[Execute.scala 117:10]
  wire  _GEN_2174; // @[Execute.scala 117:10]
  wire  _GEN_2175; // @[Execute.scala 117:10]
  wire  _GEN_2176; // @[Execute.scala 117:10]
  wire  _GEN_2177; // @[Execute.scala 117:10]
  wire  _T_251; // @[Execute.scala 117:10]
  wire  _T_252; // @[Execute.scala 117:15]
  wire [5:0] _T_254; // @[Execute.scala 117:37]
  wire [5:0] _T_258; // @[Execute.scala 117:60]
  wire  _GEN_2179; // @[Execute.scala 117:10]
  wire  _GEN_2180; // @[Execute.scala 117:10]
  wire  _GEN_2181; // @[Execute.scala 117:10]
  wire  _GEN_2182; // @[Execute.scala 117:10]
  wire  _GEN_2183; // @[Execute.scala 117:10]
  wire  _GEN_2184; // @[Execute.scala 117:10]
  wire  _GEN_2185; // @[Execute.scala 117:10]
  wire  _GEN_2186; // @[Execute.scala 117:10]
  wire  _GEN_2187; // @[Execute.scala 117:10]
  wire  _GEN_2188; // @[Execute.scala 117:10]
  wire  _GEN_2189; // @[Execute.scala 117:10]
  wire  _GEN_2190; // @[Execute.scala 117:10]
  wire  _GEN_2191; // @[Execute.scala 117:10]
  wire  _GEN_2192; // @[Execute.scala 117:10]
  wire  _GEN_2193; // @[Execute.scala 117:10]
  wire  _GEN_2194; // @[Execute.scala 117:10]
  wire  _GEN_2195; // @[Execute.scala 117:10]
  wire  _GEN_2196; // @[Execute.scala 117:10]
  wire  _GEN_2197; // @[Execute.scala 117:10]
  wire  _GEN_2198; // @[Execute.scala 117:10]
  wire  _GEN_2199; // @[Execute.scala 117:10]
  wire  _GEN_2200; // @[Execute.scala 117:10]
  wire  _GEN_2201; // @[Execute.scala 117:10]
  wire  _GEN_2202; // @[Execute.scala 117:10]
  wire  _GEN_2203; // @[Execute.scala 117:10]
  wire  _GEN_2204; // @[Execute.scala 117:10]
  wire  _GEN_2205; // @[Execute.scala 117:10]
  wire  _GEN_2206; // @[Execute.scala 117:10]
  wire  _GEN_2207; // @[Execute.scala 117:10]
  wire  _GEN_2208; // @[Execute.scala 117:10]
  wire  _GEN_2209; // @[Execute.scala 117:10]
  wire  _GEN_2210; // @[Execute.scala 117:10]
  wire  _GEN_2211; // @[Execute.scala 117:10]
  wire  _GEN_2212; // @[Execute.scala 117:10]
  wire  _GEN_2213; // @[Execute.scala 117:10]
  wire  _GEN_2214; // @[Execute.scala 117:10]
  wire  _GEN_2215; // @[Execute.scala 117:10]
  wire  _GEN_2216; // @[Execute.scala 117:10]
  wire  _GEN_2217; // @[Execute.scala 117:10]
  wire  _GEN_2218; // @[Execute.scala 117:10]
  wire  _GEN_2219; // @[Execute.scala 117:10]
  wire  _GEN_2220; // @[Execute.scala 117:10]
  wire  _GEN_2221; // @[Execute.scala 117:10]
  wire  _GEN_2222; // @[Execute.scala 117:10]
  wire  _GEN_2223; // @[Execute.scala 117:10]
  wire  _GEN_2224; // @[Execute.scala 117:10]
  wire  _GEN_2225; // @[Execute.scala 117:10]
  wire  _GEN_2226; // @[Execute.scala 117:10]
  wire  _GEN_2227; // @[Execute.scala 117:10]
  wire  _GEN_2228; // @[Execute.scala 117:10]
  wire  _GEN_2229; // @[Execute.scala 117:10]
  wire  _GEN_2230; // @[Execute.scala 117:10]
  wire  _GEN_2231; // @[Execute.scala 117:10]
  wire  _GEN_2232; // @[Execute.scala 117:10]
  wire  _GEN_2233; // @[Execute.scala 117:10]
  wire  _GEN_2234; // @[Execute.scala 117:10]
  wire  _GEN_2235; // @[Execute.scala 117:10]
  wire  _GEN_2236; // @[Execute.scala 117:10]
  wire  _GEN_2237; // @[Execute.scala 117:10]
  wire  _GEN_2238; // @[Execute.scala 117:10]
  wire  _GEN_2239; // @[Execute.scala 117:10]
  wire  _GEN_2240; // @[Execute.scala 117:10]
  wire  _GEN_2241; // @[Execute.scala 117:10]
  wire  _GEN_2243; // @[Execute.scala 117:10]
  wire  _GEN_2244; // @[Execute.scala 117:10]
  wire  _GEN_2245; // @[Execute.scala 117:10]
  wire  _GEN_2246; // @[Execute.scala 117:10]
  wire  _GEN_2247; // @[Execute.scala 117:10]
  wire  _GEN_2248; // @[Execute.scala 117:10]
  wire  _GEN_2249; // @[Execute.scala 117:10]
  wire  _GEN_2250; // @[Execute.scala 117:10]
  wire  _GEN_2251; // @[Execute.scala 117:10]
  wire  _GEN_2252; // @[Execute.scala 117:10]
  wire  _GEN_2253; // @[Execute.scala 117:10]
  wire  _GEN_2254; // @[Execute.scala 117:10]
  wire  _GEN_2255; // @[Execute.scala 117:10]
  wire  _GEN_2256; // @[Execute.scala 117:10]
  wire  _GEN_2257; // @[Execute.scala 117:10]
  wire  _GEN_2258; // @[Execute.scala 117:10]
  wire  _GEN_2259; // @[Execute.scala 117:10]
  wire  _GEN_2260; // @[Execute.scala 117:10]
  wire  _GEN_2261; // @[Execute.scala 117:10]
  wire  _GEN_2262; // @[Execute.scala 117:10]
  wire  _GEN_2263; // @[Execute.scala 117:10]
  wire  _GEN_2264; // @[Execute.scala 117:10]
  wire  _GEN_2265; // @[Execute.scala 117:10]
  wire  _GEN_2266; // @[Execute.scala 117:10]
  wire  _GEN_2267; // @[Execute.scala 117:10]
  wire  _GEN_2268; // @[Execute.scala 117:10]
  wire  _GEN_2269; // @[Execute.scala 117:10]
  wire  _GEN_2270; // @[Execute.scala 117:10]
  wire  _GEN_2271; // @[Execute.scala 117:10]
  wire  _GEN_2272; // @[Execute.scala 117:10]
  wire  _GEN_2273; // @[Execute.scala 117:10]
  wire  _GEN_2274; // @[Execute.scala 117:10]
  wire  _GEN_2275; // @[Execute.scala 117:10]
  wire  _GEN_2276; // @[Execute.scala 117:10]
  wire  _GEN_2277; // @[Execute.scala 117:10]
  wire  _GEN_2278; // @[Execute.scala 117:10]
  wire  _GEN_2279; // @[Execute.scala 117:10]
  wire  _GEN_2280; // @[Execute.scala 117:10]
  wire  _GEN_2281; // @[Execute.scala 117:10]
  wire  _GEN_2282; // @[Execute.scala 117:10]
  wire  _GEN_2283; // @[Execute.scala 117:10]
  wire  _GEN_2284; // @[Execute.scala 117:10]
  wire  _GEN_2285; // @[Execute.scala 117:10]
  wire  _GEN_2286; // @[Execute.scala 117:10]
  wire  _GEN_2287; // @[Execute.scala 117:10]
  wire  _GEN_2288; // @[Execute.scala 117:10]
  wire  _GEN_2289; // @[Execute.scala 117:10]
  wire  _GEN_2290; // @[Execute.scala 117:10]
  wire  _GEN_2291; // @[Execute.scala 117:10]
  wire  _GEN_2292; // @[Execute.scala 117:10]
  wire  _GEN_2293; // @[Execute.scala 117:10]
  wire  _GEN_2294; // @[Execute.scala 117:10]
  wire  _GEN_2295; // @[Execute.scala 117:10]
  wire  _GEN_2296; // @[Execute.scala 117:10]
  wire  _GEN_2297; // @[Execute.scala 117:10]
  wire  _GEN_2298; // @[Execute.scala 117:10]
  wire  _GEN_2299; // @[Execute.scala 117:10]
  wire  _GEN_2300; // @[Execute.scala 117:10]
  wire  _GEN_2301; // @[Execute.scala 117:10]
  wire  _GEN_2302; // @[Execute.scala 117:10]
  wire  _GEN_2303; // @[Execute.scala 117:10]
  wire  _GEN_2304; // @[Execute.scala 117:10]
  wire  _GEN_2305; // @[Execute.scala 117:10]
  wire  _T_261; // @[Execute.scala 117:10]
  wire  _T_262; // @[Execute.scala 117:15]
  wire [5:0] _T_264; // @[Execute.scala 117:37]
  wire [5:0] _T_268; // @[Execute.scala 117:60]
  wire  _GEN_2307; // @[Execute.scala 117:10]
  wire  _GEN_2308; // @[Execute.scala 117:10]
  wire  _GEN_2309; // @[Execute.scala 117:10]
  wire  _GEN_2310; // @[Execute.scala 117:10]
  wire  _GEN_2311; // @[Execute.scala 117:10]
  wire  _GEN_2312; // @[Execute.scala 117:10]
  wire  _GEN_2313; // @[Execute.scala 117:10]
  wire  _GEN_2314; // @[Execute.scala 117:10]
  wire  _GEN_2315; // @[Execute.scala 117:10]
  wire  _GEN_2316; // @[Execute.scala 117:10]
  wire  _GEN_2317; // @[Execute.scala 117:10]
  wire  _GEN_2318; // @[Execute.scala 117:10]
  wire  _GEN_2319; // @[Execute.scala 117:10]
  wire  _GEN_2320; // @[Execute.scala 117:10]
  wire  _GEN_2321; // @[Execute.scala 117:10]
  wire  _GEN_2322; // @[Execute.scala 117:10]
  wire  _GEN_2323; // @[Execute.scala 117:10]
  wire  _GEN_2324; // @[Execute.scala 117:10]
  wire  _GEN_2325; // @[Execute.scala 117:10]
  wire  _GEN_2326; // @[Execute.scala 117:10]
  wire  _GEN_2327; // @[Execute.scala 117:10]
  wire  _GEN_2328; // @[Execute.scala 117:10]
  wire  _GEN_2329; // @[Execute.scala 117:10]
  wire  _GEN_2330; // @[Execute.scala 117:10]
  wire  _GEN_2331; // @[Execute.scala 117:10]
  wire  _GEN_2332; // @[Execute.scala 117:10]
  wire  _GEN_2333; // @[Execute.scala 117:10]
  wire  _GEN_2334; // @[Execute.scala 117:10]
  wire  _GEN_2335; // @[Execute.scala 117:10]
  wire  _GEN_2336; // @[Execute.scala 117:10]
  wire  _GEN_2337; // @[Execute.scala 117:10]
  wire  _GEN_2338; // @[Execute.scala 117:10]
  wire  _GEN_2339; // @[Execute.scala 117:10]
  wire  _GEN_2340; // @[Execute.scala 117:10]
  wire  _GEN_2341; // @[Execute.scala 117:10]
  wire  _GEN_2342; // @[Execute.scala 117:10]
  wire  _GEN_2343; // @[Execute.scala 117:10]
  wire  _GEN_2344; // @[Execute.scala 117:10]
  wire  _GEN_2345; // @[Execute.scala 117:10]
  wire  _GEN_2346; // @[Execute.scala 117:10]
  wire  _GEN_2347; // @[Execute.scala 117:10]
  wire  _GEN_2348; // @[Execute.scala 117:10]
  wire  _GEN_2349; // @[Execute.scala 117:10]
  wire  _GEN_2350; // @[Execute.scala 117:10]
  wire  _GEN_2351; // @[Execute.scala 117:10]
  wire  _GEN_2352; // @[Execute.scala 117:10]
  wire  _GEN_2353; // @[Execute.scala 117:10]
  wire  _GEN_2354; // @[Execute.scala 117:10]
  wire  _GEN_2355; // @[Execute.scala 117:10]
  wire  _GEN_2356; // @[Execute.scala 117:10]
  wire  _GEN_2357; // @[Execute.scala 117:10]
  wire  _GEN_2358; // @[Execute.scala 117:10]
  wire  _GEN_2359; // @[Execute.scala 117:10]
  wire  _GEN_2360; // @[Execute.scala 117:10]
  wire  _GEN_2361; // @[Execute.scala 117:10]
  wire  _GEN_2362; // @[Execute.scala 117:10]
  wire  _GEN_2363; // @[Execute.scala 117:10]
  wire  _GEN_2364; // @[Execute.scala 117:10]
  wire  _GEN_2365; // @[Execute.scala 117:10]
  wire  _GEN_2366; // @[Execute.scala 117:10]
  wire  _GEN_2367; // @[Execute.scala 117:10]
  wire  _GEN_2368; // @[Execute.scala 117:10]
  wire  _GEN_2369; // @[Execute.scala 117:10]
  wire  _GEN_2371; // @[Execute.scala 117:10]
  wire  _GEN_2372; // @[Execute.scala 117:10]
  wire  _GEN_2373; // @[Execute.scala 117:10]
  wire  _GEN_2374; // @[Execute.scala 117:10]
  wire  _GEN_2375; // @[Execute.scala 117:10]
  wire  _GEN_2376; // @[Execute.scala 117:10]
  wire  _GEN_2377; // @[Execute.scala 117:10]
  wire  _GEN_2378; // @[Execute.scala 117:10]
  wire  _GEN_2379; // @[Execute.scala 117:10]
  wire  _GEN_2380; // @[Execute.scala 117:10]
  wire  _GEN_2381; // @[Execute.scala 117:10]
  wire  _GEN_2382; // @[Execute.scala 117:10]
  wire  _GEN_2383; // @[Execute.scala 117:10]
  wire  _GEN_2384; // @[Execute.scala 117:10]
  wire  _GEN_2385; // @[Execute.scala 117:10]
  wire  _GEN_2386; // @[Execute.scala 117:10]
  wire  _GEN_2387; // @[Execute.scala 117:10]
  wire  _GEN_2388; // @[Execute.scala 117:10]
  wire  _GEN_2389; // @[Execute.scala 117:10]
  wire  _GEN_2390; // @[Execute.scala 117:10]
  wire  _GEN_2391; // @[Execute.scala 117:10]
  wire  _GEN_2392; // @[Execute.scala 117:10]
  wire  _GEN_2393; // @[Execute.scala 117:10]
  wire  _GEN_2394; // @[Execute.scala 117:10]
  wire  _GEN_2395; // @[Execute.scala 117:10]
  wire  _GEN_2396; // @[Execute.scala 117:10]
  wire  _GEN_2397; // @[Execute.scala 117:10]
  wire  _GEN_2398; // @[Execute.scala 117:10]
  wire  _GEN_2399; // @[Execute.scala 117:10]
  wire  _GEN_2400; // @[Execute.scala 117:10]
  wire  _GEN_2401; // @[Execute.scala 117:10]
  wire  _GEN_2402; // @[Execute.scala 117:10]
  wire  _GEN_2403; // @[Execute.scala 117:10]
  wire  _GEN_2404; // @[Execute.scala 117:10]
  wire  _GEN_2405; // @[Execute.scala 117:10]
  wire  _GEN_2406; // @[Execute.scala 117:10]
  wire  _GEN_2407; // @[Execute.scala 117:10]
  wire  _GEN_2408; // @[Execute.scala 117:10]
  wire  _GEN_2409; // @[Execute.scala 117:10]
  wire  _GEN_2410; // @[Execute.scala 117:10]
  wire  _GEN_2411; // @[Execute.scala 117:10]
  wire  _GEN_2412; // @[Execute.scala 117:10]
  wire  _GEN_2413; // @[Execute.scala 117:10]
  wire  _GEN_2414; // @[Execute.scala 117:10]
  wire  _GEN_2415; // @[Execute.scala 117:10]
  wire  _GEN_2416; // @[Execute.scala 117:10]
  wire  _GEN_2417; // @[Execute.scala 117:10]
  wire  _GEN_2418; // @[Execute.scala 117:10]
  wire  _GEN_2419; // @[Execute.scala 117:10]
  wire  _GEN_2420; // @[Execute.scala 117:10]
  wire  _GEN_2421; // @[Execute.scala 117:10]
  wire  _GEN_2422; // @[Execute.scala 117:10]
  wire  _GEN_2423; // @[Execute.scala 117:10]
  wire  _GEN_2424; // @[Execute.scala 117:10]
  wire  _GEN_2425; // @[Execute.scala 117:10]
  wire  _GEN_2426; // @[Execute.scala 117:10]
  wire  _GEN_2427; // @[Execute.scala 117:10]
  wire  _GEN_2428; // @[Execute.scala 117:10]
  wire  _GEN_2429; // @[Execute.scala 117:10]
  wire  _GEN_2430; // @[Execute.scala 117:10]
  wire  _GEN_2431; // @[Execute.scala 117:10]
  wire  _GEN_2432; // @[Execute.scala 117:10]
  wire  _GEN_2433; // @[Execute.scala 117:10]
  wire  _T_271; // @[Execute.scala 117:10]
  wire  _T_272; // @[Execute.scala 117:15]
  wire [5:0] _T_274; // @[Execute.scala 117:37]
  wire [5:0] _T_278; // @[Execute.scala 117:60]
  wire  _GEN_2435; // @[Execute.scala 117:10]
  wire  _GEN_2436; // @[Execute.scala 117:10]
  wire  _GEN_2437; // @[Execute.scala 117:10]
  wire  _GEN_2438; // @[Execute.scala 117:10]
  wire  _GEN_2439; // @[Execute.scala 117:10]
  wire  _GEN_2440; // @[Execute.scala 117:10]
  wire  _GEN_2441; // @[Execute.scala 117:10]
  wire  _GEN_2442; // @[Execute.scala 117:10]
  wire  _GEN_2443; // @[Execute.scala 117:10]
  wire  _GEN_2444; // @[Execute.scala 117:10]
  wire  _GEN_2445; // @[Execute.scala 117:10]
  wire  _GEN_2446; // @[Execute.scala 117:10]
  wire  _GEN_2447; // @[Execute.scala 117:10]
  wire  _GEN_2448; // @[Execute.scala 117:10]
  wire  _GEN_2449; // @[Execute.scala 117:10]
  wire  _GEN_2450; // @[Execute.scala 117:10]
  wire  _GEN_2451; // @[Execute.scala 117:10]
  wire  _GEN_2452; // @[Execute.scala 117:10]
  wire  _GEN_2453; // @[Execute.scala 117:10]
  wire  _GEN_2454; // @[Execute.scala 117:10]
  wire  _GEN_2455; // @[Execute.scala 117:10]
  wire  _GEN_2456; // @[Execute.scala 117:10]
  wire  _GEN_2457; // @[Execute.scala 117:10]
  wire  _GEN_2458; // @[Execute.scala 117:10]
  wire  _GEN_2459; // @[Execute.scala 117:10]
  wire  _GEN_2460; // @[Execute.scala 117:10]
  wire  _GEN_2461; // @[Execute.scala 117:10]
  wire  _GEN_2462; // @[Execute.scala 117:10]
  wire  _GEN_2463; // @[Execute.scala 117:10]
  wire  _GEN_2464; // @[Execute.scala 117:10]
  wire  _GEN_2465; // @[Execute.scala 117:10]
  wire  _GEN_2466; // @[Execute.scala 117:10]
  wire  _GEN_2467; // @[Execute.scala 117:10]
  wire  _GEN_2468; // @[Execute.scala 117:10]
  wire  _GEN_2469; // @[Execute.scala 117:10]
  wire  _GEN_2470; // @[Execute.scala 117:10]
  wire  _GEN_2471; // @[Execute.scala 117:10]
  wire  _GEN_2472; // @[Execute.scala 117:10]
  wire  _GEN_2473; // @[Execute.scala 117:10]
  wire  _GEN_2474; // @[Execute.scala 117:10]
  wire  _GEN_2475; // @[Execute.scala 117:10]
  wire  _GEN_2476; // @[Execute.scala 117:10]
  wire  _GEN_2477; // @[Execute.scala 117:10]
  wire  _GEN_2478; // @[Execute.scala 117:10]
  wire  _GEN_2479; // @[Execute.scala 117:10]
  wire  _GEN_2480; // @[Execute.scala 117:10]
  wire  _GEN_2481; // @[Execute.scala 117:10]
  wire  _GEN_2482; // @[Execute.scala 117:10]
  wire  _GEN_2483; // @[Execute.scala 117:10]
  wire  _GEN_2484; // @[Execute.scala 117:10]
  wire  _GEN_2485; // @[Execute.scala 117:10]
  wire  _GEN_2486; // @[Execute.scala 117:10]
  wire  _GEN_2487; // @[Execute.scala 117:10]
  wire  _GEN_2488; // @[Execute.scala 117:10]
  wire  _GEN_2489; // @[Execute.scala 117:10]
  wire  _GEN_2490; // @[Execute.scala 117:10]
  wire  _GEN_2491; // @[Execute.scala 117:10]
  wire  _GEN_2492; // @[Execute.scala 117:10]
  wire  _GEN_2493; // @[Execute.scala 117:10]
  wire  _GEN_2494; // @[Execute.scala 117:10]
  wire  _GEN_2495; // @[Execute.scala 117:10]
  wire  _GEN_2496; // @[Execute.scala 117:10]
  wire  _GEN_2497; // @[Execute.scala 117:10]
  wire  _GEN_2499; // @[Execute.scala 117:10]
  wire  _GEN_2500; // @[Execute.scala 117:10]
  wire  _GEN_2501; // @[Execute.scala 117:10]
  wire  _GEN_2502; // @[Execute.scala 117:10]
  wire  _GEN_2503; // @[Execute.scala 117:10]
  wire  _GEN_2504; // @[Execute.scala 117:10]
  wire  _GEN_2505; // @[Execute.scala 117:10]
  wire  _GEN_2506; // @[Execute.scala 117:10]
  wire  _GEN_2507; // @[Execute.scala 117:10]
  wire  _GEN_2508; // @[Execute.scala 117:10]
  wire  _GEN_2509; // @[Execute.scala 117:10]
  wire  _GEN_2510; // @[Execute.scala 117:10]
  wire  _GEN_2511; // @[Execute.scala 117:10]
  wire  _GEN_2512; // @[Execute.scala 117:10]
  wire  _GEN_2513; // @[Execute.scala 117:10]
  wire  _GEN_2514; // @[Execute.scala 117:10]
  wire  _GEN_2515; // @[Execute.scala 117:10]
  wire  _GEN_2516; // @[Execute.scala 117:10]
  wire  _GEN_2517; // @[Execute.scala 117:10]
  wire  _GEN_2518; // @[Execute.scala 117:10]
  wire  _GEN_2519; // @[Execute.scala 117:10]
  wire  _GEN_2520; // @[Execute.scala 117:10]
  wire  _GEN_2521; // @[Execute.scala 117:10]
  wire  _GEN_2522; // @[Execute.scala 117:10]
  wire  _GEN_2523; // @[Execute.scala 117:10]
  wire  _GEN_2524; // @[Execute.scala 117:10]
  wire  _GEN_2525; // @[Execute.scala 117:10]
  wire  _GEN_2526; // @[Execute.scala 117:10]
  wire  _GEN_2527; // @[Execute.scala 117:10]
  wire  _GEN_2528; // @[Execute.scala 117:10]
  wire  _GEN_2529; // @[Execute.scala 117:10]
  wire  _GEN_2530; // @[Execute.scala 117:10]
  wire  _GEN_2531; // @[Execute.scala 117:10]
  wire  _GEN_2532; // @[Execute.scala 117:10]
  wire  _GEN_2533; // @[Execute.scala 117:10]
  wire  _GEN_2534; // @[Execute.scala 117:10]
  wire  _GEN_2535; // @[Execute.scala 117:10]
  wire  _GEN_2536; // @[Execute.scala 117:10]
  wire  _GEN_2537; // @[Execute.scala 117:10]
  wire  _GEN_2538; // @[Execute.scala 117:10]
  wire  _GEN_2539; // @[Execute.scala 117:10]
  wire  _GEN_2540; // @[Execute.scala 117:10]
  wire  _GEN_2541; // @[Execute.scala 117:10]
  wire  _GEN_2542; // @[Execute.scala 117:10]
  wire  _GEN_2543; // @[Execute.scala 117:10]
  wire  _GEN_2544; // @[Execute.scala 117:10]
  wire  _GEN_2545; // @[Execute.scala 117:10]
  wire  _GEN_2546; // @[Execute.scala 117:10]
  wire  _GEN_2547; // @[Execute.scala 117:10]
  wire  _GEN_2548; // @[Execute.scala 117:10]
  wire  _GEN_2549; // @[Execute.scala 117:10]
  wire  _GEN_2550; // @[Execute.scala 117:10]
  wire  _GEN_2551; // @[Execute.scala 117:10]
  wire  _GEN_2552; // @[Execute.scala 117:10]
  wire  _GEN_2553; // @[Execute.scala 117:10]
  wire  _GEN_2554; // @[Execute.scala 117:10]
  wire  _GEN_2555; // @[Execute.scala 117:10]
  wire  _GEN_2556; // @[Execute.scala 117:10]
  wire  _GEN_2557; // @[Execute.scala 117:10]
  wire  _GEN_2558; // @[Execute.scala 117:10]
  wire  _GEN_2559; // @[Execute.scala 117:10]
  wire  _GEN_2560; // @[Execute.scala 117:10]
  wire  _GEN_2561; // @[Execute.scala 117:10]
  wire  _T_281; // @[Execute.scala 117:10]
  wire  _T_282; // @[Execute.scala 117:15]
  wire [5:0] _T_284; // @[Execute.scala 117:37]
  wire [5:0] _T_288; // @[Execute.scala 117:60]
  wire  _GEN_2563; // @[Execute.scala 117:10]
  wire  _GEN_2564; // @[Execute.scala 117:10]
  wire  _GEN_2565; // @[Execute.scala 117:10]
  wire  _GEN_2566; // @[Execute.scala 117:10]
  wire  _GEN_2567; // @[Execute.scala 117:10]
  wire  _GEN_2568; // @[Execute.scala 117:10]
  wire  _GEN_2569; // @[Execute.scala 117:10]
  wire  _GEN_2570; // @[Execute.scala 117:10]
  wire  _GEN_2571; // @[Execute.scala 117:10]
  wire  _GEN_2572; // @[Execute.scala 117:10]
  wire  _GEN_2573; // @[Execute.scala 117:10]
  wire  _GEN_2574; // @[Execute.scala 117:10]
  wire  _GEN_2575; // @[Execute.scala 117:10]
  wire  _GEN_2576; // @[Execute.scala 117:10]
  wire  _GEN_2577; // @[Execute.scala 117:10]
  wire  _GEN_2578; // @[Execute.scala 117:10]
  wire  _GEN_2579; // @[Execute.scala 117:10]
  wire  _GEN_2580; // @[Execute.scala 117:10]
  wire  _GEN_2581; // @[Execute.scala 117:10]
  wire  _GEN_2582; // @[Execute.scala 117:10]
  wire  _GEN_2583; // @[Execute.scala 117:10]
  wire  _GEN_2584; // @[Execute.scala 117:10]
  wire  _GEN_2585; // @[Execute.scala 117:10]
  wire  _GEN_2586; // @[Execute.scala 117:10]
  wire  _GEN_2587; // @[Execute.scala 117:10]
  wire  _GEN_2588; // @[Execute.scala 117:10]
  wire  _GEN_2589; // @[Execute.scala 117:10]
  wire  _GEN_2590; // @[Execute.scala 117:10]
  wire  _GEN_2591; // @[Execute.scala 117:10]
  wire  _GEN_2592; // @[Execute.scala 117:10]
  wire  _GEN_2593; // @[Execute.scala 117:10]
  wire  _GEN_2594; // @[Execute.scala 117:10]
  wire  _GEN_2595; // @[Execute.scala 117:10]
  wire  _GEN_2596; // @[Execute.scala 117:10]
  wire  _GEN_2597; // @[Execute.scala 117:10]
  wire  _GEN_2598; // @[Execute.scala 117:10]
  wire  _GEN_2599; // @[Execute.scala 117:10]
  wire  _GEN_2600; // @[Execute.scala 117:10]
  wire  _GEN_2601; // @[Execute.scala 117:10]
  wire  _GEN_2602; // @[Execute.scala 117:10]
  wire  _GEN_2603; // @[Execute.scala 117:10]
  wire  _GEN_2604; // @[Execute.scala 117:10]
  wire  _GEN_2605; // @[Execute.scala 117:10]
  wire  _GEN_2606; // @[Execute.scala 117:10]
  wire  _GEN_2607; // @[Execute.scala 117:10]
  wire  _GEN_2608; // @[Execute.scala 117:10]
  wire  _GEN_2609; // @[Execute.scala 117:10]
  wire  _GEN_2610; // @[Execute.scala 117:10]
  wire  _GEN_2611; // @[Execute.scala 117:10]
  wire  _GEN_2612; // @[Execute.scala 117:10]
  wire  _GEN_2613; // @[Execute.scala 117:10]
  wire  _GEN_2614; // @[Execute.scala 117:10]
  wire  _GEN_2615; // @[Execute.scala 117:10]
  wire  _GEN_2616; // @[Execute.scala 117:10]
  wire  _GEN_2617; // @[Execute.scala 117:10]
  wire  _GEN_2618; // @[Execute.scala 117:10]
  wire  _GEN_2619; // @[Execute.scala 117:10]
  wire  _GEN_2620; // @[Execute.scala 117:10]
  wire  _GEN_2621; // @[Execute.scala 117:10]
  wire  _GEN_2622; // @[Execute.scala 117:10]
  wire  _GEN_2623; // @[Execute.scala 117:10]
  wire  _GEN_2624; // @[Execute.scala 117:10]
  wire  _GEN_2625; // @[Execute.scala 117:10]
  wire  _GEN_2627; // @[Execute.scala 117:10]
  wire  _GEN_2628; // @[Execute.scala 117:10]
  wire  _GEN_2629; // @[Execute.scala 117:10]
  wire  _GEN_2630; // @[Execute.scala 117:10]
  wire  _GEN_2631; // @[Execute.scala 117:10]
  wire  _GEN_2632; // @[Execute.scala 117:10]
  wire  _GEN_2633; // @[Execute.scala 117:10]
  wire  _GEN_2634; // @[Execute.scala 117:10]
  wire  _GEN_2635; // @[Execute.scala 117:10]
  wire  _GEN_2636; // @[Execute.scala 117:10]
  wire  _GEN_2637; // @[Execute.scala 117:10]
  wire  _GEN_2638; // @[Execute.scala 117:10]
  wire  _GEN_2639; // @[Execute.scala 117:10]
  wire  _GEN_2640; // @[Execute.scala 117:10]
  wire  _GEN_2641; // @[Execute.scala 117:10]
  wire  _GEN_2642; // @[Execute.scala 117:10]
  wire  _GEN_2643; // @[Execute.scala 117:10]
  wire  _GEN_2644; // @[Execute.scala 117:10]
  wire  _GEN_2645; // @[Execute.scala 117:10]
  wire  _GEN_2646; // @[Execute.scala 117:10]
  wire  _GEN_2647; // @[Execute.scala 117:10]
  wire  _GEN_2648; // @[Execute.scala 117:10]
  wire  _GEN_2649; // @[Execute.scala 117:10]
  wire  _GEN_2650; // @[Execute.scala 117:10]
  wire  _GEN_2651; // @[Execute.scala 117:10]
  wire  _GEN_2652; // @[Execute.scala 117:10]
  wire  _GEN_2653; // @[Execute.scala 117:10]
  wire  _GEN_2654; // @[Execute.scala 117:10]
  wire  _GEN_2655; // @[Execute.scala 117:10]
  wire  _GEN_2656; // @[Execute.scala 117:10]
  wire  _GEN_2657; // @[Execute.scala 117:10]
  wire  _GEN_2658; // @[Execute.scala 117:10]
  wire  _GEN_2659; // @[Execute.scala 117:10]
  wire  _GEN_2660; // @[Execute.scala 117:10]
  wire  _GEN_2661; // @[Execute.scala 117:10]
  wire  _GEN_2662; // @[Execute.scala 117:10]
  wire  _GEN_2663; // @[Execute.scala 117:10]
  wire  _GEN_2664; // @[Execute.scala 117:10]
  wire  _GEN_2665; // @[Execute.scala 117:10]
  wire  _GEN_2666; // @[Execute.scala 117:10]
  wire  _GEN_2667; // @[Execute.scala 117:10]
  wire  _GEN_2668; // @[Execute.scala 117:10]
  wire  _GEN_2669; // @[Execute.scala 117:10]
  wire  _GEN_2670; // @[Execute.scala 117:10]
  wire  _GEN_2671; // @[Execute.scala 117:10]
  wire  _GEN_2672; // @[Execute.scala 117:10]
  wire  _GEN_2673; // @[Execute.scala 117:10]
  wire  _GEN_2674; // @[Execute.scala 117:10]
  wire  _GEN_2675; // @[Execute.scala 117:10]
  wire  _GEN_2676; // @[Execute.scala 117:10]
  wire  _GEN_2677; // @[Execute.scala 117:10]
  wire  _GEN_2678; // @[Execute.scala 117:10]
  wire  _GEN_2679; // @[Execute.scala 117:10]
  wire  _GEN_2680; // @[Execute.scala 117:10]
  wire  _GEN_2681; // @[Execute.scala 117:10]
  wire  _GEN_2682; // @[Execute.scala 117:10]
  wire  _GEN_2683; // @[Execute.scala 117:10]
  wire  _GEN_2684; // @[Execute.scala 117:10]
  wire  _GEN_2685; // @[Execute.scala 117:10]
  wire  _GEN_2686; // @[Execute.scala 117:10]
  wire  _GEN_2687; // @[Execute.scala 117:10]
  wire  _GEN_2688; // @[Execute.scala 117:10]
  wire  _GEN_2689; // @[Execute.scala 117:10]
  wire  _T_291; // @[Execute.scala 117:10]
  wire  _T_292; // @[Execute.scala 117:15]
  wire [5:0] _T_294; // @[Execute.scala 117:37]
  wire [5:0] _T_298; // @[Execute.scala 117:60]
  wire  _GEN_2691; // @[Execute.scala 117:10]
  wire  _GEN_2692; // @[Execute.scala 117:10]
  wire  _GEN_2693; // @[Execute.scala 117:10]
  wire  _GEN_2694; // @[Execute.scala 117:10]
  wire  _GEN_2695; // @[Execute.scala 117:10]
  wire  _GEN_2696; // @[Execute.scala 117:10]
  wire  _GEN_2697; // @[Execute.scala 117:10]
  wire  _GEN_2698; // @[Execute.scala 117:10]
  wire  _GEN_2699; // @[Execute.scala 117:10]
  wire  _GEN_2700; // @[Execute.scala 117:10]
  wire  _GEN_2701; // @[Execute.scala 117:10]
  wire  _GEN_2702; // @[Execute.scala 117:10]
  wire  _GEN_2703; // @[Execute.scala 117:10]
  wire  _GEN_2704; // @[Execute.scala 117:10]
  wire  _GEN_2705; // @[Execute.scala 117:10]
  wire  _GEN_2706; // @[Execute.scala 117:10]
  wire  _GEN_2707; // @[Execute.scala 117:10]
  wire  _GEN_2708; // @[Execute.scala 117:10]
  wire  _GEN_2709; // @[Execute.scala 117:10]
  wire  _GEN_2710; // @[Execute.scala 117:10]
  wire  _GEN_2711; // @[Execute.scala 117:10]
  wire  _GEN_2712; // @[Execute.scala 117:10]
  wire  _GEN_2713; // @[Execute.scala 117:10]
  wire  _GEN_2714; // @[Execute.scala 117:10]
  wire  _GEN_2715; // @[Execute.scala 117:10]
  wire  _GEN_2716; // @[Execute.scala 117:10]
  wire  _GEN_2717; // @[Execute.scala 117:10]
  wire  _GEN_2718; // @[Execute.scala 117:10]
  wire  _GEN_2719; // @[Execute.scala 117:10]
  wire  _GEN_2720; // @[Execute.scala 117:10]
  wire  _GEN_2721; // @[Execute.scala 117:10]
  wire  _GEN_2722; // @[Execute.scala 117:10]
  wire  _GEN_2723; // @[Execute.scala 117:10]
  wire  _GEN_2724; // @[Execute.scala 117:10]
  wire  _GEN_2725; // @[Execute.scala 117:10]
  wire  _GEN_2726; // @[Execute.scala 117:10]
  wire  _GEN_2727; // @[Execute.scala 117:10]
  wire  _GEN_2728; // @[Execute.scala 117:10]
  wire  _GEN_2729; // @[Execute.scala 117:10]
  wire  _GEN_2730; // @[Execute.scala 117:10]
  wire  _GEN_2731; // @[Execute.scala 117:10]
  wire  _GEN_2732; // @[Execute.scala 117:10]
  wire  _GEN_2733; // @[Execute.scala 117:10]
  wire  _GEN_2734; // @[Execute.scala 117:10]
  wire  _GEN_2735; // @[Execute.scala 117:10]
  wire  _GEN_2736; // @[Execute.scala 117:10]
  wire  _GEN_2737; // @[Execute.scala 117:10]
  wire  _GEN_2738; // @[Execute.scala 117:10]
  wire  _GEN_2739; // @[Execute.scala 117:10]
  wire  _GEN_2740; // @[Execute.scala 117:10]
  wire  _GEN_2741; // @[Execute.scala 117:10]
  wire  _GEN_2742; // @[Execute.scala 117:10]
  wire  _GEN_2743; // @[Execute.scala 117:10]
  wire  _GEN_2744; // @[Execute.scala 117:10]
  wire  _GEN_2745; // @[Execute.scala 117:10]
  wire  _GEN_2746; // @[Execute.scala 117:10]
  wire  _GEN_2747; // @[Execute.scala 117:10]
  wire  _GEN_2748; // @[Execute.scala 117:10]
  wire  _GEN_2749; // @[Execute.scala 117:10]
  wire  _GEN_2750; // @[Execute.scala 117:10]
  wire  _GEN_2751; // @[Execute.scala 117:10]
  wire  _GEN_2752; // @[Execute.scala 117:10]
  wire  _GEN_2753; // @[Execute.scala 117:10]
  wire  _GEN_2755; // @[Execute.scala 117:10]
  wire  _GEN_2756; // @[Execute.scala 117:10]
  wire  _GEN_2757; // @[Execute.scala 117:10]
  wire  _GEN_2758; // @[Execute.scala 117:10]
  wire  _GEN_2759; // @[Execute.scala 117:10]
  wire  _GEN_2760; // @[Execute.scala 117:10]
  wire  _GEN_2761; // @[Execute.scala 117:10]
  wire  _GEN_2762; // @[Execute.scala 117:10]
  wire  _GEN_2763; // @[Execute.scala 117:10]
  wire  _GEN_2764; // @[Execute.scala 117:10]
  wire  _GEN_2765; // @[Execute.scala 117:10]
  wire  _GEN_2766; // @[Execute.scala 117:10]
  wire  _GEN_2767; // @[Execute.scala 117:10]
  wire  _GEN_2768; // @[Execute.scala 117:10]
  wire  _GEN_2769; // @[Execute.scala 117:10]
  wire  _GEN_2770; // @[Execute.scala 117:10]
  wire  _GEN_2771; // @[Execute.scala 117:10]
  wire  _GEN_2772; // @[Execute.scala 117:10]
  wire  _GEN_2773; // @[Execute.scala 117:10]
  wire  _GEN_2774; // @[Execute.scala 117:10]
  wire  _GEN_2775; // @[Execute.scala 117:10]
  wire  _GEN_2776; // @[Execute.scala 117:10]
  wire  _GEN_2777; // @[Execute.scala 117:10]
  wire  _GEN_2778; // @[Execute.scala 117:10]
  wire  _GEN_2779; // @[Execute.scala 117:10]
  wire  _GEN_2780; // @[Execute.scala 117:10]
  wire  _GEN_2781; // @[Execute.scala 117:10]
  wire  _GEN_2782; // @[Execute.scala 117:10]
  wire  _GEN_2783; // @[Execute.scala 117:10]
  wire  _GEN_2784; // @[Execute.scala 117:10]
  wire  _GEN_2785; // @[Execute.scala 117:10]
  wire  _GEN_2786; // @[Execute.scala 117:10]
  wire  _GEN_2787; // @[Execute.scala 117:10]
  wire  _GEN_2788; // @[Execute.scala 117:10]
  wire  _GEN_2789; // @[Execute.scala 117:10]
  wire  _GEN_2790; // @[Execute.scala 117:10]
  wire  _GEN_2791; // @[Execute.scala 117:10]
  wire  _GEN_2792; // @[Execute.scala 117:10]
  wire  _GEN_2793; // @[Execute.scala 117:10]
  wire  _GEN_2794; // @[Execute.scala 117:10]
  wire  _GEN_2795; // @[Execute.scala 117:10]
  wire  _GEN_2796; // @[Execute.scala 117:10]
  wire  _GEN_2797; // @[Execute.scala 117:10]
  wire  _GEN_2798; // @[Execute.scala 117:10]
  wire  _GEN_2799; // @[Execute.scala 117:10]
  wire  _GEN_2800; // @[Execute.scala 117:10]
  wire  _GEN_2801; // @[Execute.scala 117:10]
  wire  _GEN_2802; // @[Execute.scala 117:10]
  wire  _GEN_2803; // @[Execute.scala 117:10]
  wire  _GEN_2804; // @[Execute.scala 117:10]
  wire  _GEN_2805; // @[Execute.scala 117:10]
  wire  _GEN_2806; // @[Execute.scala 117:10]
  wire  _GEN_2807; // @[Execute.scala 117:10]
  wire  _GEN_2808; // @[Execute.scala 117:10]
  wire  _GEN_2809; // @[Execute.scala 117:10]
  wire  _GEN_2810; // @[Execute.scala 117:10]
  wire  _GEN_2811; // @[Execute.scala 117:10]
  wire  _GEN_2812; // @[Execute.scala 117:10]
  wire  _GEN_2813; // @[Execute.scala 117:10]
  wire  _GEN_2814; // @[Execute.scala 117:10]
  wire  _GEN_2815; // @[Execute.scala 117:10]
  wire  _GEN_2816; // @[Execute.scala 117:10]
  wire  _GEN_2817; // @[Execute.scala 117:10]
  wire  _T_301; // @[Execute.scala 117:10]
  wire  _T_302; // @[Execute.scala 117:15]
  wire [5:0] _T_304; // @[Execute.scala 117:37]
  wire [5:0] _T_308; // @[Execute.scala 117:60]
  wire  _GEN_2819; // @[Execute.scala 117:10]
  wire  _GEN_2820; // @[Execute.scala 117:10]
  wire  _GEN_2821; // @[Execute.scala 117:10]
  wire  _GEN_2822; // @[Execute.scala 117:10]
  wire  _GEN_2823; // @[Execute.scala 117:10]
  wire  _GEN_2824; // @[Execute.scala 117:10]
  wire  _GEN_2825; // @[Execute.scala 117:10]
  wire  _GEN_2826; // @[Execute.scala 117:10]
  wire  _GEN_2827; // @[Execute.scala 117:10]
  wire  _GEN_2828; // @[Execute.scala 117:10]
  wire  _GEN_2829; // @[Execute.scala 117:10]
  wire  _GEN_2830; // @[Execute.scala 117:10]
  wire  _GEN_2831; // @[Execute.scala 117:10]
  wire  _GEN_2832; // @[Execute.scala 117:10]
  wire  _GEN_2833; // @[Execute.scala 117:10]
  wire  _GEN_2834; // @[Execute.scala 117:10]
  wire  _GEN_2835; // @[Execute.scala 117:10]
  wire  _GEN_2836; // @[Execute.scala 117:10]
  wire  _GEN_2837; // @[Execute.scala 117:10]
  wire  _GEN_2838; // @[Execute.scala 117:10]
  wire  _GEN_2839; // @[Execute.scala 117:10]
  wire  _GEN_2840; // @[Execute.scala 117:10]
  wire  _GEN_2841; // @[Execute.scala 117:10]
  wire  _GEN_2842; // @[Execute.scala 117:10]
  wire  _GEN_2843; // @[Execute.scala 117:10]
  wire  _GEN_2844; // @[Execute.scala 117:10]
  wire  _GEN_2845; // @[Execute.scala 117:10]
  wire  _GEN_2846; // @[Execute.scala 117:10]
  wire  _GEN_2847; // @[Execute.scala 117:10]
  wire  _GEN_2848; // @[Execute.scala 117:10]
  wire  _GEN_2849; // @[Execute.scala 117:10]
  wire  _GEN_2850; // @[Execute.scala 117:10]
  wire  _GEN_2851; // @[Execute.scala 117:10]
  wire  _GEN_2852; // @[Execute.scala 117:10]
  wire  _GEN_2853; // @[Execute.scala 117:10]
  wire  _GEN_2854; // @[Execute.scala 117:10]
  wire  _GEN_2855; // @[Execute.scala 117:10]
  wire  _GEN_2856; // @[Execute.scala 117:10]
  wire  _GEN_2857; // @[Execute.scala 117:10]
  wire  _GEN_2858; // @[Execute.scala 117:10]
  wire  _GEN_2859; // @[Execute.scala 117:10]
  wire  _GEN_2860; // @[Execute.scala 117:10]
  wire  _GEN_2861; // @[Execute.scala 117:10]
  wire  _GEN_2862; // @[Execute.scala 117:10]
  wire  _GEN_2863; // @[Execute.scala 117:10]
  wire  _GEN_2864; // @[Execute.scala 117:10]
  wire  _GEN_2865; // @[Execute.scala 117:10]
  wire  _GEN_2866; // @[Execute.scala 117:10]
  wire  _GEN_2867; // @[Execute.scala 117:10]
  wire  _GEN_2868; // @[Execute.scala 117:10]
  wire  _GEN_2869; // @[Execute.scala 117:10]
  wire  _GEN_2870; // @[Execute.scala 117:10]
  wire  _GEN_2871; // @[Execute.scala 117:10]
  wire  _GEN_2872; // @[Execute.scala 117:10]
  wire  _GEN_2873; // @[Execute.scala 117:10]
  wire  _GEN_2874; // @[Execute.scala 117:10]
  wire  _GEN_2875; // @[Execute.scala 117:10]
  wire  _GEN_2876; // @[Execute.scala 117:10]
  wire  _GEN_2877; // @[Execute.scala 117:10]
  wire  _GEN_2878; // @[Execute.scala 117:10]
  wire  _GEN_2879; // @[Execute.scala 117:10]
  wire  _GEN_2880; // @[Execute.scala 117:10]
  wire  _GEN_2881; // @[Execute.scala 117:10]
  wire  _GEN_2883; // @[Execute.scala 117:10]
  wire  _GEN_2884; // @[Execute.scala 117:10]
  wire  _GEN_2885; // @[Execute.scala 117:10]
  wire  _GEN_2886; // @[Execute.scala 117:10]
  wire  _GEN_2887; // @[Execute.scala 117:10]
  wire  _GEN_2888; // @[Execute.scala 117:10]
  wire  _GEN_2889; // @[Execute.scala 117:10]
  wire  _GEN_2890; // @[Execute.scala 117:10]
  wire  _GEN_2891; // @[Execute.scala 117:10]
  wire  _GEN_2892; // @[Execute.scala 117:10]
  wire  _GEN_2893; // @[Execute.scala 117:10]
  wire  _GEN_2894; // @[Execute.scala 117:10]
  wire  _GEN_2895; // @[Execute.scala 117:10]
  wire  _GEN_2896; // @[Execute.scala 117:10]
  wire  _GEN_2897; // @[Execute.scala 117:10]
  wire  _GEN_2898; // @[Execute.scala 117:10]
  wire  _GEN_2899; // @[Execute.scala 117:10]
  wire  _GEN_2900; // @[Execute.scala 117:10]
  wire  _GEN_2901; // @[Execute.scala 117:10]
  wire  _GEN_2902; // @[Execute.scala 117:10]
  wire  _GEN_2903; // @[Execute.scala 117:10]
  wire  _GEN_2904; // @[Execute.scala 117:10]
  wire  _GEN_2905; // @[Execute.scala 117:10]
  wire  _GEN_2906; // @[Execute.scala 117:10]
  wire  _GEN_2907; // @[Execute.scala 117:10]
  wire  _GEN_2908; // @[Execute.scala 117:10]
  wire  _GEN_2909; // @[Execute.scala 117:10]
  wire  _GEN_2910; // @[Execute.scala 117:10]
  wire  _GEN_2911; // @[Execute.scala 117:10]
  wire  _GEN_2912; // @[Execute.scala 117:10]
  wire  _GEN_2913; // @[Execute.scala 117:10]
  wire  _GEN_2914; // @[Execute.scala 117:10]
  wire  _GEN_2915; // @[Execute.scala 117:10]
  wire  _GEN_2916; // @[Execute.scala 117:10]
  wire  _GEN_2917; // @[Execute.scala 117:10]
  wire  _GEN_2918; // @[Execute.scala 117:10]
  wire  _GEN_2919; // @[Execute.scala 117:10]
  wire  _GEN_2920; // @[Execute.scala 117:10]
  wire  _GEN_2921; // @[Execute.scala 117:10]
  wire  _GEN_2922; // @[Execute.scala 117:10]
  wire  _GEN_2923; // @[Execute.scala 117:10]
  wire  _GEN_2924; // @[Execute.scala 117:10]
  wire  _GEN_2925; // @[Execute.scala 117:10]
  wire  _GEN_2926; // @[Execute.scala 117:10]
  wire  _GEN_2927; // @[Execute.scala 117:10]
  wire  _GEN_2928; // @[Execute.scala 117:10]
  wire  _GEN_2929; // @[Execute.scala 117:10]
  wire  _GEN_2930; // @[Execute.scala 117:10]
  wire  _GEN_2931; // @[Execute.scala 117:10]
  wire  _GEN_2932; // @[Execute.scala 117:10]
  wire  _GEN_2933; // @[Execute.scala 117:10]
  wire  _GEN_2934; // @[Execute.scala 117:10]
  wire  _GEN_2935; // @[Execute.scala 117:10]
  wire  _GEN_2936; // @[Execute.scala 117:10]
  wire  _GEN_2937; // @[Execute.scala 117:10]
  wire  _GEN_2938; // @[Execute.scala 117:10]
  wire  _GEN_2939; // @[Execute.scala 117:10]
  wire  _GEN_2940; // @[Execute.scala 117:10]
  wire  _GEN_2941; // @[Execute.scala 117:10]
  wire  _GEN_2942; // @[Execute.scala 117:10]
  wire  _GEN_2943; // @[Execute.scala 117:10]
  wire  _GEN_2944; // @[Execute.scala 117:10]
  wire  _GEN_2945; // @[Execute.scala 117:10]
  wire  _T_311; // @[Execute.scala 117:10]
  wire  _T_312; // @[Execute.scala 117:15]
  wire [5:0] _T_314; // @[Execute.scala 117:37]
  wire [5:0] _T_318; // @[Execute.scala 117:60]
  wire  _GEN_2947; // @[Execute.scala 117:10]
  wire  _GEN_2948; // @[Execute.scala 117:10]
  wire  _GEN_2949; // @[Execute.scala 117:10]
  wire  _GEN_2950; // @[Execute.scala 117:10]
  wire  _GEN_2951; // @[Execute.scala 117:10]
  wire  _GEN_2952; // @[Execute.scala 117:10]
  wire  _GEN_2953; // @[Execute.scala 117:10]
  wire  _GEN_2954; // @[Execute.scala 117:10]
  wire  _GEN_2955; // @[Execute.scala 117:10]
  wire  _GEN_2956; // @[Execute.scala 117:10]
  wire  _GEN_2957; // @[Execute.scala 117:10]
  wire  _GEN_2958; // @[Execute.scala 117:10]
  wire  _GEN_2959; // @[Execute.scala 117:10]
  wire  _GEN_2960; // @[Execute.scala 117:10]
  wire  _GEN_2961; // @[Execute.scala 117:10]
  wire  _GEN_2962; // @[Execute.scala 117:10]
  wire  _GEN_2963; // @[Execute.scala 117:10]
  wire  _GEN_2964; // @[Execute.scala 117:10]
  wire  _GEN_2965; // @[Execute.scala 117:10]
  wire  _GEN_2966; // @[Execute.scala 117:10]
  wire  _GEN_2967; // @[Execute.scala 117:10]
  wire  _GEN_2968; // @[Execute.scala 117:10]
  wire  _GEN_2969; // @[Execute.scala 117:10]
  wire  _GEN_2970; // @[Execute.scala 117:10]
  wire  _GEN_2971; // @[Execute.scala 117:10]
  wire  _GEN_2972; // @[Execute.scala 117:10]
  wire  _GEN_2973; // @[Execute.scala 117:10]
  wire  _GEN_2974; // @[Execute.scala 117:10]
  wire  _GEN_2975; // @[Execute.scala 117:10]
  wire  _GEN_2976; // @[Execute.scala 117:10]
  wire  _GEN_2977; // @[Execute.scala 117:10]
  wire  _GEN_2978; // @[Execute.scala 117:10]
  wire  _GEN_2979; // @[Execute.scala 117:10]
  wire  _GEN_2980; // @[Execute.scala 117:10]
  wire  _GEN_2981; // @[Execute.scala 117:10]
  wire  _GEN_2982; // @[Execute.scala 117:10]
  wire  _GEN_2983; // @[Execute.scala 117:10]
  wire  _GEN_2984; // @[Execute.scala 117:10]
  wire  _GEN_2985; // @[Execute.scala 117:10]
  wire  _GEN_2986; // @[Execute.scala 117:10]
  wire  _GEN_2987; // @[Execute.scala 117:10]
  wire  _GEN_2988; // @[Execute.scala 117:10]
  wire  _GEN_2989; // @[Execute.scala 117:10]
  wire  _GEN_2990; // @[Execute.scala 117:10]
  wire  _GEN_2991; // @[Execute.scala 117:10]
  wire  _GEN_2992; // @[Execute.scala 117:10]
  wire  _GEN_2993; // @[Execute.scala 117:10]
  wire  _GEN_2994; // @[Execute.scala 117:10]
  wire  _GEN_2995; // @[Execute.scala 117:10]
  wire  _GEN_2996; // @[Execute.scala 117:10]
  wire  _GEN_2997; // @[Execute.scala 117:10]
  wire  _GEN_2998; // @[Execute.scala 117:10]
  wire  _GEN_2999; // @[Execute.scala 117:10]
  wire  _GEN_3000; // @[Execute.scala 117:10]
  wire  _GEN_3001; // @[Execute.scala 117:10]
  wire  _GEN_3002; // @[Execute.scala 117:10]
  wire  _GEN_3003; // @[Execute.scala 117:10]
  wire  _GEN_3004; // @[Execute.scala 117:10]
  wire  _GEN_3005; // @[Execute.scala 117:10]
  wire  _GEN_3006; // @[Execute.scala 117:10]
  wire  _GEN_3007; // @[Execute.scala 117:10]
  wire  _GEN_3008; // @[Execute.scala 117:10]
  wire  _GEN_3009; // @[Execute.scala 117:10]
  wire  _GEN_3011; // @[Execute.scala 117:10]
  wire  _GEN_3012; // @[Execute.scala 117:10]
  wire  _GEN_3013; // @[Execute.scala 117:10]
  wire  _GEN_3014; // @[Execute.scala 117:10]
  wire  _GEN_3015; // @[Execute.scala 117:10]
  wire  _GEN_3016; // @[Execute.scala 117:10]
  wire  _GEN_3017; // @[Execute.scala 117:10]
  wire  _GEN_3018; // @[Execute.scala 117:10]
  wire  _GEN_3019; // @[Execute.scala 117:10]
  wire  _GEN_3020; // @[Execute.scala 117:10]
  wire  _GEN_3021; // @[Execute.scala 117:10]
  wire  _GEN_3022; // @[Execute.scala 117:10]
  wire  _GEN_3023; // @[Execute.scala 117:10]
  wire  _GEN_3024; // @[Execute.scala 117:10]
  wire  _GEN_3025; // @[Execute.scala 117:10]
  wire  _GEN_3026; // @[Execute.scala 117:10]
  wire  _GEN_3027; // @[Execute.scala 117:10]
  wire  _GEN_3028; // @[Execute.scala 117:10]
  wire  _GEN_3029; // @[Execute.scala 117:10]
  wire  _GEN_3030; // @[Execute.scala 117:10]
  wire  _GEN_3031; // @[Execute.scala 117:10]
  wire  _GEN_3032; // @[Execute.scala 117:10]
  wire  _GEN_3033; // @[Execute.scala 117:10]
  wire  _GEN_3034; // @[Execute.scala 117:10]
  wire  _GEN_3035; // @[Execute.scala 117:10]
  wire  _GEN_3036; // @[Execute.scala 117:10]
  wire  _GEN_3037; // @[Execute.scala 117:10]
  wire  _GEN_3038; // @[Execute.scala 117:10]
  wire  _GEN_3039; // @[Execute.scala 117:10]
  wire  _GEN_3040; // @[Execute.scala 117:10]
  wire  _GEN_3041; // @[Execute.scala 117:10]
  wire  _GEN_3042; // @[Execute.scala 117:10]
  wire  _GEN_3043; // @[Execute.scala 117:10]
  wire  _GEN_3044; // @[Execute.scala 117:10]
  wire  _GEN_3045; // @[Execute.scala 117:10]
  wire  _GEN_3046; // @[Execute.scala 117:10]
  wire  _GEN_3047; // @[Execute.scala 117:10]
  wire  _GEN_3048; // @[Execute.scala 117:10]
  wire  _GEN_3049; // @[Execute.scala 117:10]
  wire  _GEN_3050; // @[Execute.scala 117:10]
  wire  _GEN_3051; // @[Execute.scala 117:10]
  wire  _GEN_3052; // @[Execute.scala 117:10]
  wire  _GEN_3053; // @[Execute.scala 117:10]
  wire  _GEN_3054; // @[Execute.scala 117:10]
  wire  _GEN_3055; // @[Execute.scala 117:10]
  wire  _GEN_3056; // @[Execute.scala 117:10]
  wire  _GEN_3057; // @[Execute.scala 117:10]
  wire  _GEN_3058; // @[Execute.scala 117:10]
  wire  _GEN_3059; // @[Execute.scala 117:10]
  wire  _GEN_3060; // @[Execute.scala 117:10]
  wire  _GEN_3061; // @[Execute.scala 117:10]
  wire  _GEN_3062; // @[Execute.scala 117:10]
  wire  _GEN_3063; // @[Execute.scala 117:10]
  wire  _GEN_3064; // @[Execute.scala 117:10]
  wire  _GEN_3065; // @[Execute.scala 117:10]
  wire  _GEN_3066; // @[Execute.scala 117:10]
  wire  _GEN_3067; // @[Execute.scala 117:10]
  wire  _GEN_3068; // @[Execute.scala 117:10]
  wire  _GEN_3069; // @[Execute.scala 117:10]
  wire  _GEN_3070; // @[Execute.scala 117:10]
  wire  _GEN_3071; // @[Execute.scala 117:10]
  wire  _GEN_3072; // @[Execute.scala 117:10]
  wire  _GEN_3073; // @[Execute.scala 117:10]
  wire  _T_321; // @[Execute.scala 117:10]
  wire  _T_322; // @[Execute.scala 117:15]
  wire [5:0] _T_324; // @[Execute.scala 117:37]
  wire [5:0] _T_328; // @[Execute.scala 117:60]
  wire  _GEN_3075; // @[Execute.scala 117:10]
  wire  _GEN_3076; // @[Execute.scala 117:10]
  wire  _GEN_3077; // @[Execute.scala 117:10]
  wire  _GEN_3078; // @[Execute.scala 117:10]
  wire  _GEN_3079; // @[Execute.scala 117:10]
  wire  _GEN_3080; // @[Execute.scala 117:10]
  wire  _GEN_3081; // @[Execute.scala 117:10]
  wire  _GEN_3082; // @[Execute.scala 117:10]
  wire  _GEN_3083; // @[Execute.scala 117:10]
  wire  _GEN_3084; // @[Execute.scala 117:10]
  wire  _GEN_3085; // @[Execute.scala 117:10]
  wire  _GEN_3086; // @[Execute.scala 117:10]
  wire  _GEN_3087; // @[Execute.scala 117:10]
  wire  _GEN_3088; // @[Execute.scala 117:10]
  wire  _GEN_3089; // @[Execute.scala 117:10]
  wire  _GEN_3090; // @[Execute.scala 117:10]
  wire  _GEN_3091; // @[Execute.scala 117:10]
  wire  _GEN_3092; // @[Execute.scala 117:10]
  wire  _GEN_3093; // @[Execute.scala 117:10]
  wire  _GEN_3094; // @[Execute.scala 117:10]
  wire  _GEN_3095; // @[Execute.scala 117:10]
  wire  _GEN_3096; // @[Execute.scala 117:10]
  wire  _GEN_3097; // @[Execute.scala 117:10]
  wire  _GEN_3098; // @[Execute.scala 117:10]
  wire  _GEN_3099; // @[Execute.scala 117:10]
  wire  _GEN_3100; // @[Execute.scala 117:10]
  wire  _GEN_3101; // @[Execute.scala 117:10]
  wire  _GEN_3102; // @[Execute.scala 117:10]
  wire  _GEN_3103; // @[Execute.scala 117:10]
  wire  _GEN_3104; // @[Execute.scala 117:10]
  wire  _GEN_3105; // @[Execute.scala 117:10]
  wire  _GEN_3106; // @[Execute.scala 117:10]
  wire  _GEN_3107; // @[Execute.scala 117:10]
  wire  _GEN_3108; // @[Execute.scala 117:10]
  wire  _GEN_3109; // @[Execute.scala 117:10]
  wire  _GEN_3110; // @[Execute.scala 117:10]
  wire  _GEN_3111; // @[Execute.scala 117:10]
  wire  _GEN_3112; // @[Execute.scala 117:10]
  wire  _GEN_3113; // @[Execute.scala 117:10]
  wire  _GEN_3114; // @[Execute.scala 117:10]
  wire  _GEN_3115; // @[Execute.scala 117:10]
  wire  _GEN_3116; // @[Execute.scala 117:10]
  wire  _GEN_3117; // @[Execute.scala 117:10]
  wire  _GEN_3118; // @[Execute.scala 117:10]
  wire  _GEN_3119; // @[Execute.scala 117:10]
  wire  _GEN_3120; // @[Execute.scala 117:10]
  wire  _GEN_3121; // @[Execute.scala 117:10]
  wire  _GEN_3122; // @[Execute.scala 117:10]
  wire  _GEN_3123; // @[Execute.scala 117:10]
  wire  _GEN_3124; // @[Execute.scala 117:10]
  wire  _GEN_3125; // @[Execute.scala 117:10]
  wire  _GEN_3126; // @[Execute.scala 117:10]
  wire  _GEN_3127; // @[Execute.scala 117:10]
  wire  _GEN_3128; // @[Execute.scala 117:10]
  wire  _GEN_3129; // @[Execute.scala 117:10]
  wire  _GEN_3130; // @[Execute.scala 117:10]
  wire  _GEN_3131; // @[Execute.scala 117:10]
  wire  _GEN_3132; // @[Execute.scala 117:10]
  wire  _GEN_3133; // @[Execute.scala 117:10]
  wire  _GEN_3134; // @[Execute.scala 117:10]
  wire  _GEN_3135; // @[Execute.scala 117:10]
  wire  _GEN_3136; // @[Execute.scala 117:10]
  wire  _GEN_3137; // @[Execute.scala 117:10]
  wire  _GEN_3139; // @[Execute.scala 117:10]
  wire  _GEN_3140; // @[Execute.scala 117:10]
  wire  _GEN_3141; // @[Execute.scala 117:10]
  wire  _GEN_3142; // @[Execute.scala 117:10]
  wire  _GEN_3143; // @[Execute.scala 117:10]
  wire  _GEN_3144; // @[Execute.scala 117:10]
  wire  _GEN_3145; // @[Execute.scala 117:10]
  wire  _GEN_3146; // @[Execute.scala 117:10]
  wire  _GEN_3147; // @[Execute.scala 117:10]
  wire  _GEN_3148; // @[Execute.scala 117:10]
  wire  _GEN_3149; // @[Execute.scala 117:10]
  wire  _GEN_3150; // @[Execute.scala 117:10]
  wire  _GEN_3151; // @[Execute.scala 117:10]
  wire  _GEN_3152; // @[Execute.scala 117:10]
  wire  _GEN_3153; // @[Execute.scala 117:10]
  wire  _GEN_3154; // @[Execute.scala 117:10]
  wire  _GEN_3155; // @[Execute.scala 117:10]
  wire  _GEN_3156; // @[Execute.scala 117:10]
  wire  _GEN_3157; // @[Execute.scala 117:10]
  wire  _GEN_3158; // @[Execute.scala 117:10]
  wire  _GEN_3159; // @[Execute.scala 117:10]
  wire  _GEN_3160; // @[Execute.scala 117:10]
  wire  _GEN_3161; // @[Execute.scala 117:10]
  wire  _GEN_3162; // @[Execute.scala 117:10]
  wire  _GEN_3163; // @[Execute.scala 117:10]
  wire  _GEN_3164; // @[Execute.scala 117:10]
  wire  _GEN_3165; // @[Execute.scala 117:10]
  wire  _GEN_3166; // @[Execute.scala 117:10]
  wire  _GEN_3167; // @[Execute.scala 117:10]
  wire  _GEN_3168; // @[Execute.scala 117:10]
  wire  _GEN_3169; // @[Execute.scala 117:10]
  wire  _GEN_3170; // @[Execute.scala 117:10]
  wire  _GEN_3171; // @[Execute.scala 117:10]
  wire  _GEN_3172; // @[Execute.scala 117:10]
  wire  _GEN_3173; // @[Execute.scala 117:10]
  wire  _GEN_3174; // @[Execute.scala 117:10]
  wire  _GEN_3175; // @[Execute.scala 117:10]
  wire  _GEN_3176; // @[Execute.scala 117:10]
  wire  _GEN_3177; // @[Execute.scala 117:10]
  wire  _GEN_3178; // @[Execute.scala 117:10]
  wire  _GEN_3179; // @[Execute.scala 117:10]
  wire  _GEN_3180; // @[Execute.scala 117:10]
  wire  _GEN_3181; // @[Execute.scala 117:10]
  wire  _GEN_3182; // @[Execute.scala 117:10]
  wire  _GEN_3183; // @[Execute.scala 117:10]
  wire  _GEN_3184; // @[Execute.scala 117:10]
  wire  _GEN_3185; // @[Execute.scala 117:10]
  wire  _GEN_3186; // @[Execute.scala 117:10]
  wire  _GEN_3187; // @[Execute.scala 117:10]
  wire  _GEN_3188; // @[Execute.scala 117:10]
  wire  _GEN_3189; // @[Execute.scala 117:10]
  wire  _GEN_3190; // @[Execute.scala 117:10]
  wire  _GEN_3191; // @[Execute.scala 117:10]
  wire  _GEN_3192; // @[Execute.scala 117:10]
  wire  _GEN_3193; // @[Execute.scala 117:10]
  wire  _GEN_3194; // @[Execute.scala 117:10]
  wire  _GEN_3195; // @[Execute.scala 117:10]
  wire  _GEN_3196; // @[Execute.scala 117:10]
  wire  _GEN_3197; // @[Execute.scala 117:10]
  wire  _GEN_3198; // @[Execute.scala 117:10]
  wire  _GEN_3199; // @[Execute.scala 117:10]
  wire  _GEN_3200; // @[Execute.scala 117:10]
  wire  _GEN_3201; // @[Execute.scala 117:10]
  wire  _T_331; // @[Execute.scala 117:10]
  wire  _T_332; // @[Execute.scala 117:15]
  wire [5:0] _T_334; // @[Execute.scala 117:37]
  wire [5:0] _T_338; // @[Execute.scala 117:60]
  wire  _GEN_3203; // @[Execute.scala 117:10]
  wire  _GEN_3204; // @[Execute.scala 117:10]
  wire  _GEN_3205; // @[Execute.scala 117:10]
  wire  _GEN_3206; // @[Execute.scala 117:10]
  wire  _GEN_3207; // @[Execute.scala 117:10]
  wire  _GEN_3208; // @[Execute.scala 117:10]
  wire  _GEN_3209; // @[Execute.scala 117:10]
  wire  _GEN_3210; // @[Execute.scala 117:10]
  wire  _GEN_3211; // @[Execute.scala 117:10]
  wire  _GEN_3212; // @[Execute.scala 117:10]
  wire  _GEN_3213; // @[Execute.scala 117:10]
  wire  _GEN_3214; // @[Execute.scala 117:10]
  wire  _GEN_3215; // @[Execute.scala 117:10]
  wire  _GEN_3216; // @[Execute.scala 117:10]
  wire  _GEN_3217; // @[Execute.scala 117:10]
  wire  _GEN_3218; // @[Execute.scala 117:10]
  wire  _GEN_3219; // @[Execute.scala 117:10]
  wire  _GEN_3220; // @[Execute.scala 117:10]
  wire  _GEN_3221; // @[Execute.scala 117:10]
  wire  _GEN_3222; // @[Execute.scala 117:10]
  wire  _GEN_3223; // @[Execute.scala 117:10]
  wire  _GEN_3224; // @[Execute.scala 117:10]
  wire  _GEN_3225; // @[Execute.scala 117:10]
  wire  _GEN_3226; // @[Execute.scala 117:10]
  wire  _GEN_3227; // @[Execute.scala 117:10]
  wire  _GEN_3228; // @[Execute.scala 117:10]
  wire  _GEN_3229; // @[Execute.scala 117:10]
  wire  _GEN_3230; // @[Execute.scala 117:10]
  wire  _GEN_3231; // @[Execute.scala 117:10]
  wire  _GEN_3232; // @[Execute.scala 117:10]
  wire  _GEN_3233; // @[Execute.scala 117:10]
  wire  _GEN_3234; // @[Execute.scala 117:10]
  wire  _GEN_3235; // @[Execute.scala 117:10]
  wire  _GEN_3236; // @[Execute.scala 117:10]
  wire  _GEN_3237; // @[Execute.scala 117:10]
  wire  _GEN_3238; // @[Execute.scala 117:10]
  wire  _GEN_3239; // @[Execute.scala 117:10]
  wire  _GEN_3240; // @[Execute.scala 117:10]
  wire  _GEN_3241; // @[Execute.scala 117:10]
  wire  _GEN_3242; // @[Execute.scala 117:10]
  wire  _GEN_3243; // @[Execute.scala 117:10]
  wire  _GEN_3244; // @[Execute.scala 117:10]
  wire  _GEN_3245; // @[Execute.scala 117:10]
  wire  _GEN_3246; // @[Execute.scala 117:10]
  wire  _GEN_3247; // @[Execute.scala 117:10]
  wire  _GEN_3248; // @[Execute.scala 117:10]
  wire  _GEN_3249; // @[Execute.scala 117:10]
  wire  _GEN_3250; // @[Execute.scala 117:10]
  wire  _GEN_3251; // @[Execute.scala 117:10]
  wire  _GEN_3252; // @[Execute.scala 117:10]
  wire  _GEN_3253; // @[Execute.scala 117:10]
  wire  _GEN_3254; // @[Execute.scala 117:10]
  wire  _GEN_3255; // @[Execute.scala 117:10]
  wire  _GEN_3256; // @[Execute.scala 117:10]
  wire  _GEN_3257; // @[Execute.scala 117:10]
  wire  _GEN_3258; // @[Execute.scala 117:10]
  wire  _GEN_3259; // @[Execute.scala 117:10]
  wire  _GEN_3260; // @[Execute.scala 117:10]
  wire  _GEN_3261; // @[Execute.scala 117:10]
  wire  _GEN_3262; // @[Execute.scala 117:10]
  wire  _GEN_3263; // @[Execute.scala 117:10]
  wire  _GEN_3264; // @[Execute.scala 117:10]
  wire  _GEN_3265; // @[Execute.scala 117:10]
  wire  _GEN_3267; // @[Execute.scala 117:10]
  wire  _GEN_3268; // @[Execute.scala 117:10]
  wire  _GEN_3269; // @[Execute.scala 117:10]
  wire  _GEN_3270; // @[Execute.scala 117:10]
  wire  _GEN_3271; // @[Execute.scala 117:10]
  wire  _GEN_3272; // @[Execute.scala 117:10]
  wire  _GEN_3273; // @[Execute.scala 117:10]
  wire  _GEN_3274; // @[Execute.scala 117:10]
  wire  _GEN_3275; // @[Execute.scala 117:10]
  wire  _GEN_3276; // @[Execute.scala 117:10]
  wire  _GEN_3277; // @[Execute.scala 117:10]
  wire  _GEN_3278; // @[Execute.scala 117:10]
  wire  _GEN_3279; // @[Execute.scala 117:10]
  wire  _GEN_3280; // @[Execute.scala 117:10]
  wire  _GEN_3281; // @[Execute.scala 117:10]
  wire  _GEN_3282; // @[Execute.scala 117:10]
  wire  _GEN_3283; // @[Execute.scala 117:10]
  wire  _GEN_3284; // @[Execute.scala 117:10]
  wire  _GEN_3285; // @[Execute.scala 117:10]
  wire  _GEN_3286; // @[Execute.scala 117:10]
  wire  _GEN_3287; // @[Execute.scala 117:10]
  wire  _GEN_3288; // @[Execute.scala 117:10]
  wire  _GEN_3289; // @[Execute.scala 117:10]
  wire  _GEN_3290; // @[Execute.scala 117:10]
  wire  _GEN_3291; // @[Execute.scala 117:10]
  wire  _GEN_3292; // @[Execute.scala 117:10]
  wire  _GEN_3293; // @[Execute.scala 117:10]
  wire  _GEN_3294; // @[Execute.scala 117:10]
  wire  _GEN_3295; // @[Execute.scala 117:10]
  wire  _GEN_3296; // @[Execute.scala 117:10]
  wire  _GEN_3297; // @[Execute.scala 117:10]
  wire  _GEN_3298; // @[Execute.scala 117:10]
  wire  _GEN_3299; // @[Execute.scala 117:10]
  wire  _GEN_3300; // @[Execute.scala 117:10]
  wire  _GEN_3301; // @[Execute.scala 117:10]
  wire  _GEN_3302; // @[Execute.scala 117:10]
  wire  _GEN_3303; // @[Execute.scala 117:10]
  wire  _GEN_3304; // @[Execute.scala 117:10]
  wire  _GEN_3305; // @[Execute.scala 117:10]
  wire  _GEN_3306; // @[Execute.scala 117:10]
  wire  _GEN_3307; // @[Execute.scala 117:10]
  wire  _GEN_3308; // @[Execute.scala 117:10]
  wire  _GEN_3309; // @[Execute.scala 117:10]
  wire  _GEN_3310; // @[Execute.scala 117:10]
  wire  _GEN_3311; // @[Execute.scala 117:10]
  wire  _GEN_3312; // @[Execute.scala 117:10]
  wire  _GEN_3313; // @[Execute.scala 117:10]
  wire  _GEN_3314; // @[Execute.scala 117:10]
  wire  _GEN_3315; // @[Execute.scala 117:10]
  wire  _GEN_3316; // @[Execute.scala 117:10]
  wire  _GEN_3317; // @[Execute.scala 117:10]
  wire  _GEN_3318; // @[Execute.scala 117:10]
  wire  _GEN_3319; // @[Execute.scala 117:10]
  wire  _GEN_3320; // @[Execute.scala 117:10]
  wire  _GEN_3321; // @[Execute.scala 117:10]
  wire  _GEN_3322; // @[Execute.scala 117:10]
  wire  _GEN_3323; // @[Execute.scala 117:10]
  wire  _GEN_3324; // @[Execute.scala 117:10]
  wire  _GEN_3325; // @[Execute.scala 117:10]
  wire  _GEN_3326; // @[Execute.scala 117:10]
  wire  _GEN_3327; // @[Execute.scala 117:10]
  wire  _GEN_3328; // @[Execute.scala 117:10]
  wire  _GEN_3329; // @[Execute.scala 117:10]
  wire  _T_341; // @[Execute.scala 117:10]
  wire  _T_342; // @[Execute.scala 117:15]
  wire [5:0] _T_344; // @[Execute.scala 117:37]
  wire [5:0] _T_348; // @[Execute.scala 117:60]
  wire  _GEN_3331; // @[Execute.scala 117:10]
  wire  _GEN_3332; // @[Execute.scala 117:10]
  wire  _GEN_3333; // @[Execute.scala 117:10]
  wire  _GEN_3334; // @[Execute.scala 117:10]
  wire  _GEN_3335; // @[Execute.scala 117:10]
  wire  _GEN_3336; // @[Execute.scala 117:10]
  wire  _GEN_3337; // @[Execute.scala 117:10]
  wire  _GEN_3338; // @[Execute.scala 117:10]
  wire  _GEN_3339; // @[Execute.scala 117:10]
  wire  _GEN_3340; // @[Execute.scala 117:10]
  wire  _GEN_3341; // @[Execute.scala 117:10]
  wire  _GEN_3342; // @[Execute.scala 117:10]
  wire  _GEN_3343; // @[Execute.scala 117:10]
  wire  _GEN_3344; // @[Execute.scala 117:10]
  wire  _GEN_3345; // @[Execute.scala 117:10]
  wire  _GEN_3346; // @[Execute.scala 117:10]
  wire  _GEN_3347; // @[Execute.scala 117:10]
  wire  _GEN_3348; // @[Execute.scala 117:10]
  wire  _GEN_3349; // @[Execute.scala 117:10]
  wire  _GEN_3350; // @[Execute.scala 117:10]
  wire  _GEN_3351; // @[Execute.scala 117:10]
  wire  _GEN_3352; // @[Execute.scala 117:10]
  wire  _GEN_3353; // @[Execute.scala 117:10]
  wire  _GEN_3354; // @[Execute.scala 117:10]
  wire  _GEN_3355; // @[Execute.scala 117:10]
  wire  _GEN_3356; // @[Execute.scala 117:10]
  wire  _GEN_3357; // @[Execute.scala 117:10]
  wire  _GEN_3358; // @[Execute.scala 117:10]
  wire  _GEN_3359; // @[Execute.scala 117:10]
  wire  _GEN_3360; // @[Execute.scala 117:10]
  wire  _GEN_3361; // @[Execute.scala 117:10]
  wire  _GEN_3362; // @[Execute.scala 117:10]
  wire  _GEN_3363; // @[Execute.scala 117:10]
  wire  _GEN_3364; // @[Execute.scala 117:10]
  wire  _GEN_3365; // @[Execute.scala 117:10]
  wire  _GEN_3366; // @[Execute.scala 117:10]
  wire  _GEN_3367; // @[Execute.scala 117:10]
  wire  _GEN_3368; // @[Execute.scala 117:10]
  wire  _GEN_3369; // @[Execute.scala 117:10]
  wire  _GEN_3370; // @[Execute.scala 117:10]
  wire  _GEN_3371; // @[Execute.scala 117:10]
  wire  _GEN_3372; // @[Execute.scala 117:10]
  wire  _GEN_3373; // @[Execute.scala 117:10]
  wire  _GEN_3374; // @[Execute.scala 117:10]
  wire  _GEN_3375; // @[Execute.scala 117:10]
  wire  _GEN_3376; // @[Execute.scala 117:10]
  wire  _GEN_3377; // @[Execute.scala 117:10]
  wire  _GEN_3378; // @[Execute.scala 117:10]
  wire  _GEN_3379; // @[Execute.scala 117:10]
  wire  _GEN_3380; // @[Execute.scala 117:10]
  wire  _GEN_3381; // @[Execute.scala 117:10]
  wire  _GEN_3382; // @[Execute.scala 117:10]
  wire  _GEN_3383; // @[Execute.scala 117:10]
  wire  _GEN_3384; // @[Execute.scala 117:10]
  wire  _GEN_3385; // @[Execute.scala 117:10]
  wire  _GEN_3386; // @[Execute.scala 117:10]
  wire  _GEN_3387; // @[Execute.scala 117:10]
  wire  _GEN_3388; // @[Execute.scala 117:10]
  wire  _GEN_3389; // @[Execute.scala 117:10]
  wire  _GEN_3390; // @[Execute.scala 117:10]
  wire  _GEN_3391; // @[Execute.scala 117:10]
  wire  _GEN_3392; // @[Execute.scala 117:10]
  wire  _GEN_3393; // @[Execute.scala 117:10]
  wire  _GEN_3395; // @[Execute.scala 117:10]
  wire  _GEN_3396; // @[Execute.scala 117:10]
  wire  _GEN_3397; // @[Execute.scala 117:10]
  wire  _GEN_3398; // @[Execute.scala 117:10]
  wire  _GEN_3399; // @[Execute.scala 117:10]
  wire  _GEN_3400; // @[Execute.scala 117:10]
  wire  _GEN_3401; // @[Execute.scala 117:10]
  wire  _GEN_3402; // @[Execute.scala 117:10]
  wire  _GEN_3403; // @[Execute.scala 117:10]
  wire  _GEN_3404; // @[Execute.scala 117:10]
  wire  _GEN_3405; // @[Execute.scala 117:10]
  wire  _GEN_3406; // @[Execute.scala 117:10]
  wire  _GEN_3407; // @[Execute.scala 117:10]
  wire  _GEN_3408; // @[Execute.scala 117:10]
  wire  _GEN_3409; // @[Execute.scala 117:10]
  wire  _GEN_3410; // @[Execute.scala 117:10]
  wire  _GEN_3411; // @[Execute.scala 117:10]
  wire  _GEN_3412; // @[Execute.scala 117:10]
  wire  _GEN_3413; // @[Execute.scala 117:10]
  wire  _GEN_3414; // @[Execute.scala 117:10]
  wire  _GEN_3415; // @[Execute.scala 117:10]
  wire  _GEN_3416; // @[Execute.scala 117:10]
  wire  _GEN_3417; // @[Execute.scala 117:10]
  wire  _GEN_3418; // @[Execute.scala 117:10]
  wire  _GEN_3419; // @[Execute.scala 117:10]
  wire  _GEN_3420; // @[Execute.scala 117:10]
  wire  _GEN_3421; // @[Execute.scala 117:10]
  wire  _GEN_3422; // @[Execute.scala 117:10]
  wire  _GEN_3423; // @[Execute.scala 117:10]
  wire  _GEN_3424; // @[Execute.scala 117:10]
  wire  _GEN_3425; // @[Execute.scala 117:10]
  wire  _GEN_3426; // @[Execute.scala 117:10]
  wire  _GEN_3427; // @[Execute.scala 117:10]
  wire  _GEN_3428; // @[Execute.scala 117:10]
  wire  _GEN_3429; // @[Execute.scala 117:10]
  wire  _GEN_3430; // @[Execute.scala 117:10]
  wire  _GEN_3431; // @[Execute.scala 117:10]
  wire  _GEN_3432; // @[Execute.scala 117:10]
  wire  _GEN_3433; // @[Execute.scala 117:10]
  wire  _GEN_3434; // @[Execute.scala 117:10]
  wire  _GEN_3435; // @[Execute.scala 117:10]
  wire  _GEN_3436; // @[Execute.scala 117:10]
  wire  _GEN_3437; // @[Execute.scala 117:10]
  wire  _GEN_3438; // @[Execute.scala 117:10]
  wire  _GEN_3439; // @[Execute.scala 117:10]
  wire  _GEN_3440; // @[Execute.scala 117:10]
  wire  _GEN_3441; // @[Execute.scala 117:10]
  wire  _GEN_3442; // @[Execute.scala 117:10]
  wire  _GEN_3443; // @[Execute.scala 117:10]
  wire  _GEN_3444; // @[Execute.scala 117:10]
  wire  _GEN_3445; // @[Execute.scala 117:10]
  wire  _GEN_3446; // @[Execute.scala 117:10]
  wire  _GEN_3447; // @[Execute.scala 117:10]
  wire  _GEN_3448; // @[Execute.scala 117:10]
  wire  _GEN_3449; // @[Execute.scala 117:10]
  wire  _GEN_3450; // @[Execute.scala 117:10]
  wire  _GEN_3451; // @[Execute.scala 117:10]
  wire  _GEN_3452; // @[Execute.scala 117:10]
  wire  _GEN_3453; // @[Execute.scala 117:10]
  wire  _GEN_3454; // @[Execute.scala 117:10]
  wire  _GEN_3455; // @[Execute.scala 117:10]
  wire  _GEN_3456; // @[Execute.scala 117:10]
  wire  _GEN_3457; // @[Execute.scala 117:10]
  wire  _T_351; // @[Execute.scala 117:10]
  wire  _T_352; // @[Execute.scala 117:15]
  wire [5:0] _T_354; // @[Execute.scala 117:37]
  wire [5:0] _T_358; // @[Execute.scala 117:60]
  wire  _GEN_3459; // @[Execute.scala 117:10]
  wire  _GEN_3460; // @[Execute.scala 117:10]
  wire  _GEN_3461; // @[Execute.scala 117:10]
  wire  _GEN_3462; // @[Execute.scala 117:10]
  wire  _GEN_3463; // @[Execute.scala 117:10]
  wire  _GEN_3464; // @[Execute.scala 117:10]
  wire  _GEN_3465; // @[Execute.scala 117:10]
  wire  _GEN_3466; // @[Execute.scala 117:10]
  wire  _GEN_3467; // @[Execute.scala 117:10]
  wire  _GEN_3468; // @[Execute.scala 117:10]
  wire  _GEN_3469; // @[Execute.scala 117:10]
  wire  _GEN_3470; // @[Execute.scala 117:10]
  wire  _GEN_3471; // @[Execute.scala 117:10]
  wire  _GEN_3472; // @[Execute.scala 117:10]
  wire  _GEN_3473; // @[Execute.scala 117:10]
  wire  _GEN_3474; // @[Execute.scala 117:10]
  wire  _GEN_3475; // @[Execute.scala 117:10]
  wire  _GEN_3476; // @[Execute.scala 117:10]
  wire  _GEN_3477; // @[Execute.scala 117:10]
  wire  _GEN_3478; // @[Execute.scala 117:10]
  wire  _GEN_3479; // @[Execute.scala 117:10]
  wire  _GEN_3480; // @[Execute.scala 117:10]
  wire  _GEN_3481; // @[Execute.scala 117:10]
  wire  _GEN_3482; // @[Execute.scala 117:10]
  wire  _GEN_3483; // @[Execute.scala 117:10]
  wire  _GEN_3484; // @[Execute.scala 117:10]
  wire  _GEN_3485; // @[Execute.scala 117:10]
  wire  _GEN_3486; // @[Execute.scala 117:10]
  wire  _GEN_3487; // @[Execute.scala 117:10]
  wire  _GEN_3488; // @[Execute.scala 117:10]
  wire  _GEN_3489; // @[Execute.scala 117:10]
  wire  _GEN_3490; // @[Execute.scala 117:10]
  wire  _GEN_3491; // @[Execute.scala 117:10]
  wire  _GEN_3492; // @[Execute.scala 117:10]
  wire  _GEN_3493; // @[Execute.scala 117:10]
  wire  _GEN_3494; // @[Execute.scala 117:10]
  wire  _GEN_3495; // @[Execute.scala 117:10]
  wire  _GEN_3496; // @[Execute.scala 117:10]
  wire  _GEN_3497; // @[Execute.scala 117:10]
  wire  _GEN_3498; // @[Execute.scala 117:10]
  wire  _GEN_3499; // @[Execute.scala 117:10]
  wire  _GEN_3500; // @[Execute.scala 117:10]
  wire  _GEN_3501; // @[Execute.scala 117:10]
  wire  _GEN_3502; // @[Execute.scala 117:10]
  wire  _GEN_3503; // @[Execute.scala 117:10]
  wire  _GEN_3504; // @[Execute.scala 117:10]
  wire  _GEN_3505; // @[Execute.scala 117:10]
  wire  _GEN_3506; // @[Execute.scala 117:10]
  wire  _GEN_3507; // @[Execute.scala 117:10]
  wire  _GEN_3508; // @[Execute.scala 117:10]
  wire  _GEN_3509; // @[Execute.scala 117:10]
  wire  _GEN_3510; // @[Execute.scala 117:10]
  wire  _GEN_3511; // @[Execute.scala 117:10]
  wire  _GEN_3512; // @[Execute.scala 117:10]
  wire  _GEN_3513; // @[Execute.scala 117:10]
  wire  _GEN_3514; // @[Execute.scala 117:10]
  wire  _GEN_3515; // @[Execute.scala 117:10]
  wire  _GEN_3516; // @[Execute.scala 117:10]
  wire  _GEN_3517; // @[Execute.scala 117:10]
  wire  _GEN_3518; // @[Execute.scala 117:10]
  wire  _GEN_3519; // @[Execute.scala 117:10]
  wire  _GEN_3520; // @[Execute.scala 117:10]
  wire  _GEN_3521; // @[Execute.scala 117:10]
  wire  _GEN_3523; // @[Execute.scala 117:10]
  wire  _GEN_3524; // @[Execute.scala 117:10]
  wire  _GEN_3525; // @[Execute.scala 117:10]
  wire  _GEN_3526; // @[Execute.scala 117:10]
  wire  _GEN_3527; // @[Execute.scala 117:10]
  wire  _GEN_3528; // @[Execute.scala 117:10]
  wire  _GEN_3529; // @[Execute.scala 117:10]
  wire  _GEN_3530; // @[Execute.scala 117:10]
  wire  _GEN_3531; // @[Execute.scala 117:10]
  wire  _GEN_3532; // @[Execute.scala 117:10]
  wire  _GEN_3533; // @[Execute.scala 117:10]
  wire  _GEN_3534; // @[Execute.scala 117:10]
  wire  _GEN_3535; // @[Execute.scala 117:10]
  wire  _GEN_3536; // @[Execute.scala 117:10]
  wire  _GEN_3537; // @[Execute.scala 117:10]
  wire  _GEN_3538; // @[Execute.scala 117:10]
  wire  _GEN_3539; // @[Execute.scala 117:10]
  wire  _GEN_3540; // @[Execute.scala 117:10]
  wire  _GEN_3541; // @[Execute.scala 117:10]
  wire  _GEN_3542; // @[Execute.scala 117:10]
  wire  _GEN_3543; // @[Execute.scala 117:10]
  wire  _GEN_3544; // @[Execute.scala 117:10]
  wire  _GEN_3545; // @[Execute.scala 117:10]
  wire  _GEN_3546; // @[Execute.scala 117:10]
  wire  _GEN_3547; // @[Execute.scala 117:10]
  wire  _GEN_3548; // @[Execute.scala 117:10]
  wire  _GEN_3549; // @[Execute.scala 117:10]
  wire  _GEN_3550; // @[Execute.scala 117:10]
  wire  _GEN_3551; // @[Execute.scala 117:10]
  wire  _GEN_3552; // @[Execute.scala 117:10]
  wire  _GEN_3553; // @[Execute.scala 117:10]
  wire  _GEN_3554; // @[Execute.scala 117:10]
  wire  _GEN_3555; // @[Execute.scala 117:10]
  wire  _GEN_3556; // @[Execute.scala 117:10]
  wire  _GEN_3557; // @[Execute.scala 117:10]
  wire  _GEN_3558; // @[Execute.scala 117:10]
  wire  _GEN_3559; // @[Execute.scala 117:10]
  wire  _GEN_3560; // @[Execute.scala 117:10]
  wire  _GEN_3561; // @[Execute.scala 117:10]
  wire  _GEN_3562; // @[Execute.scala 117:10]
  wire  _GEN_3563; // @[Execute.scala 117:10]
  wire  _GEN_3564; // @[Execute.scala 117:10]
  wire  _GEN_3565; // @[Execute.scala 117:10]
  wire  _GEN_3566; // @[Execute.scala 117:10]
  wire  _GEN_3567; // @[Execute.scala 117:10]
  wire  _GEN_3568; // @[Execute.scala 117:10]
  wire  _GEN_3569; // @[Execute.scala 117:10]
  wire  _GEN_3570; // @[Execute.scala 117:10]
  wire  _GEN_3571; // @[Execute.scala 117:10]
  wire  _GEN_3572; // @[Execute.scala 117:10]
  wire  _GEN_3573; // @[Execute.scala 117:10]
  wire  _GEN_3574; // @[Execute.scala 117:10]
  wire  _GEN_3575; // @[Execute.scala 117:10]
  wire  _GEN_3576; // @[Execute.scala 117:10]
  wire  _GEN_3577; // @[Execute.scala 117:10]
  wire  _GEN_3578; // @[Execute.scala 117:10]
  wire  _GEN_3579; // @[Execute.scala 117:10]
  wire  _GEN_3580; // @[Execute.scala 117:10]
  wire  _GEN_3581; // @[Execute.scala 117:10]
  wire  _GEN_3582; // @[Execute.scala 117:10]
  wire  _GEN_3583; // @[Execute.scala 117:10]
  wire  _GEN_3584; // @[Execute.scala 117:10]
  wire  _GEN_3585; // @[Execute.scala 117:10]
  wire  _T_361; // @[Execute.scala 117:10]
  wire  _T_362; // @[Execute.scala 117:15]
  wire [5:0] _T_364; // @[Execute.scala 117:37]
  wire [5:0] _T_368; // @[Execute.scala 117:60]
  wire  _GEN_3587; // @[Execute.scala 117:10]
  wire  _GEN_3588; // @[Execute.scala 117:10]
  wire  _GEN_3589; // @[Execute.scala 117:10]
  wire  _GEN_3590; // @[Execute.scala 117:10]
  wire  _GEN_3591; // @[Execute.scala 117:10]
  wire  _GEN_3592; // @[Execute.scala 117:10]
  wire  _GEN_3593; // @[Execute.scala 117:10]
  wire  _GEN_3594; // @[Execute.scala 117:10]
  wire  _GEN_3595; // @[Execute.scala 117:10]
  wire  _GEN_3596; // @[Execute.scala 117:10]
  wire  _GEN_3597; // @[Execute.scala 117:10]
  wire  _GEN_3598; // @[Execute.scala 117:10]
  wire  _GEN_3599; // @[Execute.scala 117:10]
  wire  _GEN_3600; // @[Execute.scala 117:10]
  wire  _GEN_3601; // @[Execute.scala 117:10]
  wire  _GEN_3602; // @[Execute.scala 117:10]
  wire  _GEN_3603; // @[Execute.scala 117:10]
  wire  _GEN_3604; // @[Execute.scala 117:10]
  wire  _GEN_3605; // @[Execute.scala 117:10]
  wire  _GEN_3606; // @[Execute.scala 117:10]
  wire  _GEN_3607; // @[Execute.scala 117:10]
  wire  _GEN_3608; // @[Execute.scala 117:10]
  wire  _GEN_3609; // @[Execute.scala 117:10]
  wire  _GEN_3610; // @[Execute.scala 117:10]
  wire  _GEN_3611; // @[Execute.scala 117:10]
  wire  _GEN_3612; // @[Execute.scala 117:10]
  wire  _GEN_3613; // @[Execute.scala 117:10]
  wire  _GEN_3614; // @[Execute.scala 117:10]
  wire  _GEN_3615; // @[Execute.scala 117:10]
  wire  _GEN_3616; // @[Execute.scala 117:10]
  wire  _GEN_3617; // @[Execute.scala 117:10]
  wire  _GEN_3618; // @[Execute.scala 117:10]
  wire  _GEN_3619; // @[Execute.scala 117:10]
  wire  _GEN_3620; // @[Execute.scala 117:10]
  wire  _GEN_3621; // @[Execute.scala 117:10]
  wire  _GEN_3622; // @[Execute.scala 117:10]
  wire  _GEN_3623; // @[Execute.scala 117:10]
  wire  _GEN_3624; // @[Execute.scala 117:10]
  wire  _GEN_3625; // @[Execute.scala 117:10]
  wire  _GEN_3626; // @[Execute.scala 117:10]
  wire  _GEN_3627; // @[Execute.scala 117:10]
  wire  _GEN_3628; // @[Execute.scala 117:10]
  wire  _GEN_3629; // @[Execute.scala 117:10]
  wire  _GEN_3630; // @[Execute.scala 117:10]
  wire  _GEN_3631; // @[Execute.scala 117:10]
  wire  _GEN_3632; // @[Execute.scala 117:10]
  wire  _GEN_3633; // @[Execute.scala 117:10]
  wire  _GEN_3634; // @[Execute.scala 117:10]
  wire  _GEN_3635; // @[Execute.scala 117:10]
  wire  _GEN_3636; // @[Execute.scala 117:10]
  wire  _GEN_3637; // @[Execute.scala 117:10]
  wire  _GEN_3638; // @[Execute.scala 117:10]
  wire  _GEN_3639; // @[Execute.scala 117:10]
  wire  _GEN_3640; // @[Execute.scala 117:10]
  wire  _GEN_3641; // @[Execute.scala 117:10]
  wire  _GEN_3642; // @[Execute.scala 117:10]
  wire  _GEN_3643; // @[Execute.scala 117:10]
  wire  _GEN_3644; // @[Execute.scala 117:10]
  wire  _GEN_3645; // @[Execute.scala 117:10]
  wire  _GEN_3646; // @[Execute.scala 117:10]
  wire  _GEN_3647; // @[Execute.scala 117:10]
  wire  _GEN_3648; // @[Execute.scala 117:10]
  wire  _GEN_3649; // @[Execute.scala 117:10]
  wire  _GEN_3651; // @[Execute.scala 117:10]
  wire  _GEN_3652; // @[Execute.scala 117:10]
  wire  _GEN_3653; // @[Execute.scala 117:10]
  wire  _GEN_3654; // @[Execute.scala 117:10]
  wire  _GEN_3655; // @[Execute.scala 117:10]
  wire  _GEN_3656; // @[Execute.scala 117:10]
  wire  _GEN_3657; // @[Execute.scala 117:10]
  wire  _GEN_3658; // @[Execute.scala 117:10]
  wire  _GEN_3659; // @[Execute.scala 117:10]
  wire  _GEN_3660; // @[Execute.scala 117:10]
  wire  _GEN_3661; // @[Execute.scala 117:10]
  wire  _GEN_3662; // @[Execute.scala 117:10]
  wire  _GEN_3663; // @[Execute.scala 117:10]
  wire  _GEN_3664; // @[Execute.scala 117:10]
  wire  _GEN_3665; // @[Execute.scala 117:10]
  wire  _GEN_3666; // @[Execute.scala 117:10]
  wire  _GEN_3667; // @[Execute.scala 117:10]
  wire  _GEN_3668; // @[Execute.scala 117:10]
  wire  _GEN_3669; // @[Execute.scala 117:10]
  wire  _GEN_3670; // @[Execute.scala 117:10]
  wire  _GEN_3671; // @[Execute.scala 117:10]
  wire  _GEN_3672; // @[Execute.scala 117:10]
  wire  _GEN_3673; // @[Execute.scala 117:10]
  wire  _GEN_3674; // @[Execute.scala 117:10]
  wire  _GEN_3675; // @[Execute.scala 117:10]
  wire  _GEN_3676; // @[Execute.scala 117:10]
  wire  _GEN_3677; // @[Execute.scala 117:10]
  wire  _GEN_3678; // @[Execute.scala 117:10]
  wire  _GEN_3679; // @[Execute.scala 117:10]
  wire  _GEN_3680; // @[Execute.scala 117:10]
  wire  _GEN_3681; // @[Execute.scala 117:10]
  wire  _GEN_3682; // @[Execute.scala 117:10]
  wire  _GEN_3683; // @[Execute.scala 117:10]
  wire  _GEN_3684; // @[Execute.scala 117:10]
  wire  _GEN_3685; // @[Execute.scala 117:10]
  wire  _GEN_3686; // @[Execute.scala 117:10]
  wire  _GEN_3687; // @[Execute.scala 117:10]
  wire  _GEN_3688; // @[Execute.scala 117:10]
  wire  _GEN_3689; // @[Execute.scala 117:10]
  wire  _GEN_3690; // @[Execute.scala 117:10]
  wire  _GEN_3691; // @[Execute.scala 117:10]
  wire  _GEN_3692; // @[Execute.scala 117:10]
  wire  _GEN_3693; // @[Execute.scala 117:10]
  wire  _GEN_3694; // @[Execute.scala 117:10]
  wire  _GEN_3695; // @[Execute.scala 117:10]
  wire  _GEN_3696; // @[Execute.scala 117:10]
  wire  _GEN_3697; // @[Execute.scala 117:10]
  wire  _GEN_3698; // @[Execute.scala 117:10]
  wire  _GEN_3699; // @[Execute.scala 117:10]
  wire  _GEN_3700; // @[Execute.scala 117:10]
  wire  _GEN_3701; // @[Execute.scala 117:10]
  wire  _GEN_3702; // @[Execute.scala 117:10]
  wire  _GEN_3703; // @[Execute.scala 117:10]
  wire  _GEN_3704; // @[Execute.scala 117:10]
  wire  _GEN_3705; // @[Execute.scala 117:10]
  wire  _GEN_3706; // @[Execute.scala 117:10]
  wire  _GEN_3707; // @[Execute.scala 117:10]
  wire  _GEN_3708; // @[Execute.scala 117:10]
  wire  _GEN_3709; // @[Execute.scala 117:10]
  wire  _GEN_3710; // @[Execute.scala 117:10]
  wire  _GEN_3711; // @[Execute.scala 117:10]
  wire  _GEN_3712; // @[Execute.scala 117:10]
  wire  _GEN_3713; // @[Execute.scala 117:10]
  wire  _T_371; // @[Execute.scala 117:10]
  wire  _T_372; // @[Execute.scala 117:15]
  wire [5:0] _T_374; // @[Execute.scala 117:37]
  wire [5:0] _T_378; // @[Execute.scala 117:60]
  wire  _GEN_3715; // @[Execute.scala 117:10]
  wire  _GEN_3716; // @[Execute.scala 117:10]
  wire  _GEN_3717; // @[Execute.scala 117:10]
  wire  _GEN_3718; // @[Execute.scala 117:10]
  wire  _GEN_3719; // @[Execute.scala 117:10]
  wire  _GEN_3720; // @[Execute.scala 117:10]
  wire  _GEN_3721; // @[Execute.scala 117:10]
  wire  _GEN_3722; // @[Execute.scala 117:10]
  wire  _GEN_3723; // @[Execute.scala 117:10]
  wire  _GEN_3724; // @[Execute.scala 117:10]
  wire  _GEN_3725; // @[Execute.scala 117:10]
  wire  _GEN_3726; // @[Execute.scala 117:10]
  wire  _GEN_3727; // @[Execute.scala 117:10]
  wire  _GEN_3728; // @[Execute.scala 117:10]
  wire  _GEN_3729; // @[Execute.scala 117:10]
  wire  _GEN_3730; // @[Execute.scala 117:10]
  wire  _GEN_3731; // @[Execute.scala 117:10]
  wire  _GEN_3732; // @[Execute.scala 117:10]
  wire  _GEN_3733; // @[Execute.scala 117:10]
  wire  _GEN_3734; // @[Execute.scala 117:10]
  wire  _GEN_3735; // @[Execute.scala 117:10]
  wire  _GEN_3736; // @[Execute.scala 117:10]
  wire  _GEN_3737; // @[Execute.scala 117:10]
  wire  _GEN_3738; // @[Execute.scala 117:10]
  wire  _GEN_3739; // @[Execute.scala 117:10]
  wire  _GEN_3740; // @[Execute.scala 117:10]
  wire  _GEN_3741; // @[Execute.scala 117:10]
  wire  _GEN_3742; // @[Execute.scala 117:10]
  wire  _GEN_3743; // @[Execute.scala 117:10]
  wire  _GEN_3744; // @[Execute.scala 117:10]
  wire  _GEN_3745; // @[Execute.scala 117:10]
  wire  _GEN_3746; // @[Execute.scala 117:10]
  wire  _GEN_3747; // @[Execute.scala 117:10]
  wire  _GEN_3748; // @[Execute.scala 117:10]
  wire  _GEN_3749; // @[Execute.scala 117:10]
  wire  _GEN_3750; // @[Execute.scala 117:10]
  wire  _GEN_3751; // @[Execute.scala 117:10]
  wire  _GEN_3752; // @[Execute.scala 117:10]
  wire  _GEN_3753; // @[Execute.scala 117:10]
  wire  _GEN_3754; // @[Execute.scala 117:10]
  wire  _GEN_3755; // @[Execute.scala 117:10]
  wire  _GEN_3756; // @[Execute.scala 117:10]
  wire  _GEN_3757; // @[Execute.scala 117:10]
  wire  _GEN_3758; // @[Execute.scala 117:10]
  wire  _GEN_3759; // @[Execute.scala 117:10]
  wire  _GEN_3760; // @[Execute.scala 117:10]
  wire  _GEN_3761; // @[Execute.scala 117:10]
  wire  _GEN_3762; // @[Execute.scala 117:10]
  wire  _GEN_3763; // @[Execute.scala 117:10]
  wire  _GEN_3764; // @[Execute.scala 117:10]
  wire  _GEN_3765; // @[Execute.scala 117:10]
  wire  _GEN_3766; // @[Execute.scala 117:10]
  wire  _GEN_3767; // @[Execute.scala 117:10]
  wire  _GEN_3768; // @[Execute.scala 117:10]
  wire  _GEN_3769; // @[Execute.scala 117:10]
  wire  _GEN_3770; // @[Execute.scala 117:10]
  wire  _GEN_3771; // @[Execute.scala 117:10]
  wire  _GEN_3772; // @[Execute.scala 117:10]
  wire  _GEN_3773; // @[Execute.scala 117:10]
  wire  _GEN_3774; // @[Execute.scala 117:10]
  wire  _GEN_3775; // @[Execute.scala 117:10]
  wire  _GEN_3776; // @[Execute.scala 117:10]
  wire  _GEN_3777; // @[Execute.scala 117:10]
  wire  _GEN_3779; // @[Execute.scala 117:10]
  wire  _GEN_3780; // @[Execute.scala 117:10]
  wire  _GEN_3781; // @[Execute.scala 117:10]
  wire  _GEN_3782; // @[Execute.scala 117:10]
  wire  _GEN_3783; // @[Execute.scala 117:10]
  wire  _GEN_3784; // @[Execute.scala 117:10]
  wire  _GEN_3785; // @[Execute.scala 117:10]
  wire  _GEN_3786; // @[Execute.scala 117:10]
  wire  _GEN_3787; // @[Execute.scala 117:10]
  wire  _GEN_3788; // @[Execute.scala 117:10]
  wire  _GEN_3789; // @[Execute.scala 117:10]
  wire  _GEN_3790; // @[Execute.scala 117:10]
  wire  _GEN_3791; // @[Execute.scala 117:10]
  wire  _GEN_3792; // @[Execute.scala 117:10]
  wire  _GEN_3793; // @[Execute.scala 117:10]
  wire  _GEN_3794; // @[Execute.scala 117:10]
  wire  _GEN_3795; // @[Execute.scala 117:10]
  wire  _GEN_3796; // @[Execute.scala 117:10]
  wire  _GEN_3797; // @[Execute.scala 117:10]
  wire  _GEN_3798; // @[Execute.scala 117:10]
  wire  _GEN_3799; // @[Execute.scala 117:10]
  wire  _GEN_3800; // @[Execute.scala 117:10]
  wire  _GEN_3801; // @[Execute.scala 117:10]
  wire  _GEN_3802; // @[Execute.scala 117:10]
  wire  _GEN_3803; // @[Execute.scala 117:10]
  wire  _GEN_3804; // @[Execute.scala 117:10]
  wire  _GEN_3805; // @[Execute.scala 117:10]
  wire  _GEN_3806; // @[Execute.scala 117:10]
  wire  _GEN_3807; // @[Execute.scala 117:10]
  wire  _GEN_3808; // @[Execute.scala 117:10]
  wire  _GEN_3809; // @[Execute.scala 117:10]
  wire  _GEN_3810; // @[Execute.scala 117:10]
  wire  _GEN_3811; // @[Execute.scala 117:10]
  wire  _GEN_3812; // @[Execute.scala 117:10]
  wire  _GEN_3813; // @[Execute.scala 117:10]
  wire  _GEN_3814; // @[Execute.scala 117:10]
  wire  _GEN_3815; // @[Execute.scala 117:10]
  wire  _GEN_3816; // @[Execute.scala 117:10]
  wire  _GEN_3817; // @[Execute.scala 117:10]
  wire  _GEN_3818; // @[Execute.scala 117:10]
  wire  _GEN_3819; // @[Execute.scala 117:10]
  wire  _GEN_3820; // @[Execute.scala 117:10]
  wire  _GEN_3821; // @[Execute.scala 117:10]
  wire  _GEN_3822; // @[Execute.scala 117:10]
  wire  _GEN_3823; // @[Execute.scala 117:10]
  wire  _GEN_3824; // @[Execute.scala 117:10]
  wire  _GEN_3825; // @[Execute.scala 117:10]
  wire  _GEN_3826; // @[Execute.scala 117:10]
  wire  _GEN_3827; // @[Execute.scala 117:10]
  wire  _GEN_3828; // @[Execute.scala 117:10]
  wire  _GEN_3829; // @[Execute.scala 117:10]
  wire  _GEN_3830; // @[Execute.scala 117:10]
  wire  _GEN_3831; // @[Execute.scala 117:10]
  wire  _GEN_3832; // @[Execute.scala 117:10]
  wire  _GEN_3833; // @[Execute.scala 117:10]
  wire  _GEN_3834; // @[Execute.scala 117:10]
  wire  _GEN_3835; // @[Execute.scala 117:10]
  wire  _GEN_3836; // @[Execute.scala 117:10]
  wire  _GEN_3837; // @[Execute.scala 117:10]
  wire  _GEN_3838; // @[Execute.scala 117:10]
  wire  _GEN_3839; // @[Execute.scala 117:10]
  wire  _GEN_3840; // @[Execute.scala 117:10]
  wire  _GEN_3841; // @[Execute.scala 117:10]
  wire  _T_381; // @[Execute.scala 117:10]
  wire  _T_382; // @[Execute.scala 117:15]
  wire [5:0] _T_384; // @[Execute.scala 117:37]
  wire [5:0] _T_388; // @[Execute.scala 117:60]
  wire  _GEN_3843; // @[Execute.scala 117:10]
  wire  _GEN_3844; // @[Execute.scala 117:10]
  wire  _GEN_3845; // @[Execute.scala 117:10]
  wire  _GEN_3846; // @[Execute.scala 117:10]
  wire  _GEN_3847; // @[Execute.scala 117:10]
  wire  _GEN_3848; // @[Execute.scala 117:10]
  wire  _GEN_3849; // @[Execute.scala 117:10]
  wire  _GEN_3850; // @[Execute.scala 117:10]
  wire  _GEN_3851; // @[Execute.scala 117:10]
  wire  _GEN_3852; // @[Execute.scala 117:10]
  wire  _GEN_3853; // @[Execute.scala 117:10]
  wire  _GEN_3854; // @[Execute.scala 117:10]
  wire  _GEN_3855; // @[Execute.scala 117:10]
  wire  _GEN_3856; // @[Execute.scala 117:10]
  wire  _GEN_3857; // @[Execute.scala 117:10]
  wire  _GEN_3858; // @[Execute.scala 117:10]
  wire  _GEN_3859; // @[Execute.scala 117:10]
  wire  _GEN_3860; // @[Execute.scala 117:10]
  wire  _GEN_3861; // @[Execute.scala 117:10]
  wire  _GEN_3862; // @[Execute.scala 117:10]
  wire  _GEN_3863; // @[Execute.scala 117:10]
  wire  _GEN_3864; // @[Execute.scala 117:10]
  wire  _GEN_3865; // @[Execute.scala 117:10]
  wire  _GEN_3866; // @[Execute.scala 117:10]
  wire  _GEN_3867; // @[Execute.scala 117:10]
  wire  _GEN_3868; // @[Execute.scala 117:10]
  wire  _GEN_3869; // @[Execute.scala 117:10]
  wire  _GEN_3870; // @[Execute.scala 117:10]
  wire  _GEN_3871; // @[Execute.scala 117:10]
  wire  _GEN_3872; // @[Execute.scala 117:10]
  wire  _GEN_3873; // @[Execute.scala 117:10]
  wire  _GEN_3874; // @[Execute.scala 117:10]
  wire  _GEN_3875; // @[Execute.scala 117:10]
  wire  _GEN_3876; // @[Execute.scala 117:10]
  wire  _GEN_3877; // @[Execute.scala 117:10]
  wire  _GEN_3878; // @[Execute.scala 117:10]
  wire  _GEN_3879; // @[Execute.scala 117:10]
  wire  _GEN_3880; // @[Execute.scala 117:10]
  wire  _GEN_3881; // @[Execute.scala 117:10]
  wire  _GEN_3882; // @[Execute.scala 117:10]
  wire  _GEN_3883; // @[Execute.scala 117:10]
  wire  _GEN_3884; // @[Execute.scala 117:10]
  wire  _GEN_3885; // @[Execute.scala 117:10]
  wire  _GEN_3886; // @[Execute.scala 117:10]
  wire  _GEN_3887; // @[Execute.scala 117:10]
  wire  _GEN_3888; // @[Execute.scala 117:10]
  wire  _GEN_3889; // @[Execute.scala 117:10]
  wire  _GEN_3890; // @[Execute.scala 117:10]
  wire  _GEN_3891; // @[Execute.scala 117:10]
  wire  _GEN_3892; // @[Execute.scala 117:10]
  wire  _GEN_3893; // @[Execute.scala 117:10]
  wire  _GEN_3894; // @[Execute.scala 117:10]
  wire  _GEN_3895; // @[Execute.scala 117:10]
  wire  _GEN_3896; // @[Execute.scala 117:10]
  wire  _GEN_3897; // @[Execute.scala 117:10]
  wire  _GEN_3898; // @[Execute.scala 117:10]
  wire  _GEN_3899; // @[Execute.scala 117:10]
  wire  _GEN_3900; // @[Execute.scala 117:10]
  wire  _GEN_3901; // @[Execute.scala 117:10]
  wire  _GEN_3902; // @[Execute.scala 117:10]
  wire  _GEN_3903; // @[Execute.scala 117:10]
  wire  _GEN_3904; // @[Execute.scala 117:10]
  wire  _GEN_3905; // @[Execute.scala 117:10]
  wire  _GEN_3907; // @[Execute.scala 117:10]
  wire  _GEN_3908; // @[Execute.scala 117:10]
  wire  _GEN_3909; // @[Execute.scala 117:10]
  wire  _GEN_3910; // @[Execute.scala 117:10]
  wire  _GEN_3911; // @[Execute.scala 117:10]
  wire  _GEN_3912; // @[Execute.scala 117:10]
  wire  _GEN_3913; // @[Execute.scala 117:10]
  wire  _GEN_3914; // @[Execute.scala 117:10]
  wire  _GEN_3915; // @[Execute.scala 117:10]
  wire  _GEN_3916; // @[Execute.scala 117:10]
  wire  _GEN_3917; // @[Execute.scala 117:10]
  wire  _GEN_3918; // @[Execute.scala 117:10]
  wire  _GEN_3919; // @[Execute.scala 117:10]
  wire  _GEN_3920; // @[Execute.scala 117:10]
  wire  _GEN_3921; // @[Execute.scala 117:10]
  wire  _GEN_3922; // @[Execute.scala 117:10]
  wire  _GEN_3923; // @[Execute.scala 117:10]
  wire  _GEN_3924; // @[Execute.scala 117:10]
  wire  _GEN_3925; // @[Execute.scala 117:10]
  wire  _GEN_3926; // @[Execute.scala 117:10]
  wire  _GEN_3927; // @[Execute.scala 117:10]
  wire  _GEN_3928; // @[Execute.scala 117:10]
  wire  _GEN_3929; // @[Execute.scala 117:10]
  wire  _GEN_3930; // @[Execute.scala 117:10]
  wire  _GEN_3931; // @[Execute.scala 117:10]
  wire  _GEN_3932; // @[Execute.scala 117:10]
  wire  _GEN_3933; // @[Execute.scala 117:10]
  wire  _GEN_3934; // @[Execute.scala 117:10]
  wire  _GEN_3935; // @[Execute.scala 117:10]
  wire  _GEN_3936; // @[Execute.scala 117:10]
  wire  _GEN_3937; // @[Execute.scala 117:10]
  wire  _GEN_3938; // @[Execute.scala 117:10]
  wire  _GEN_3939; // @[Execute.scala 117:10]
  wire  _GEN_3940; // @[Execute.scala 117:10]
  wire  _GEN_3941; // @[Execute.scala 117:10]
  wire  _GEN_3942; // @[Execute.scala 117:10]
  wire  _GEN_3943; // @[Execute.scala 117:10]
  wire  _GEN_3944; // @[Execute.scala 117:10]
  wire  _GEN_3945; // @[Execute.scala 117:10]
  wire  _GEN_3946; // @[Execute.scala 117:10]
  wire  _GEN_3947; // @[Execute.scala 117:10]
  wire  _GEN_3948; // @[Execute.scala 117:10]
  wire  _GEN_3949; // @[Execute.scala 117:10]
  wire  _GEN_3950; // @[Execute.scala 117:10]
  wire  _GEN_3951; // @[Execute.scala 117:10]
  wire  _GEN_3952; // @[Execute.scala 117:10]
  wire  _GEN_3953; // @[Execute.scala 117:10]
  wire  _GEN_3954; // @[Execute.scala 117:10]
  wire  _GEN_3955; // @[Execute.scala 117:10]
  wire  _GEN_3956; // @[Execute.scala 117:10]
  wire  _GEN_3957; // @[Execute.scala 117:10]
  wire  _GEN_3958; // @[Execute.scala 117:10]
  wire  _GEN_3959; // @[Execute.scala 117:10]
  wire  _GEN_3960; // @[Execute.scala 117:10]
  wire  _GEN_3961; // @[Execute.scala 117:10]
  wire  _GEN_3962; // @[Execute.scala 117:10]
  wire  _GEN_3963; // @[Execute.scala 117:10]
  wire  _GEN_3964; // @[Execute.scala 117:10]
  wire  _GEN_3965; // @[Execute.scala 117:10]
  wire  _GEN_3966; // @[Execute.scala 117:10]
  wire  _GEN_3967; // @[Execute.scala 117:10]
  wire  _GEN_3968; // @[Execute.scala 117:10]
  wire  _GEN_3969; // @[Execute.scala 117:10]
  wire  _T_391; // @[Execute.scala 117:10]
  wire  _T_392; // @[Execute.scala 117:15]
  wire [5:0] _T_394; // @[Execute.scala 117:37]
  wire [5:0] _T_398; // @[Execute.scala 117:60]
  wire  _GEN_3971; // @[Execute.scala 117:10]
  wire  _GEN_3972; // @[Execute.scala 117:10]
  wire  _GEN_3973; // @[Execute.scala 117:10]
  wire  _GEN_3974; // @[Execute.scala 117:10]
  wire  _GEN_3975; // @[Execute.scala 117:10]
  wire  _GEN_3976; // @[Execute.scala 117:10]
  wire  _GEN_3977; // @[Execute.scala 117:10]
  wire  _GEN_3978; // @[Execute.scala 117:10]
  wire  _GEN_3979; // @[Execute.scala 117:10]
  wire  _GEN_3980; // @[Execute.scala 117:10]
  wire  _GEN_3981; // @[Execute.scala 117:10]
  wire  _GEN_3982; // @[Execute.scala 117:10]
  wire  _GEN_3983; // @[Execute.scala 117:10]
  wire  _GEN_3984; // @[Execute.scala 117:10]
  wire  _GEN_3985; // @[Execute.scala 117:10]
  wire  _GEN_3986; // @[Execute.scala 117:10]
  wire  _GEN_3987; // @[Execute.scala 117:10]
  wire  _GEN_3988; // @[Execute.scala 117:10]
  wire  _GEN_3989; // @[Execute.scala 117:10]
  wire  _GEN_3990; // @[Execute.scala 117:10]
  wire  _GEN_3991; // @[Execute.scala 117:10]
  wire  _GEN_3992; // @[Execute.scala 117:10]
  wire  _GEN_3993; // @[Execute.scala 117:10]
  wire  _GEN_3994; // @[Execute.scala 117:10]
  wire  _GEN_3995; // @[Execute.scala 117:10]
  wire  _GEN_3996; // @[Execute.scala 117:10]
  wire  _GEN_3997; // @[Execute.scala 117:10]
  wire  _GEN_3998; // @[Execute.scala 117:10]
  wire  _GEN_3999; // @[Execute.scala 117:10]
  wire  _GEN_4000; // @[Execute.scala 117:10]
  wire  _GEN_4001; // @[Execute.scala 117:10]
  wire  _GEN_4002; // @[Execute.scala 117:10]
  wire  _GEN_4003; // @[Execute.scala 117:10]
  wire  _GEN_4004; // @[Execute.scala 117:10]
  wire  _GEN_4005; // @[Execute.scala 117:10]
  wire  _GEN_4006; // @[Execute.scala 117:10]
  wire  _GEN_4007; // @[Execute.scala 117:10]
  wire  _GEN_4008; // @[Execute.scala 117:10]
  wire  _GEN_4009; // @[Execute.scala 117:10]
  wire  _GEN_4010; // @[Execute.scala 117:10]
  wire  _GEN_4011; // @[Execute.scala 117:10]
  wire  _GEN_4012; // @[Execute.scala 117:10]
  wire  _GEN_4013; // @[Execute.scala 117:10]
  wire  _GEN_4014; // @[Execute.scala 117:10]
  wire  _GEN_4015; // @[Execute.scala 117:10]
  wire  _GEN_4016; // @[Execute.scala 117:10]
  wire  _GEN_4017; // @[Execute.scala 117:10]
  wire  _GEN_4018; // @[Execute.scala 117:10]
  wire  _GEN_4019; // @[Execute.scala 117:10]
  wire  _GEN_4020; // @[Execute.scala 117:10]
  wire  _GEN_4021; // @[Execute.scala 117:10]
  wire  _GEN_4022; // @[Execute.scala 117:10]
  wire  _GEN_4023; // @[Execute.scala 117:10]
  wire  _GEN_4024; // @[Execute.scala 117:10]
  wire  _GEN_4025; // @[Execute.scala 117:10]
  wire  _GEN_4026; // @[Execute.scala 117:10]
  wire  _GEN_4027; // @[Execute.scala 117:10]
  wire  _GEN_4028; // @[Execute.scala 117:10]
  wire  _GEN_4029; // @[Execute.scala 117:10]
  wire  _GEN_4030; // @[Execute.scala 117:10]
  wire  _GEN_4031; // @[Execute.scala 117:10]
  wire  _GEN_4032; // @[Execute.scala 117:10]
  wire  _GEN_4033; // @[Execute.scala 117:10]
  wire  _GEN_4035; // @[Execute.scala 117:10]
  wire  _GEN_4036; // @[Execute.scala 117:10]
  wire  _GEN_4037; // @[Execute.scala 117:10]
  wire  _GEN_4038; // @[Execute.scala 117:10]
  wire  _GEN_4039; // @[Execute.scala 117:10]
  wire  _GEN_4040; // @[Execute.scala 117:10]
  wire  _GEN_4041; // @[Execute.scala 117:10]
  wire  _GEN_4042; // @[Execute.scala 117:10]
  wire  _GEN_4043; // @[Execute.scala 117:10]
  wire  _GEN_4044; // @[Execute.scala 117:10]
  wire  _GEN_4045; // @[Execute.scala 117:10]
  wire  _GEN_4046; // @[Execute.scala 117:10]
  wire  _GEN_4047; // @[Execute.scala 117:10]
  wire  _GEN_4048; // @[Execute.scala 117:10]
  wire  _GEN_4049; // @[Execute.scala 117:10]
  wire  _GEN_4050; // @[Execute.scala 117:10]
  wire  _GEN_4051; // @[Execute.scala 117:10]
  wire  _GEN_4052; // @[Execute.scala 117:10]
  wire  _GEN_4053; // @[Execute.scala 117:10]
  wire  _GEN_4054; // @[Execute.scala 117:10]
  wire  _GEN_4055; // @[Execute.scala 117:10]
  wire  _GEN_4056; // @[Execute.scala 117:10]
  wire  _GEN_4057; // @[Execute.scala 117:10]
  wire  _GEN_4058; // @[Execute.scala 117:10]
  wire  _GEN_4059; // @[Execute.scala 117:10]
  wire  _GEN_4060; // @[Execute.scala 117:10]
  wire  _GEN_4061; // @[Execute.scala 117:10]
  wire  _GEN_4062; // @[Execute.scala 117:10]
  wire  _GEN_4063; // @[Execute.scala 117:10]
  wire  _GEN_4064; // @[Execute.scala 117:10]
  wire  _GEN_4065; // @[Execute.scala 117:10]
  wire  _GEN_4066; // @[Execute.scala 117:10]
  wire  _GEN_4067; // @[Execute.scala 117:10]
  wire  _GEN_4068; // @[Execute.scala 117:10]
  wire  _GEN_4069; // @[Execute.scala 117:10]
  wire  _GEN_4070; // @[Execute.scala 117:10]
  wire  _GEN_4071; // @[Execute.scala 117:10]
  wire  _GEN_4072; // @[Execute.scala 117:10]
  wire  _GEN_4073; // @[Execute.scala 117:10]
  wire  _GEN_4074; // @[Execute.scala 117:10]
  wire  _GEN_4075; // @[Execute.scala 117:10]
  wire  _GEN_4076; // @[Execute.scala 117:10]
  wire  _GEN_4077; // @[Execute.scala 117:10]
  wire  _GEN_4078; // @[Execute.scala 117:10]
  wire  _GEN_4079; // @[Execute.scala 117:10]
  wire  _GEN_4080; // @[Execute.scala 117:10]
  wire  _GEN_4081; // @[Execute.scala 117:10]
  wire  _GEN_4082; // @[Execute.scala 117:10]
  wire  _GEN_4083; // @[Execute.scala 117:10]
  wire  _GEN_4084; // @[Execute.scala 117:10]
  wire  _GEN_4085; // @[Execute.scala 117:10]
  wire  _GEN_4086; // @[Execute.scala 117:10]
  wire  _GEN_4087; // @[Execute.scala 117:10]
  wire  _GEN_4088; // @[Execute.scala 117:10]
  wire  _GEN_4089; // @[Execute.scala 117:10]
  wire  _GEN_4090; // @[Execute.scala 117:10]
  wire  _GEN_4091; // @[Execute.scala 117:10]
  wire  _GEN_4092; // @[Execute.scala 117:10]
  wire  _GEN_4093; // @[Execute.scala 117:10]
  wire  _GEN_4094; // @[Execute.scala 117:10]
  wire  _GEN_4095; // @[Execute.scala 117:10]
  wire  _GEN_4096; // @[Execute.scala 117:10]
  wire  _GEN_4097; // @[Execute.scala 117:10]
  wire  _T_401; // @[Execute.scala 117:10]
  wire  _T_402; // @[Execute.scala 117:15]
  wire [5:0] _T_404; // @[Execute.scala 117:37]
  wire [5:0] _T_408; // @[Execute.scala 117:60]
  wire  _GEN_4099; // @[Execute.scala 117:10]
  wire  _GEN_4100; // @[Execute.scala 117:10]
  wire  _GEN_4101; // @[Execute.scala 117:10]
  wire  _GEN_4102; // @[Execute.scala 117:10]
  wire  _GEN_4103; // @[Execute.scala 117:10]
  wire  _GEN_4104; // @[Execute.scala 117:10]
  wire  _GEN_4105; // @[Execute.scala 117:10]
  wire  _GEN_4106; // @[Execute.scala 117:10]
  wire  _GEN_4107; // @[Execute.scala 117:10]
  wire  _GEN_4108; // @[Execute.scala 117:10]
  wire  _GEN_4109; // @[Execute.scala 117:10]
  wire  _GEN_4110; // @[Execute.scala 117:10]
  wire  _GEN_4111; // @[Execute.scala 117:10]
  wire  _GEN_4112; // @[Execute.scala 117:10]
  wire  _GEN_4113; // @[Execute.scala 117:10]
  wire  _GEN_4114; // @[Execute.scala 117:10]
  wire  _GEN_4115; // @[Execute.scala 117:10]
  wire  _GEN_4116; // @[Execute.scala 117:10]
  wire  _GEN_4117; // @[Execute.scala 117:10]
  wire  _GEN_4118; // @[Execute.scala 117:10]
  wire  _GEN_4119; // @[Execute.scala 117:10]
  wire  _GEN_4120; // @[Execute.scala 117:10]
  wire  _GEN_4121; // @[Execute.scala 117:10]
  wire  _GEN_4122; // @[Execute.scala 117:10]
  wire  _GEN_4123; // @[Execute.scala 117:10]
  wire  _GEN_4124; // @[Execute.scala 117:10]
  wire  _GEN_4125; // @[Execute.scala 117:10]
  wire  _GEN_4126; // @[Execute.scala 117:10]
  wire  _GEN_4127; // @[Execute.scala 117:10]
  wire  _GEN_4128; // @[Execute.scala 117:10]
  wire  _GEN_4129; // @[Execute.scala 117:10]
  wire  _GEN_4130; // @[Execute.scala 117:10]
  wire  _GEN_4131; // @[Execute.scala 117:10]
  wire  _GEN_4132; // @[Execute.scala 117:10]
  wire  _GEN_4133; // @[Execute.scala 117:10]
  wire  _GEN_4134; // @[Execute.scala 117:10]
  wire  _GEN_4135; // @[Execute.scala 117:10]
  wire  _GEN_4136; // @[Execute.scala 117:10]
  wire  _GEN_4137; // @[Execute.scala 117:10]
  wire  _GEN_4138; // @[Execute.scala 117:10]
  wire  _GEN_4139; // @[Execute.scala 117:10]
  wire  _GEN_4140; // @[Execute.scala 117:10]
  wire  _GEN_4141; // @[Execute.scala 117:10]
  wire  _GEN_4142; // @[Execute.scala 117:10]
  wire  _GEN_4143; // @[Execute.scala 117:10]
  wire  _GEN_4144; // @[Execute.scala 117:10]
  wire  _GEN_4145; // @[Execute.scala 117:10]
  wire  _GEN_4146; // @[Execute.scala 117:10]
  wire  _GEN_4147; // @[Execute.scala 117:10]
  wire  _GEN_4148; // @[Execute.scala 117:10]
  wire  _GEN_4149; // @[Execute.scala 117:10]
  wire  _GEN_4150; // @[Execute.scala 117:10]
  wire  _GEN_4151; // @[Execute.scala 117:10]
  wire  _GEN_4152; // @[Execute.scala 117:10]
  wire  _GEN_4153; // @[Execute.scala 117:10]
  wire  _GEN_4154; // @[Execute.scala 117:10]
  wire  _GEN_4155; // @[Execute.scala 117:10]
  wire  _GEN_4156; // @[Execute.scala 117:10]
  wire  _GEN_4157; // @[Execute.scala 117:10]
  wire  _GEN_4158; // @[Execute.scala 117:10]
  wire  _GEN_4159; // @[Execute.scala 117:10]
  wire  _GEN_4160; // @[Execute.scala 117:10]
  wire  _GEN_4161; // @[Execute.scala 117:10]
  wire  _GEN_4163; // @[Execute.scala 117:10]
  wire  _GEN_4164; // @[Execute.scala 117:10]
  wire  _GEN_4165; // @[Execute.scala 117:10]
  wire  _GEN_4166; // @[Execute.scala 117:10]
  wire  _GEN_4167; // @[Execute.scala 117:10]
  wire  _GEN_4168; // @[Execute.scala 117:10]
  wire  _GEN_4169; // @[Execute.scala 117:10]
  wire  _GEN_4170; // @[Execute.scala 117:10]
  wire  _GEN_4171; // @[Execute.scala 117:10]
  wire  _GEN_4172; // @[Execute.scala 117:10]
  wire  _GEN_4173; // @[Execute.scala 117:10]
  wire  _GEN_4174; // @[Execute.scala 117:10]
  wire  _GEN_4175; // @[Execute.scala 117:10]
  wire  _GEN_4176; // @[Execute.scala 117:10]
  wire  _GEN_4177; // @[Execute.scala 117:10]
  wire  _GEN_4178; // @[Execute.scala 117:10]
  wire  _GEN_4179; // @[Execute.scala 117:10]
  wire  _GEN_4180; // @[Execute.scala 117:10]
  wire  _GEN_4181; // @[Execute.scala 117:10]
  wire  _GEN_4182; // @[Execute.scala 117:10]
  wire  _GEN_4183; // @[Execute.scala 117:10]
  wire  _GEN_4184; // @[Execute.scala 117:10]
  wire  _GEN_4185; // @[Execute.scala 117:10]
  wire  _GEN_4186; // @[Execute.scala 117:10]
  wire  _GEN_4187; // @[Execute.scala 117:10]
  wire  _GEN_4188; // @[Execute.scala 117:10]
  wire  _GEN_4189; // @[Execute.scala 117:10]
  wire  _GEN_4190; // @[Execute.scala 117:10]
  wire  _GEN_4191; // @[Execute.scala 117:10]
  wire  _GEN_4192; // @[Execute.scala 117:10]
  wire  _GEN_4193; // @[Execute.scala 117:10]
  wire  _GEN_4194; // @[Execute.scala 117:10]
  wire  _GEN_4195; // @[Execute.scala 117:10]
  wire  _GEN_4196; // @[Execute.scala 117:10]
  wire  _GEN_4197; // @[Execute.scala 117:10]
  wire  _GEN_4198; // @[Execute.scala 117:10]
  wire  _GEN_4199; // @[Execute.scala 117:10]
  wire  _GEN_4200; // @[Execute.scala 117:10]
  wire  _GEN_4201; // @[Execute.scala 117:10]
  wire  _GEN_4202; // @[Execute.scala 117:10]
  wire  _GEN_4203; // @[Execute.scala 117:10]
  wire  _GEN_4204; // @[Execute.scala 117:10]
  wire  _GEN_4205; // @[Execute.scala 117:10]
  wire  _GEN_4206; // @[Execute.scala 117:10]
  wire  _GEN_4207; // @[Execute.scala 117:10]
  wire  _GEN_4208; // @[Execute.scala 117:10]
  wire  _GEN_4209; // @[Execute.scala 117:10]
  wire  _GEN_4210; // @[Execute.scala 117:10]
  wire  _GEN_4211; // @[Execute.scala 117:10]
  wire  _GEN_4212; // @[Execute.scala 117:10]
  wire  _GEN_4213; // @[Execute.scala 117:10]
  wire  _GEN_4214; // @[Execute.scala 117:10]
  wire  _GEN_4215; // @[Execute.scala 117:10]
  wire  _GEN_4216; // @[Execute.scala 117:10]
  wire  _GEN_4217; // @[Execute.scala 117:10]
  wire  _GEN_4218; // @[Execute.scala 117:10]
  wire  _GEN_4219; // @[Execute.scala 117:10]
  wire  _GEN_4220; // @[Execute.scala 117:10]
  wire  _GEN_4221; // @[Execute.scala 117:10]
  wire  _GEN_4222; // @[Execute.scala 117:10]
  wire  _GEN_4223; // @[Execute.scala 117:10]
  wire  _GEN_4224; // @[Execute.scala 117:10]
  wire  _GEN_4225; // @[Execute.scala 117:10]
  wire  _T_411; // @[Execute.scala 117:10]
  wire  _T_412; // @[Execute.scala 117:15]
  wire [5:0] _T_414; // @[Execute.scala 117:37]
  wire [5:0] _T_418; // @[Execute.scala 117:60]
  wire  _GEN_4227; // @[Execute.scala 117:10]
  wire  _GEN_4228; // @[Execute.scala 117:10]
  wire  _GEN_4229; // @[Execute.scala 117:10]
  wire  _GEN_4230; // @[Execute.scala 117:10]
  wire  _GEN_4231; // @[Execute.scala 117:10]
  wire  _GEN_4232; // @[Execute.scala 117:10]
  wire  _GEN_4233; // @[Execute.scala 117:10]
  wire  _GEN_4234; // @[Execute.scala 117:10]
  wire  _GEN_4235; // @[Execute.scala 117:10]
  wire  _GEN_4236; // @[Execute.scala 117:10]
  wire  _GEN_4237; // @[Execute.scala 117:10]
  wire  _GEN_4238; // @[Execute.scala 117:10]
  wire  _GEN_4239; // @[Execute.scala 117:10]
  wire  _GEN_4240; // @[Execute.scala 117:10]
  wire  _GEN_4241; // @[Execute.scala 117:10]
  wire  _GEN_4242; // @[Execute.scala 117:10]
  wire  _GEN_4243; // @[Execute.scala 117:10]
  wire  _GEN_4244; // @[Execute.scala 117:10]
  wire  _GEN_4245; // @[Execute.scala 117:10]
  wire  _GEN_4246; // @[Execute.scala 117:10]
  wire  _GEN_4247; // @[Execute.scala 117:10]
  wire  _GEN_4248; // @[Execute.scala 117:10]
  wire  _GEN_4249; // @[Execute.scala 117:10]
  wire  _GEN_4250; // @[Execute.scala 117:10]
  wire  _GEN_4251; // @[Execute.scala 117:10]
  wire  _GEN_4252; // @[Execute.scala 117:10]
  wire  _GEN_4253; // @[Execute.scala 117:10]
  wire  _GEN_4254; // @[Execute.scala 117:10]
  wire  _GEN_4255; // @[Execute.scala 117:10]
  wire  _GEN_4256; // @[Execute.scala 117:10]
  wire  _GEN_4257; // @[Execute.scala 117:10]
  wire  _GEN_4258; // @[Execute.scala 117:10]
  wire  _GEN_4259; // @[Execute.scala 117:10]
  wire  _GEN_4260; // @[Execute.scala 117:10]
  wire  _GEN_4261; // @[Execute.scala 117:10]
  wire  _GEN_4262; // @[Execute.scala 117:10]
  wire  _GEN_4263; // @[Execute.scala 117:10]
  wire  _GEN_4264; // @[Execute.scala 117:10]
  wire  _GEN_4265; // @[Execute.scala 117:10]
  wire  _GEN_4266; // @[Execute.scala 117:10]
  wire  _GEN_4267; // @[Execute.scala 117:10]
  wire  _GEN_4268; // @[Execute.scala 117:10]
  wire  _GEN_4269; // @[Execute.scala 117:10]
  wire  _GEN_4270; // @[Execute.scala 117:10]
  wire  _GEN_4271; // @[Execute.scala 117:10]
  wire  _GEN_4272; // @[Execute.scala 117:10]
  wire  _GEN_4273; // @[Execute.scala 117:10]
  wire  _GEN_4274; // @[Execute.scala 117:10]
  wire  _GEN_4275; // @[Execute.scala 117:10]
  wire  _GEN_4276; // @[Execute.scala 117:10]
  wire  _GEN_4277; // @[Execute.scala 117:10]
  wire  _GEN_4278; // @[Execute.scala 117:10]
  wire  _GEN_4279; // @[Execute.scala 117:10]
  wire  _GEN_4280; // @[Execute.scala 117:10]
  wire  _GEN_4281; // @[Execute.scala 117:10]
  wire  _GEN_4282; // @[Execute.scala 117:10]
  wire  _GEN_4283; // @[Execute.scala 117:10]
  wire  _GEN_4284; // @[Execute.scala 117:10]
  wire  _GEN_4285; // @[Execute.scala 117:10]
  wire  _GEN_4286; // @[Execute.scala 117:10]
  wire  _GEN_4287; // @[Execute.scala 117:10]
  wire  _GEN_4288; // @[Execute.scala 117:10]
  wire  _GEN_4289; // @[Execute.scala 117:10]
  wire  _GEN_4291; // @[Execute.scala 117:10]
  wire  _GEN_4292; // @[Execute.scala 117:10]
  wire  _GEN_4293; // @[Execute.scala 117:10]
  wire  _GEN_4294; // @[Execute.scala 117:10]
  wire  _GEN_4295; // @[Execute.scala 117:10]
  wire  _GEN_4296; // @[Execute.scala 117:10]
  wire  _GEN_4297; // @[Execute.scala 117:10]
  wire  _GEN_4298; // @[Execute.scala 117:10]
  wire  _GEN_4299; // @[Execute.scala 117:10]
  wire  _GEN_4300; // @[Execute.scala 117:10]
  wire  _GEN_4301; // @[Execute.scala 117:10]
  wire  _GEN_4302; // @[Execute.scala 117:10]
  wire  _GEN_4303; // @[Execute.scala 117:10]
  wire  _GEN_4304; // @[Execute.scala 117:10]
  wire  _GEN_4305; // @[Execute.scala 117:10]
  wire  _GEN_4306; // @[Execute.scala 117:10]
  wire  _GEN_4307; // @[Execute.scala 117:10]
  wire  _GEN_4308; // @[Execute.scala 117:10]
  wire  _GEN_4309; // @[Execute.scala 117:10]
  wire  _GEN_4310; // @[Execute.scala 117:10]
  wire  _GEN_4311; // @[Execute.scala 117:10]
  wire  _GEN_4312; // @[Execute.scala 117:10]
  wire  _GEN_4313; // @[Execute.scala 117:10]
  wire  _GEN_4314; // @[Execute.scala 117:10]
  wire  _GEN_4315; // @[Execute.scala 117:10]
  wire  _GEN_4316; // @[Execute.scala 117:10]
  wire  _GEN_4317; // @[Execute.scala 117:10]
  wire  _GEN_4318; // @[Execute.scala 117:10]
  wire  _GEN_4319; // @[Execute.scala 117:10]
  wire  _GEN_4320; // @[Execute.scala 117:10]
  wire  _GEN_4321; // @[Execute.scala 117:10]
  wire  _GEN_4322; // @[Execute.scala 117:10]
  wire  _GEN_4323; // @[Execute.scala 117:10]
  wire  _GEN_4324; // @[Execute.scala 117:10]
  wire  _GEN_4325; // @[Execute.scala 117:10]
  wire  _GEN_4326; // @[Execute.scala 117:10]
  wire  _GEN_4327; // @[Execute.scala 117:10]
  wire  _GEN_4328; // @[Execute.scala 117:10]
  wire  _GEN_4329; // @[Execute.scala 117:10]
  wire  _GEN_4330; // @[Execute.scala 117:10]
  wire  _GEN_4331; // @[Execute.scala 117:10]
  wire  _GEN_4332; // @[Execute.scala 117:10]
  wire  _GEN_4333; // @[Execute.scala 117:10]
  wire  _GEN_4334; // @[Execute.scala 117:10]
  wire  _GEN_4335; // @[Execute.scala 117:10]
  wire  _GEN_4336; // @[Execute.scala 117:10]
  wire  _GEN_4337; // @[Execute.scala 117:10]
  wire  _GEN_4338; // @[Execute.scala 117:10]
  wire  _GEN_4339; // @[Execute.scala 117:10]
  wire  _GEN_4340; // @[Execute.scala 117:10]
  wire  _GEN_4341; // @[Execute.scala 117:10]
  wire  _GEN_4342; // @[Execute.scala 117:10]
  wire  _GEN_4343; // @[Execute.scala 117:10]
  wire  _GEN_4344; // @[Execute.scala 117:10]
  wire  _GEN_4345; // @[Execute.scala 117:10]
  wire  _GEN_4346; // @[Execute.scala 117:10]
  wire  _GEN_4347; // @[Execute.scala 117:10]
  wire  _GEN_4348; // @[Execute.scala 117:10]
  wire  _GEN_4349; // @[Execute.scala 117:10]
  wire  _GEN_4350; // @[Execute.scala 117:10]
  wire  _GEN_4351; // @[Execute.scala 117:10]
  wire  _GEN_4352; // @[Execute.scala 117:10]
  wire  _GEN_4353; // @[Execute.scala 117:10]
  wire  _T_421; // @[Execute.scala 117:10]
  wire  _T_422; // @[Execute.scala 117:15]
  wire [5:0] _T_424; // @[Execute.scala 117:37]
  wire [5:0] _T_428; // @[Execute.scala 117:60]
  wire  _GEN_4355; // @[Execute.scala 117:10]
  wire  _GEN_4356; // @[Execute.scala 117:10]
  wire  _GEN_4357; // @[Execute.scala 117:10]
  wire  _GEN_4358; // @[Execute.scala 117:10]
  wire  _GEN_4359; // @[Execute.scala 117:10]
  wire  _GEN_4360; // @[Execute.scala 117:10]
  wire  _GEN_4361; // @[Execute.scala 117:10]
  wire  _GEN_4362; // @[Execute.scala 117:10]
  wire  _GEN_4363; // @[Execute.scala 117:10]
  wire  _GEN_4364; // @[Execute.scala 117:10]
  wire  _GEN_4365; // @[Execute.scala 117:10]
  wire  _GEN_4366; // @[Execute.scala 117:10]
  wire  _GEN_4367; // @[Execute.scala 117:10]
  wire  _GEN_4368; // @[Execute.scala 117:10]
  wire  _GEN_4369; // @[Execute.scala 117:10]
  wire  _GEN_4370; // @[Execute.scala 117:10]
  wire  _GEN_4371; // @[Execute.scala 117:10]
  wire  _GEN_4372; // @[Execute.scala 117:10]
  wire  _GEN_4373; // @[Execute.scala 117:10]
  wire  _GEN_4374; // @[Execute.scala 117:10]
  wire  _GEN_4375; // @[Execute.scala 117:10]
  wire  _GEN_4376; // @[Execute.scala 117:10]
  wire  _GEN_4377; // @[Execute.scala 117:10]
  wire  _GEN_4378; // @[Execute.scala 117:10]
  wire  _GEN_4379; // @[Execute.scala 117:10]
  wire  _GEN_4380; // @[Execute.scala 117:10]
  wire  _GEN_4381; // @[Execute.scala 117:10]
  wire  _GEN_4382; // @[Execute.scala 117:10]
  wire  _GEN_4383; // @[Execute.scala 117:10]
  wire  _GEN_4384; // @[Execute.scala 117:10]
  wire  _GEN_4385; // @[Execute.scala 117:10]
  wire  _GEN_4386; // @[Execute.scala 117:10]
  wire  _GEN_4387; // @[Execute.scala 117:10]
  wire  _GEN_4388; // @[Execute.scala 117:10]
  wire  _GEN_4389; // @[Execute.scala 117:10]
  wire  _GEN_4390; // @[Execute.scala 117:10]
  wire  _GEN_4391; // @[Execute.scala 117:10]
  wire  _GEN_4392; // @[Execute.scala 117:10]
  wire  _GEN_4393; // @[Execute.scala 117:10]
  wire  _GEN_4394; // @[Execute.scala 117:10]
  wire  _GEN_4395; // @[Execute.scala 117:10]
  wire  _GEN_4396; // @[Execute.scala 117:10]
  wire  _GEN_4397; // @[Execute.scala 117:10]
  wire  _GEN_4398; // @[Execute.scala 117:10]
  wire  _GEN_4399; // @[Execute.scala 117:10]
  wire  _GEN_4400; // @[Execute.scala 117:10]
  wire  _GEN_4401; // @[Execute.scala 117:10]
  wire  _GEN_4402; // @[Execute.scala 117:10]
  wire  _GEN_4403; // @[Execute.scala 117:10]
  wire  _GEN_4404; // @[Execute.scala 117:10]
  wire  _GEN_4405; // @[Execute.scala 117:10]
  wire  _GEN_4406; // @[Execute.scala 117:10]
  wire  _GEN_4407; // @[Execute.scala 117:10]
  wire  _GEN_4408; // @[Execute.scala 117:10]
  wire  _GEN_4409; // @[Execute.scala 117:10]
  wire  _GEN_4410; // @[Execute.scala 117:10]
  wire  _GEN_4411; // @[Execute.scala 117:10]
  wire  _GEN_4412; // @[Execute.scala 117:10]
  wire  _GEN_4413; // @[Execute.scala 117:10]
  wire  _GEN_4414; // @[Execute.scala 117:10]
  wire  _GEN_4415; // @[Execute.scala 117:10]
  wire  _GEN_4416; // @[Execute.scala 117:10]
  wire  _GEN_4417; // @[Execute.scala 117:10]
  wire  _GEN_4419; // @[Execute.scala 117:10]
  wire  _GEN_4420; // @[Execute.scala 117:10]
  wire  _GEN_4421; // @[Execute.scala 117:10]
  wire  _GEN_4422; // @[Execute.scala 117:10]
  wire  _GEN_4423; // @[Execute.scala 117:10]
  wire  _GEN_4424; // @[Execute.scala 117:10]
  wire  _GEN_4425; // @[Execute.scala 117:10]
  wire  _GEN_4426; // @[Execute.scala 117:10]
  wire  _GEN_4427; // @[Execute.scala 117:10]
  wire  _GEN_4428; // @[Execute.scala 117:10]
  wire  _GEN_4429; // @[Execute.scala 117:10]
  wire  _GEN_4430; // @[Execute.scala 117:10]
  wire  _GEN_4431; // @[Execute.scala 117:10]
  wire  _GEN_4432; // @[Execute.scala 117:10]
  wire  _GEN_4433; // @[Execute.scala 117:10]
  wire  _GEN_4434; // @[Execute.scala 117:10]
  wire  _GEN_4435; // @[Execute.scala 117:10]
  wire  _GEN_4436; // @[Execute.scala 117:10]
  wire  _GEN_4437; // @[Execute.scala 117:10]
  wire  _GEN_4438; // @[Execute.scala 117:10]
  wire  _GEN_4439; // @[Execute.scala 117:10]
  wire  _GEN_4440; // @[Execute.scala 117:10]
  wire  _GEN_4441; // @[Execute.scala 117:10]
  wire  _GEN_4442; // @[Execute.scala 117:10]
  wire  _GEN_4443; // @[Execute.scala 117:10]
  wire  _GEN_4444; // @[Execute.scala 117:10]
  wire  _GEN_4445; // @[Execute.scala 117:10]
  wire  _GEN_4446; // @[Execute.scala 117:10]
  wire  _GEN_4447; // @[Execute.scala 117:10]
  wire  _GEN_4448; // @[Execute.scala 117:10]
  wire  _GEN_4449; // @[Execute.scala 117:10]
  wire  _GEN_4450; // @[Execute.scala 117:10]
  wire  _GEN_4451; // @[Execute.scala 117:10]
  wire  _GEN_4452; // @[Execute.scala 117:10]
  wire  _GEN_4453; // @[Execute.scala 117:10]
  wire  _GEN_4454; // @[Execute.scala 117:10]
  wire  _GEN_4455; // @[Execute.scala 117:10]
  wire  _GEN_4456; // @[Execute.scala 117:10]
  wire  _GEN_4457; // @[Execute.scala 117:10]
  wire  _GEN_4458; // @[Execute.scala 117:10]
  wire  _GEN_4459; // @[Execute.scala 117:10]
  wire  _GEN_4460; // @[Execute.scala 117:10]
  wire  _GEN_4461; // @[Execute.scala 117:10]
  wire  _GEN_4462; // @[Execute.scala 117:10]
  wire  _GEN_4463; // @[Execute.scala 117:10]
  wire  _GEN_4464; // @[Execute.scala 117:10]
  wire  _GEN_4465; // @[Execute.scala 117:10]
  wire  _GEN_4466; // @[Execute.scala 117:10]
  wire  _GEN_4467; // @[Execute.scala 117:10]
  wire  _GEN_4468; // @[Execute.scala 117:10]
  wire  _GEN_4469; // @[Execute.scala 117:10]
  wire  _GEN_4470; // @[Execute.scala 117:10]
  wire  _GEN_4471; // @[Execute.scala 117:10]
  wire  _GEN_4472; // @[Execute.scala 117:10]
  wire  _GEN_4473; // @[Execute.scala 117:10]
  wire  _GEN_4474; // @[Execute.scala 117:10]
  wire  _GEN_4475; // @[Execute.scala 117:10]
  wire  _GEN_4476; // @[Execute.scala 117:10]
  wire  _GEN_4477; // @[Execute.scala 117:10]
  wire  _GEN_4478; // @[Execute.scala 117:10]
  wire  _GEN_4479; // @[Execute.scala 117:10]
  wire  _GEN_4480; // @[Execute.scala 117:10]
  wire  _GEN_4481; // @[Execute.scala 117:10]
  wire  _T_431; // @[Execute.scala 117:10]
  wire  _T_432; // @[Execute.scala 117:15]
  wire [5:0] _T_434; // @[Execute.scala 117:37]
  wire [5:0] _T_438; // @[Execute.scala 117:60]
  wire  _GEN_4483; // @[Execute.scala 117:10]
  wire  _GEN_4484; // @[Execute.scala 117:10]
  wire  _GEN_4485; // @[Execute.scala 117:10]
  wire  _GEN_4486; // @[Execute.scala 117:10]
  wire  _GEN_4487; // @[Execute.scala 117:10]
  wire  _GEN_4488; // @[Execute.scala 117:10]
  wire  _GEN_4489; // @[Execute.scala 117:10]
  wire  _GEN_4490; // @[Execute.scala 117:10]
  wire  _GEN_4491; // @[Execute.scala 117:10]
  wire  _GEN_4492; // @[Execute.scala 117:10]
  wire  _GEN_4493; // @[Execute.scala 117:10]
  wire  _GEN_4494; // @[Execute.scala 117:10]
  wire  _GEN_4495; // @[Execute.scala 117:10]
  wire  _GEN_4496; // @[Execute.scala 117:10]
  wire  _GEN_4497; // @[Execute.scala 117:10]
  wire  _GEN_4498; // @[Execute.scala 117:10]
  wire  _GEN_4499; // @[Execute.scala 117:10]
  wire  _GEN_4500; // @[Execute.scala 117:10]
  wire  _GEN_4501; // @[Execute.scala 117:10]
  wire  _GEN_4502; // @[Execute.scala 117:10]
  wire  _GEN_4503; // @[Execute.scala 117:10]
  wire  _GEN_4504; // @[Execute.scala 117:10]
  wire  _GEN_4505; // @[Execute.scala 117:10]
  wire  _GEN_4506; // @[Execute.scala 117:10]
  wire  _GEN_4507; // @[Execute.scala 117:10]
  wire  _GEN_4508; // @[Execute.scala 117:10]
  wire  _GEN_4509; // @[Execute.scala 117:10]
  wire  _GEN_4510; // @[Execute.scala 117:10]
  wire  _GEN_4511; // @[Execute.scala 117:10]
  wire  _GEN_4512; // @[Execute.scala 117:10]
  wire  _GEN_4513; // @[Execute.scala 117:10]
  wire  _GEN_4514; // @[Execute.scala 117:10]
  wire  _GEN_4515; // @[Execute.scala 117:10]
  wire  _GEN_4516; // @[Execute.scala 117:10]
  wire  _GEN_4517; // @[Execute.scala 117:10]
  wire  _GEN_4518; // @[Execute.scala 117:10]
  wire  _GEN_4519; // @[Execute.scala 117:10]
  wire  _GEN_4520; // @[Execute.scala 117:10]
  wire  _GEN_4521; // @[Execute.scala 117:10]
  wire  _GEN_4522; // @[Execute.scala 117:10]
  wire  _GEN_4523; // @[Execute.scala 117:10]
  wire  _GEN_4524; // @[Execute.scala 117:10]
  wire  _GEN_4525; // @[Execute.scala 117:10]
  wire  _GEN_4526; // @[Execute.scala 117:10]
  wire  _GEN_4527; // @[Execute.scala 117:10]
  wire  _GEN_4528; // @[Execute.scala 117:10]
  wire  _GEN_4529; // @[Execute.scala 117:10]
  wire  _GEN_4530; // @[Execute.scala 117:10]
  wire  _GEN_4531; // @[Execute.scala 117:10]
  wire  _GEN_4532; // @[Execute.scala 117:10]
  wire  _GEN_4533; // @[Execute.scala 117:10]
  wire  _GEN_4534; // @[Execute.scala 117:10]
  wire  _GEN_4535; // @[Execute.scala 117:10]
  wire  _GEN_4536; // @[Execute.scala 117:10]
  wire  _GEN_4537; // @[Execute.scala 117:10]
  wire  _GEN_4538; // @[Execute.scala 117:10]
  wire  _GEN_4539; // @[Execute.scala 117:10]
  wire  _GEN_4540; // @[Execute.scala 117:10]
  wire  _GEN_4541; // @[Execute.scala 117:10]
  wire  _GEN_4542; // @[Execute.scala 117:10]
  wire  _GEN_4543; // @[Execute.scala 117:10]
  wire  _GEN_4544; // @[Execute.scala 117:10]
  wire  _GEN_4545; // @[Execute.scala 117:10]
  wire  _GEN_4547; // @[Execute.scala 117:10]
  wire  _GEN_4548; // @[Execute.scala 117:10]
  wire  _GEN_4549; // @[Execute.scala 117:10]
  wire  _GEN_4550; // @[Execute.scala 117:10]
  wire  _GEN_4551; // @[Execute.scala 117:10]
  wire  _GEN_4552; // @[Execute.scala 117:10]
  wire  _GEN_4553; // @[Execute.scala 117:10]
  wire  _GEN_4554; // @[Execute.scala 117:10]
  wire  _GEN_4555; // @[Execute.scala 117:10]
  wire  _GEN_4556; // @[Execute.scala 117:10]
  wire  _GEN_4557; // @[Execute.scala 117:10]
  wire  _GEN_4558; // @[Execute.scala 117:10]
  wire  _GEN_4559; // @[Execute.scala 117:10]
  wire  _GEN_4560; // @[Execute.scala 117:10]
  wire  _GEN_4561; // @[Execute.scala 117:10]
  wire  _GEN_4562; // @[Execute.scala 117:10]
  wire  _GEN_4563; // @[Execute.scala 117:10]
  wire  _GEN_4564; // @[Execute.scala 117:10]
  wire  _GEN_4565; // @[Execute.scala 117:10]
  wire  _GEN_4566; // @[Execute.scala 117:10]
  wire  _GEN_4567; // @[Execute.scala 117:10]
  wire  _GEN_4568; // @[Execute.scala 117:10]
  wire  _GEN_4569; // @[Execute.scala 117:10]
  wire  _GEN_4570; // @[Execute.scala 117:10]
  wire  _GEN_4571; // @[Execute.scala 117:10]
  wire  _GEN_4572; // @[Execute.scala 117:10]
  wire  _GEN_4573; // @[Execute.scala 117:10]
  wire  _GEN_4574; // @[Execute.scala 117:10]
  wire  _GEN_4575; // @[Execute.scala 117:10]
  wire  _GEN_4576; // @[Execute.scala 117:10]
  wire  _GEN_4577; // @[Execute.scala 117:10]
  wire  _GEN_4578; // @[Execute.scala 117:10]
  wire  _GEN_4579; // @[Execute.scala 117:10]
  wire  _GEN_4580; // @[Execute.scala 117:10]
  wire  _GEN_4581; // @[Execute.scala 117:10]
  wire  _GEN_4582; // @[Execute.scala 117:10]
  wire  _GEN_4583; // @[Execute.scala 117:10]
  wire  _GEN_4584; // @[Execute.scala 117:10]
  wire  _GEN_4585; // @[Execute.scala 117:10]
  wire  _GEN_4586; // @[Execute.scala 117:10]
  wire  _GEN_4587; // @[Execute.scala 117:10]
  wire  _GEN_4588; // @[Execute.scala 117:10]
  wire  _GEN_4589; // @[Execute.scala 117:10]
  wire  _GEN_4590; // @[Execute.scala 117:10]
  wire  _GEN_4591; // @[Execute.scala 117:10]
  wire  _GEN_4592; // @[Execute.scala 117:10]
  wire  _GEN_4593; // @[Execute.scala 117:10]
  wire  _GEN_4594; // @[Execute.scala 117:10]
  wire  _GEN_4595; // @[Execute.scala 117:10]
  wire  _GEN_4596; // @[Execute.scala 117:10]
  wire  _GEN_4597; // @[Execute.scala 117:10]
  wire  _GEN_4598; // @[Execute.scala 117:10]
  wire  _GEN_4599; // @[Execute.scala 117:10]
  wire  _GEN_4600; // @[Execute.scala 117:10]
  wire  _GEN_4601; // @[Execute.scala 117:10]
  wire  _GEN_4602; // @[Execute.scala 117:10]
  wire  _GEN_4603; // @[Execute.scala 117:10]
  wire  _GEN_4604; // @[Execute.scala 117:10]
  wire  _GEN_4605; // @[Execute.scala 117:10]
  wire  _GEN_4606; // @[Execute.scala 117:10]
  wire  _GEN_4607; // @[Execute.scala 117:10]
  wire  _GEN_4608; // @[Execute.scala 117:10]
  wire  _GEN_4609; // @[Execute.scala 117:10]
  wire  _T_441; // @[Execute.scala 117:10]
  wire  _T_442; // @[Execute.scala 117:15]
  wire [5:0] _T_444; // @[Execute.scala 117:37]
  wire [5:0] _T_448; // @[Execute.scala 117:60]
  wire  _GEN_4611; // @[Execute.scala 117:10]
  wire  _GEN_4612; // @[Execute.scala 117:10]
  wire  _GEN_4613; // @[Execute.scala 117:10]
  wire  _GEN_4614; // @[Execute.scala 117:10]
  wire  _GEN_4615; // @[Execute.scala 117:10]
  wire  _GEN_4616; // @[Execute.scala 117:10]
  wire  _GEN_4617; // @[Execute.scala 117:10]
  wire  _GEN_4618; // @[Execute.scala 117:10]
  wire  _GEN_4619; // @[Execute.scala 117:10]
  wire  _GEN_4620; // @[Execute.scala 117:10]
  wire  _GEN_4621; // @[Execute.scala 117:10]
  wire  _GEN_4622; // @[Execute.scala 117:10]
  wire  _GEN_4623; // @[Execute.scala 117:10]
  wire  _GEN_4624; // @[Execute.scala 117:10]
  wire  _GEN_4625; // @[Execute.scala 117:10]
  wire  _GEN_4626; // @[Execute.scala 117:10]
  wire  _GEN_4627; // @[Execute.scala 117:10]
  wire  _GEN_4628; // @[Execute.scala 117:10]
  wire  _GEN_4629; // @[Execute.scala 117:10]
  wire  _GEN_4630; // @[Execute.scala 117:10]
  wire  _GEN_4631; // @[Execute.scala 117:10]
  wire  _GEN_4632; // @[Execute.scala 117:10]
  wire  _GEN_4633; // @[Execute.scala 117:10]
  wire  _GEN_4634; // @[Execute.scala 117:10]
  wire  _GEN_4635; // @[Execute.scala 117:10]
  wire  _GEN_4636; // @[Execute.scala 117:10]
  wire  _GEN_4637; // @[Execute.scala 117:10]
  wire  _GEN_4638; // @[Execute.scala 117:10]
  wire  _GEN_4639; // @[Execute.scala 117:10]
  wire  _GEN_4640; // @[Execute.scala 117:10]
  wire  _GEN_4641; // @[Execute.scala 117:10]
  wire  _GEN_4642; // @[Execute.scala 117:10]
  wire  _GEN_4643; // @[Execute.scala 117:10]
  wire  _GEN_4644; // @[Execute.scala 117:10]
  wire  _GEN_4645; // @[Execute.scala 117:10]
  wire  _GEN_4646; // @[Execute.scala 117:10]
  wire  _GEN_4647; // @[Execute.scala 117:10]
  wire  _GEN_4648; // @[Execute.scala 117:10]
  wire  _GEN_4649; // @[Execute.scala 117:10]
  wire  _GEN_4650; // @[Execute.scala 117:10]
  wire  _GEN_4651; // @[Execute.scala 117:10]
  wire  _GEN_4652; // @[Execute.scala 117:10]
  wire  _GEN_4653; // @[Execute.scala 117:10]
  wire  _GEN_4654; // @[Execute.scala 117:10]
  wire  _GEN_4655; // @[Execute.scala 117:10]
  wire  _GEN_4656; // @[Execute.scala 117:10]
  wire  _GEN_4657; // @[Execute.scala 117:10]
  wire  _GEN_4658; // @[Execute.scala 117:10]
  wire  _GEN_4659; // @[Execute.scala 117:10]
  wire  _GEN_4660; // @[Execute.scala 117:10]
  wire  _GEN_4661; // @[Execute.scala 117:10]
  wire  _GEN_4662; // @[Execute.scala 117:10]
  wire  _GEN_4663; // @[Execute.scala 117:10]
  wire  _GEN_4664; // @[Execute.scala 117:10]
  wire  _GEN_4665; // @[Execute.scala 117:10]
  wire  _GEN_4666; // @[Execute.scala 117:10]
  wire  _GEN_4667; // @[Execute.scala 117:10]
  wire  _GEN_4668; // @[Execute.scala 117:10]
  wire  _GEN_4669; // @[Execute.scala 117:10]
  wire  _GEN_4670; // @[Execute.scala 117:10]
  wire  _GEN_4671; // @[Execute.scala 117:10]
  wire  _GEN_4672; // @[Execute.scala 117:10]
  wire  _GEN_4673; // @[Execute.scala 117:10]
  wire  _GEN_4675; // @[Execute.scala 117:10]
  wire  _GEN_4676; // @[Execute.scala 117:10]
  wire  _GEN_4677; // @[Execute.scala 117:10]
  wire  _GEN_4678; // @[Execute.scala 117:10]
  wire  _GEN_4679; // @[Execute.scala 117:10]
  wire  _GEN_4680; // @[Execute.scala 117:10]
  wire  _GEN_4681; // @[Execute.scala 117:10]
  wire  _GEN_4682; // @[Execute.scala 117:10]
  wire  _GEN_4683; // @[Execute.scala 117:10]
  wire  _GEN_4684; // @[Execute.scala 117:10]
  wire  _GEN_4685; // @[Execute.scala 117:10]
  wire  _GEN_4686; // @[Execute.scala 117:10]
  wire  _GEN_4687; // @[Execute.scala 117:10]
  wire  _GEN_4688; // @[Execute.scala 117:10]
  wire  _GEN_4689; // @[Execute.scala 117:10]
  wire  _GEN_4690; // @[Execute.scala 117:10]
  wire  _GEN_4691; // @[Execute.scala 117:10]
  wire  _GEN_4692; // @[Execute.scala 117:10]
  wire  _GEN_4693; // @[Execute.scala 117:10]
  wire  _GEN_4694; // @[Execute.scala 117:10]
  wire  _GEN_4695; // @[Execute.scala 117:10]
  wire  _GEN_4696; // @[Execute.scala 117:10]
  wire  _GEN_4697; // @[Execute.scala 117:10]
  wire  _GEN_4698; // @[Execute.scala 117:10]
  wire  _GEN_4699; // @[Execute.scala 117:10]
  wire  _GEN_4700; // @[Execute.scala 117:10]
  wire  _GEN_4701; // @[Execute.scala 117:10]
  wire  _GEN_4702; // @[Execute.scala 117:10]
  wire  _GEN_4703; // @[Execute.scala 117:10]
  wire  _GEN_4704; // @[Execute.scala 117:10]
  wire  _GEN_4705; // @[Execute.scala 117:10]
  wire  _GEN_4706; // @[Execute.scala 117:10]
  wire  _GEN_4707; // @[Execute.scala 117:10]
  wire  _GEN_4708; // @[Execute.scala 117:10]
  wire  _GEN_4709; // @[Execute.scala 117:10]
  wire  _GEN_4710; // @[Execute.scala 117:10]
  wire  _GEN_4711; // @[Execute.scala 117:10]
  wire  _GEN_4712; // @[Execute.scala 117:10]
  wire  _GEN_4713; // @[Execute.scala 117:10]
  wire  _GEN_4714; // @[Execute.scala 117:10]
  wire  _GEN_4715; // @[Execute.scala 117:10]
  wire  _GEN_4716; // @[Execute.scala 117:10]
  wire  _GEN_4717; // @[Execute.scala 117:10]
  wire  _GEN_4718; // @[Execute.scala 117:10]
  wire  _GEN_4719; // @[Execute.scala 117:10]
  wire  _GEN_4720; // @[Execute.scala 117:10]
  wire  _GEN_4721; // @[Execute.scala 117:10]
  wire  _GEN_4722; // @[Execute.scala 117:10]
  wire  _GEN_4723; // @[Execute.scala 117:10]
  wire  _GEN_4724; // @[Execute.scala 117:10]
  wire  _GEN_4725; // @[Execute.scala 117:10]
  wire  _GEN_4726; // @[Execute.scala 117:10]
  wire  _GEN_4727; // @[Execute.scala 117:10]
  wire  _GEN_4728; // @[Execute.scala 117:10]
  wire  _GEN_4729; // @[Execute.scala 117:10]
  wire  _GEN_4730; // @[Execute.scala 117:10]
  wire  _GEN_4731; // @[Execute.scala 117:10]
  wire  _GEN_4732; // @[Execute.scala 117:10]
  wire  _GEN_4733; // @[Execute.scala 117:10]
  wire  _GEN_4734; // @[Execute.scala 117:10]
  wire  _GEN_4735; // @[Execute.scala 117:10]
  wire  _GEN_4736; // @[Execute.scala 117:10]
  wire  _GEN_4737; // @[Execute.scala 117:10]
  wire  _T_451; // @[Execute.scala 117:10]
  wire  _T_452; // @[Execute.scala 117:15]
  wire [5:0] _T_454; // @[Execute.scala 117:37]
  wire [5:0] _T_458; // @[Execute.scala 117:60]
  wire  _GEN_4739; // @[Execute.scala 117:10]
  wire  _GEN_4740; // @[Execute.scala 117:10]
  wire  _GEN_4741; // @[Execute.scala 117:10]
  wire  _GEN_4742; // @[Execute.scala 117:10]
  wire  _GEN_4743; // @[Execute.scala 117:10]
  wire  _GEN_4744; // @[Execute.scala 117:10]
  wire  _GEN_4745; // @[Execute.scala 117:10]
  wire  _GEN_4746; // @[Execute.scala 117:10]
  wire  _GEN_4747; // @[Execute.scala 117:10]
  wire  _GEN_4748; // @[Execute.scala 117:10]
  wire  _GEN_4749; // @[Execute.scala 117:10]
  wire  _GEN_4750; // @[Execute.scala 117:10]
  wire  _GEN_4751; // @[Execute.scala 117:10]
  wire  _GEN_4752; // @[Execute.scala 117:10]
  wire  _GEN_4753; // @[Execute.scala 117:10]
  wire  _GEN_4754; // @[Execute.scala 117:10]
  wire  _GEN_4755; // @[Execute.scala 117:10]
  wire  _GEN_4756; // @[Execute.scala 117:10]
  wire  _GEN_4757; // @[Execute.scala 117:10]
  wire  _GEN_4758; // @[Execute.scala 117:10]
  wire  _GEN_4759; // @[Execute.scala 117:10]
  wire  _GEN_4760; // @[Execute.scala 117:10]
  wire  _GEN_4761; // @[Execute.scala 117:10]
  wire  _GEN_4762; // @[Execute.scala 117:10]
  wire  _GEN_4763; // @[Execute.scala 117:10]
  wire  _GEN_4764; // @[Execute.scala 117:10]
  wire  _GEN_4765; // @[Execute.scala 117:10]
  wire  _GEN_4766; // @[Execute.scala 117:10]
  wire  _GEN_4767; // @[Execute.scala 117:10]
  wire  _GEN_4768; // @[Execute.scala 117:10]
  wire  _GEN_4769; // @[Execute.scala 117:10]
  wire  _GEN_4770; // @[Execute.scala 117:10]
  wire  _GEN_4771; // @[Execute.scala 117:10]
  wire  _GEN_4772; // @[Execute.scala 117:10]
  wire  _GEN_4773; // @[Execute.scala 117:10]
  wire  _GEN_4774; // @[Execute.scala 117:10]
  wire  _GEN_4775; // @[Execute.scala 117:10]
  wire  _GEN_4776; // @[Execute.scala 117:10]
  wire  _GEN_4777; // @[Execute.scala 117:10]
  wire  _GEN_4778; // @[Execute.scala 117:10]
  wire  _GEN_4779; // @[Execute.scala 117:10]
  wire  _GEN_4780; // @[Execute.scala 117:10]
  wire  _GEN_4781; // @[Execute.scala 117:10]
  wire  _GEN_4782; // @[Execute.scala 117:10]
  wire  _GEN_4783; // @[Execute.scala 117:10]
  wire  _GEN_4784; // @[Execute.scala 117:10]
  wire  _GEN_4785; // @[Execute.scala 117:10]
  wire  _GEN_4786; // @[Execute.scala 117:10]
  wire  _GEN_4787; // @[Execute.scala 117:10]
  wire  _GEN_4788; // @[Execute.scala 117:10]
  wire  _GEN_4789; // @[Execute.scala 117:10]
  wire  _GEN_4790; // @[Execute.scala 117:10]
  wire  _GEN_4791; // @[Execute.scala 117:10]
  wire  _GEN_4792; // @[Execute.scala 117:10]
  wire  _GEN_4793; // @[Execute.scala 117:10]
  wire  _GEN_4794; // @[Execute.scala 117:10]
  wire  _GEN_4795; // @[Execute.scala 117:10]
  wire  _GEN_4796; // @[Execute.scala 117:10]
  wire  _GEN_4797; // @[Execute.scala 117:10]
  wire  _GEN_4798; // @[Execute.scala 117:10]
  wire  _GEN_4799; // @[Execute.scala 117:10]
  wire  _GEN_4800; // @[Execute.scala 117:10]
  wire  _GEN_4801; // @[Execute.scala 117:10]
  wire  _GEN_4803; // @[Execute.scala 117:10]
  wire  _GEN_4804; // @[Execute.scala 117:10]
  wire  _GEN_4805; // @[Execute.scala 117:10]
  wire  _GEN_4806; // @[Execute.scala 117:10]
  wire  _GEN_4807; // @[Execute.scala 117:10]
  wire  _GEN_4808; // @[Execute.scala 117:10]
  wire  _GEN_4809; // @[Execute.scala 117:10]
  wire  _GEN_4810; // @[Execute.scala 117:10]
  wire  _GEN_4811; // @[Execute.scala 117:10]
  wire  _GEN_4812; // @[Execute.scala 117:10]
  wire  _GEN_4813; // @[Execute.scala 117:10]
  wire  _GEN_4814; // @[Execute.scala 117:10]
  wire  _GEN_4815; // @[Execute.scala 117:10]
  wire  _GEN_4816; // @[Execute.scala 117:10]
  wire  _GEN_4817; // @[Execute.scala 117:10]
  wire  _GEN_4818; // @[Execute.scala 117:10]
  wire  _GEN_4819; // @[Execute.scala 117:10]
  wire  _GEN_4820; // @[Execute.scala 117:10]
  wire  _GEN_4821; // @[Execute.scala 117:10]
  wire  _GEN_4822; // @[Execute.scala 117:10]
  wire  _GEN_4823; // @[Execute.scala 117:10]
  wire  _GEN_4824; // @[Execute.scala 117:10]
  wire  _GEN_4825; // @[Execute.scala 117:10]
  wire  _GEN_4826; // @[Execute.scala 117:10]
  wire  _GEN_4827; // @[Execute.scala 117:10]
  wire  _GEN_4828; // @[Execute.scala 117:10]
  wire  _GEN_4829; // @[Execute.scala 117:10]
  wire  _GEN_4830; // @[Execute.scala 117:10]
  wire  _GEN_4831; // @[Execute.scala 117:10]
  wire  _GEN_4832; // @[Execute.scala 117:10]
  wire  _GEN_4833; // @[Execute.scala 117:10]
  wire  _GEN_4834; // @[Execute.scala 117:10]
  wire  _GEN_4835; // @[Execute.scala 117:10]
  wire  _GEN_4836; // @[Execute.scala 117:10]
  wire  _GEN_4837; // @[Execute.scala 117:10]
  wire  _GEN_4838; // @[Execute.scala 117:10]
  wire  _GEN_4839; // @[Execute.scala 117:10]
  wire  _GEN_4840; // @[Execute.scala 117:10]
  wire  _GEN_4841; // @[Execute.scala 117:10]
  wire  _GEN_4842; // @[Execute.scala 117:10]
  wire  _GEN_4843; // @[Execute.scala 117:10]
  wire  _GEN_4844; // @[Execute.scala 117:10]
  wire  _GEN_4845; // @[Execute.scala 117:10]
  wire  _GEN_4846; // @[Execute.scala 117:10]
  wire  _GEN_4847; // @[Execute.scala 117:10]
  wire  _GEN_4848; // @[Execute.scala 117:10]
  wire  _GEN_4849; // @[Execute.scala 117:10]
  wire  _GEN_4850; // @[Execute.scala 117:10]
  wire  _GEN_4851; // @[Execute.scala 117:10]
  wire  _GEN_4852; // @[Execute.scala 117:10]
  wire  _GEN_4853; // @[Execute.scala 117:10]
  wire  _GEN_4854; // @[Execute.scala 117:10]
  wire  _GEN_4855; // @[Execute.scala 117:10]
  wire  _GEN_4856; // @[Execute.scala 117:10]
  wire  _GEN_4857; // @[Execute.scala 117:10]
  wire  _GEN_4858; // @[Execute.scala 117:10]
  wire  _GEN_4859; // @[Execute.scala 117:10]
  wire  _GEN_4860; // @[Execute.scala 117:10]
  wire  _GEN_4861; // @[Execute.scala 117:10]
  wire  _GEN_4862; // @[Execute.scala 117:10]
  wire  _GEN_4863; // @[Execute.scala 117:10]
  wire  _GEN_4864; // @[Execute.scala 117:10]
  wire  _GEN_4865; // @[Execute.scala 117:10]
  wire  _T_461; // @[Execute.scala 117:10]
  wire  _T_462; // @[Execute.scala 117:15]
  wire [5:0] _T_464; // @[Execute.scala 117:37]
  wire [5:0] _T_468; // @[Execute.scala 117:60]
  wire  _GEN_4867; // @[Execute.scala 117:10]
  wire  _GEN_4868; // @[Execute.scala 117:10]
  wire  _GEN_4869; // @[Execute.scala 117:10]
  wire  _GEN_4870; // @[Execute.scala 117:10]
  wire  _GEN_4871; // @[Execute.scala 117:10]
  wire  _GEN_4872; // @[Execute.scala 117:10]
  wire  _GEN_4873; // @[Execute.scala 117:10]
  wire  _GEN_4874; // @[Execute.scala 117:10]
  wire  _GEN_4875; // @[Execute.scala 117:10]
  wire  _GEN_4876; // @[Execute.scala 117:10]
  wire  _GEN_4877; // @[Execute.scala 117:10]
  wire  _GEN_4878; // @[Execute.scala 117:10]
  wire  _GEN_4879; // @[Execute.scala 117:10]
  wire  _GEN_4880; // @[Execute.scala 117:10]
  wire  _GEN_4881; // @[Execute.scala 117:10]
  wire  _GEN_4882; // @[Execute.scala 117:10]
  wire  _GEN_4883; // @[Execute.scala 117:10]
  wire  _GEN_4884; // @[Execute.scala 117:10]
  wire  _GEN_4885; // @[Execute.scala 117:10]
  wire  _GEN_4886; // @[Execute.scala 117:10]
  wire  _GEN_4887; // @[Execute.scala 117:10]
  wire  _GEN_4888; // @[Execute.scala 117:10]
  wire  _GEN_4889; // @[Execute.scala 117:10]
  wire  _GEN_4890; // @[Execute.scala 117:10]
  wire  _GEN_4891; // @[Execute.scala 117:10]
  wire  _GEN_4892; // @[Execute.scala 117:10]
  wire  _GEN_4893; // @[Execute.scala 117:10]
  wire  _GEN_4894; // @[Execute.scala 117:10]
  wire  _GEN_4895; // @[Execute.scala 117:10]
  wire  _GEN_4896; // @[Execute.scala 117:10]
  wire  _GEN_4897; // @[Execute.scala 117:10]
  wire  _GEN_4898; // @[Execute.scala 117:10]
  wire  _GEN_4899; // @[Execute.scala 117:10]
  wire  _GEN_4900; // @[Execute.scala 117:10]
  wire  _GEN_4901; // @[Execute.scala 117:10]
  wire  _GEN_4902; // @[Execute.scala 117:10]
  wire  _GEN_4903; // @[Execute.scala 117:10]
  wire  _GEN_4904; // @[Execute.scala 117:10]
  wire  _GEN_4905; // @[Execute.scala 117:10]
  wire  _GEN_4906; // @[Execute.scala 117:10]
  wire  _GEN_4907; // @[Execute.scala 117:10]
  wire  _GEN_4908; // @[Execute.scala 117:10]
  wire  _GEN_4909; // @[Execute.scala 117:10]
  wire  _GEN_4910; // @[Execute.scala 117:10]
  wire  _GEN_4911; // @[Execute.scala 117:10]
  wire  _GEN_4912; // @[Execute.scala 117:10]
  wire  _GEN_4913; // @[Execute.scala 117:10]
  wire  _GEN_4914; // @[Execute.scala 117:10]
  wire  _GEN_4915; // @[Execute.scala 117:10]
  wire  _GEN_4916; // @[Execute.scala 117:10]
  wire  _GEN_4917; // @[Execute.scala 117:10]
  wire  _GEN_4918; // @[Execute.scala 117:10]
  wire  _GEN_4919; // @[Execute.scala 117:10]
  wire  _GEN_4920; // @[Execute.scala 117:10]
  wire  _GEN_4921; // @[Execute.scala 117:10]
  wire  _GEN_4922; // @[Execute.scala 117:10]
  wire  _GEN_4923; // @[Execute.scala 117:10]
  wire  _GEN_4924; // @[Execute.scala 117:10]
  wire  _GEN_4925; // @[Execute.scala 117:10]
  wire  _GEN_4926; // @[Execute.scala 117:10]
  wire  _GEN_4927; // @[Execute.scala 117:10]
  wire  _GEN_4928; // @[Execute.scala 117:10]
  wire  _GEN_4929; // @[Execute.scala 117:10]
  wire  _GEN_4931; // @[Execute.scala 117:10]
  wire  _GEN_4932; // @[Execute.scala 117:10]
  wire  _GEN_4933; // @[Execute.scala 117:10]
  wire  _GEN_4934; // @[Execute.scala 117:10]
  wire  _GEN_4935; // @[Execute.scala 117:10]
  wire  _GEN_4936; // @[Execute.scala 117:10]
  wire  _GEN_4937; // @[Execute.scala 117:10]
  wire  _GEN_4938; // @[Execute.scala 117:10]
  wire  _GEN_4939; // @[Execute.scala 117:10]
  wire  _GEN_4940; // @[Execute.scala 117:10]
  wire  _GEN_4941; // @[Execute.scala 117:10]
  wire  _GEN_4942; // @[Execute.scala 117:10]
  wire  _GEN_4943; // @[Execute.scala 117:10]
  wire  _GEN_4944; // @[Execute.scala 117:10]
  wire  _GEN_4945; // @[Execute.scala 117:10]
  wire  _GEN_4946; // @[Execute.scala 117:10]
  wire  _GEN_4947; // @[Execute.scala 117:10]
  wire  _GEN_4948; // @[Execute.scala 117:10]
  wire  _GEN_4949; // @[Execute.scala 117:10]
  wire  _GEN_4950; // @[Execute.scala 117:10]
  wire  _GEN_4951; // @[Execute.scala 117:10]
  wire  _GEN_4952; // @[Execute.scala 117:10]
  wire  _GEN_4953; // @[Execute.scala 117:10]
  wire  _GEN_4954; // @[Execute.scala 117:10]
  wire  _GEN_4955; // @[Execute.scala 117:10]
  wire  _GEN_4956; // @[Execute.scala 117:10]
  wire  _GEN_4957; // @[Execute.scala 117:10]
  wire  _GEN_4958; // @[Execute.scala 117:10]
  wire  _GEN_4959; // @[Execute.scala 117:10]
  wire  _GEN_4960; // @[Execute.scala 117:10]
  wire  _GEN_4961; // @[Execute.scala 117:10]
  wire  _GEN_4962; // @[Execute.scala 117:10]
  wire  _GEN_4963; // @[Execute.scala 117:10]
  wire  _GEN_4964; // @[Execute.scala 117:10]
  wire  _GEN_4965; // @[Execute.scala 117:10]
  wire  _GEN_4966; // @[Execute.scala 117:10]
  wire  _GEN_4967; // @[Execute.scala 117:10]
  wire  _GEN_4968; // @[Execute.scala 117:10]
  wire  _GEN_4969; // @[Execute.scala 117:10]
  wire  _GEN_4970; // @[Execute.scala 117:10]
  wire  _GEN_4971; // @[Execute.scala 117:10]
  wire  _GEN_4972; // @[Execute.scala 117:10]
  wire  _GEN_4973; // @[Execute.scala 117:10]
  wire  _GEN_4974; // @[Execute.scala 117:10]
  wire  _GEN_4975; // @[Execute.scala 117:10]
  wire  _GEN_4976; // @[Execute.scala 117:10]
  wire  _GEN_4977; // @[Execute.scala 117:10]
  wire  _GEN_4978; // @[Execute.scala 117:10]
  wire  _GEN_4979; // @[Execute.scala 117:10]
  wire  _GEN_4980; // @[Execute.scala 117:10]
  wire  _GEN_4981; // @[Execute.scala 117:10]
  wire  _GEN_4982; // @[Execute.scala 117:10]
  wire  _GEN_4983; // @[Execute.scala 117:10]
  wire  _GEN_4984; // @[Execute.scala 117:10]
  wire  _GEN_4985; // @[Execute.scala 117:10]
  wire  _GEN_4986; // @[Execute.scala 117:10]
  wire  _GEN_4987; // @[Execute.scala 117:10]
  wire  _GEN_4988; // @[Execute.scala 117:10]
  wire  _GEN_4989; // @[Execute.scala 117:10]
  wire  _GEN_4990; // @[Execute.scala 117:10]
  wire  _GEN_4991; // @[Execute.scala 117:10]
  wire  _GEN_4992; // @[Execute.scala 117:10]
  wire  _GEN_4993; // @[Execute.scala 117:10]
  wire  _T_471; // @[Execute.scala 117:10]
  wire  _T_472; // @[Execute.scala 117:15]
  wire [5:0] _T_474; // @[Execute.scala 117:37]
  wire [5:0] _T_478; // @[Execute.scala 117:60]
  wire  _GEN_4995; // @[Execute.scala 117:10]
  wire  _GEN_4996; // @[Execute.scala 117:10]
  wire  _GEN_4997; // @[Execute.scala 117:10]
  wire  _GEN_4998; // @[Execute.scala 117:10]
  wire  _GEN_4999; // @[Execute.scala 117:10]
  wire  _GEN_5000; // @[Execute.scala 117:10]
  wire  _GEN_5001; // @[Execute.scala 117:10]
  wire  _GEN_5002; // @[Execute.scala 117:10]
  wire  _GEN_5003; // @[Execute.scala 117:10]
  wire  _GEN_5004; // @[Execute.scala 117:10]
  wire  _GEN_5005; // @[Execute.scala 117:10]
  wire  _GEN_5006; // @[Execute.scala 117:10]
  wire  _GEN_5007; // @[Execute.scala 117:10]
  wire  _GEN_5008; // @[Execute.scala 117:10]
  wire  _GEN_5009; // @[Execute.scala 117:10]
  wire  _GEN_5010; // @[Execute.scala 117:10]
  wire  _GEN_5011; // @[Execute.scala 117:10]
  wire  _GEN_5012; // @[Execute.scala 117:10]
  wire  _GEN_5013; // @[Execute.scala 117:10]
  wire  _GEN_5014; // @[Execute.scala 117:10]
  wire  _GEN_5015; // @[Execute.scala 117:10]
  wire  _GEN_5016; // @[Execute.scala 117:10]
  wire  _GEN_5017; // @[Execute.scala 117:10]
  wire  _GEN_5018; // @[Execute.scala 117:10]
  wire  _GEN_5019; // @[Execute.scala 117:10]
  wire  _GEN_5020; // @[Execute.scala 117:10]
  wire  _GEN_5021; // @[Execute.scala 117:10]
  wire  _GEN_5022; // @[Execute.scala 117:10]
  wire  _GEN_5023; // @[Execute.scala 117:10]
  wire  _GEN_5024; // @[Execute.scala 117:10]
  wire  _GEN_5025; // @[Execute.scala 117:10]
  wire  _GEN_5026; // @[Execute.scala 117:10]
  wire  _GEN_5027; // @[Execute.scala 117:10]
  wire  _GEN_5028; // @[Execute.scala 117:10]
  wire  _GEN_5029; // @[Execute.scala 117:10]
  wire  _GEN_5030; // @[Execute.scala 117:10]
  wire  _GEN_5031; // @[Execute.scala 117:10]
  wire  _GEN_5032; // @[Execute.scala 117:10]
  wire  _GEN_5033; // @[Execute.scala 117:10]
  wire  _GEN_5034; // @[Execute.scala 117:10]
  wire  _GEN_5035; // @[Execute.scala 117:10]
  wire  _GEN_5036; // @[Execute.scala 117:10]
  wire  _GEN_5037; // @[Execute.scala 117:10]
  wire  _GEN_5038; // @[Execute.scala 117:10]
  wire  _GEN_5039; // @[Execute.scala 117:10]
  wire  _GEN_5040; // @[Execute.scala 117:10]
  wire  _GEN_5041; // @[Execute.scala 117:10]
  wire  _GEN_5042; // @[Execute.scala 117:10]
  wire  _GEN_5043; // @[Execute.scala 117:10]
  wire  _GEN_5044; // @[Execute.scala 117:10]
  wire  _GEN_5045; // @[Execute.scala 117:10]
  wire  _GEN_5046; // @[Execute.scala 117:10]
  wire  _GEN_5047; // @[Execute.scala 117:10]
  wire  _GEN_5048; // @[Execute.scala 117:10]
  wire  _GEN_5049; // @[Execute.scala 117:10]
  wire  _GEN_5050; // @[Execute.scala 117:10]
  wire  _GEN_5051; // @[Execute.scala 117:10]
  wire  _GEN_5052; // @[Execute.scala 117:10]
  wire  _GEN_5053; // @[Execute.scala 117:10]
  wire  _GEN_5054; // @[Execute.scala 117:10]
  wire  _GEN_5055; // @[Execute.scala 117:10]
  wire  _GEN_5056; // @[Execute.scala 117:10]
  wire  _GEN_5057; // @[Execute.scala 117:10]
  wire  _GEN_5059; // @[Execute.scala 117:10]
  wire  _GEN_5060; // @[Execute.scala 117:10]
  wire  _GEN_5061; // @[Execute.scala 117:10]
  wire  _GEN_5062; // @[Execute.scala 117:10]
  wire  _GEN_5063; // @[Execute.scala 117:10]
  wire  _GEN_5064; // @[Execute.scala 117:10]
  wire  _GEN_5065; // @[Execute.scala 117:10]
  wire  _GEN_5066; // @[Execute.scala 117:10]
  wire  _GEN_5067; // @[Execute.scala 117:10]
  wire  _GEN_5068; // @[Execute.scala 117:10]
  wire  _GEN_5069; // @[Execute.scala 117:10]
  wire  _GEN_5070; // @[Execute.scala 117:10]
  wire  _GEN_5071; // @[Execute.scala 117:10]
  wire  _GEN_5072; // @[Execute.scala 117:10]
  wire  _GEN_5073; // @[Execute.scala 117:10]
  wire  _GEN_5074; // @[Execute.scala 117:10]
  wire  _GEN_5075; // @[Execute.scala 117:10]
  wire  _GEN_5076; // @[Execute.scala 117:10]
  wire  _GEN_5077; // @[Execute.scala 117:10]
  wire  _GEN_5078; // @[Execute.scala 117:10]
  wire  _GEN_5079; // @[Execute.scala 117:10]
  wire  _GEN_5080; // @[Execute.scala 117:10]
  wire  _GEN_5081; // @[Execute.scala 117:10]
  wire  _GEN_5082; // @[Execute.scala 117:10]
  wire  _GEN_5083; // @[Execute.scala 117:10]
  wire  _GEN_5084; // @[Execute.scala 117:10]
  wire  _GEN_5085; // @[Execute.scala 117:10]
  wire  _GEN_5086; // @[Execute.scala 117:10]
  wire  _GEN_5087; // @[Execute.scala 117:10]
  wire  _GEN_5088; // @[Execute.scala 117:10]
  wire  _GEN_5089; // @[Execute.scala 117:10]
  wire  _GEN_5090; // @[Execute.scala 117:10]
  wire  _GEN_5091; // @[Execute.scala 117:10]
  wire  _GEN_5092; // @[Execute.scala 117:10]
  wire  _GEN_5093; // @[Execute.scala 117:10]
  wire  _GEN_5094; // @[Execute.scala 117:10]
  wire  _GEN_5095; // @[Execute.scala 117:10]
  wire  _GEN_5096; // @[Execute.scala 117:10]
  wire  _GEN_5097; // @[Execute.scala 117:10]
  wire  _GEN_5098; // @[Execute.scala 117:10]
  wire  _GEN_5099; // @[Execute.scala 117:10]
  wire  _GEN_5100; // @[Execute.scala 117:10]
  wire  _GEN_5101; // @[Execute.scala 117:10]
  wire  _GEN_5102; // @[Execute.scala 117:10]
  wire  _GEN_5103; // @[Execute.scala 117:10]
  wire  _GEN_5104; // @[Execute.scala 117:10]
  wire  _GEN_5105; // @[Execute.scala 117:10]
  wire  _GEN_5106; // @[Execute.scala 117:10]
  wire  _GEN_5107; // @[Execute.scala 117:10]
  wire  _GEN_5108; // @[Execute.scala 117:10]
  wire  _GEN_5109; // @[Execute.scala 117:10]
  wire  _GEN_5110; // @[Execute.scala 117:10]
  wire  _GEN_5111; // @[Execute.scala 117:10]
  wire  _GEN_5112; // @[Execute.scala 117:10]
  wire  _GEN_5113; // @[Execute.scala 117:10]
  wire  _GEN_5114; // @[Execute.scala 117:10]
  wire  _GEN_5115; // @[Execute.scala 117:10]
  wire  _GEN_5116; // @[Execute.scala 117:10]
  wire  _GEN_5117; // @[Execute.scala 117:10]
  wire  _GEN_5118; // @[Execute.scala 117:10]
  wire  _GEN_5119; // @[Execute.scala 117:10]
  wire  _GEN_5120; // @[Execute.scala 117:10]
  wire  _GEN_5121; // @[Execute.scala 117:10]
  wire  _T_481; // @[Execute.scala 117:10]
  wire  _T_482; // @[Execute.scala 117:15]
  wire [5:0] _T_484; // @[Execute.scala 117:37]
  wire [5:0] _T_488; // @[Execute.scala 117:60]
  wire  _GEN_5123; // @[Execute.scala 117:10]
  wire  _GEN_5124; // @[Execute.scala 117:10]
  wire  _GEN_5125; // @[Execute.scala 117:10]
  wire  _GEN_5126; // @[Execute.scala 117:10]
  wire  _GEN_5127; // @[Execute.scala 117:10]
  wire  _GEN_5128; // @[Execute.scala 117:10]
  wire  _GEN_5129; // @[Execute.scala 117:10]
  wire  _GEN_5130; // @[Execute.scala 117:10]
  wire  _GEN_5131; // @[Execute.scala 117:10]
  wire  _GEN_5132; // @[Execute.scala 117:10]
  wire  _GEN_5133; // @[Execute.scala 117:10]
  wire  _GEN_5134; // @[Execute.scala 117:10]
  wire  _GEN_5135; // @[Execute.scala 117:10]
  wire  _GEN_5136; // @[Execute.scala 117:10]
  wire  _GEN_5137; // @[Execute.scala 117:10]
  wire  _GEN_5138; // @[Execute.scala 117:10]
  wire  _GEN_5139; // @[Execute.scala 117:10]
  wire  _GEN_5140; // @[Execute.scala 117:10]
  wire  _GEN_5141; // @[Execute.scala 117:10]
  wire  _GEN_5142; // @[Execute.scala 117:10]
  wire  _GEN_5143; // @[Execute.scala 117:10]
  wire  _GEN_5144; // @[Execute.scala 117:10]
  wire  _GEN_5145; // @[Execute.scala 117:10]
  wire  _GEN_5146; // @[Execute.scala 117:10]
  wire  _GEN_5147; // @[Execute.scala 117:10]
  wire  _GEN_5148; // @[Execute.scala 117:10]
  wire  _GEN_5149; // @[Execute.scala 117:10]
  wire  _GEN_5150; // @[Execute.scala 117:10]
  wire  _GEN_5151; // @[Execute.scala 117:10]
  wire  _GEN_5152; // @[Execute.scala 117:10]
  wire  _GEN_5153; // @[Execute.scala 117:10]
  wire  _GEN_5154; // @[Execute.scala 117:10]
  wire  _GEN_5155; // @[Execute.scala 117:10]
  wire  _GEN_5156; // @[Execute.scala 117:10]
  wire  _GEN_5157; // @[Execute.scala 117:10]
  wire  _GEN_5158; // @[Execute.scala 117:10]
  wire  _GEN_5159; // @[Execute.scala 117:10]
  wire  _GEN_5160; // @[Execute.scala 117:10]
  wire  _GEN_5161; // @[Execute.scala 117:10]
  wire  _GEN_5162; // @[Execute.scala 117:10]
  wire  _GEN_5163; // @[Execute.scala 117:10]
  wire  _GEN_5164; // @[Execute.scala 117:10]
  wire  _GEN_5165; // @[Execute.scala 117:10]
  wire  _GEN_5166; // @[Execute.scala 117:10]
  wire  _GEN_5167; // @[Execute.scala 117:10]
  wire  _GEN_5168; // @[Execute.scala 117:10]
  wire  _GEN_5169; // @[Execute.scala 117:10]
  wire  _GEN_5170; // @[Execute.scala 117:10]
  wire  _GEN_5171; // @[Execute.scala 117:10]
  wire  _GEN_5172; // @[Execute.scala 117:10]
  wire  _GEN_5173; // @[Execute.scala 117:10]
  wire  _GEN_5174; // @[Execute.scala 117:10]
  wire  _GEN_5175; // @[Execute.scala 117:10]
  wire  _GEN_5176; // @[Execute.scala 117:10]
  wire  _GEN_5177; // @[Execute.scala 117:10]
  wire  _GEN_5178; // @[Execute.scala 117:10]
  wire  _GEN_5179; // @[Execute.scala 117:10]
  wire  _GEN_5180; // @[Execute.scala 117:10]
  wire  _GEN_5181; // @[Execute.scala 117:10]
  wire  _GEN_5182; // @[Execute.scala 117:10]
  wire  _GEN_5183; // @[Execute.scala 117:10]
  wire  _GEN_5184; // @[Execute.scala 117:10]
  wire  _GEN_5185; // @[Execute.scala 117:10]
  wire  _GEN_5187; // @[Execute.scala 117:10]
  wire  _GEN_5188; // @[Execute.scala 117:10]
  wire  _GEN_5189; // @[Execute.scala 117:10]
  wire  _GEN_5190; // @[Execute.scala 117:10]
  wire  _GEN_5191; // @[Execute.scala 117:10]
  wire  _GEN_5192; // @[Execute.scala 117:10]
  wire  _GEN_5193; // @[Execute.scala 117:10]
  wire  _GEN_5194; // @[Execute.scala 117:10]
  wire  _GEN_5195; // @[Execute.scala 117:10]
  wire  _GEN_5196; // @[Execute.scala 117:10]
  wire  _GEN_5197; // @[Execute.scala 117:10]
  wire  _GEN_5198; // @[Execute.scala 117:10]
  wire  _GEN_5199; // @[Execute.scala 117:10]
  wire  _GEN_5200; // @[Execute.scala 117:10]
  wire  _GEN_5201; // @[Execute.scala 117:10]
  wire  _GEN_5202; // @[Execute.scala 117:10]
  wire  _GEN_5203; // @[Execute.scala 117:10]
  wire  _GEN_5204; // @[Execute.scala 117:10]
  wire  _GEN_5205; // @[Execute.scala 117:10]
  wire  _GEN_5206; // @[Execute.scala 117:10]
  wire  _GEN_5207; // @[Execute.scala 117:10]
  wire  _GEN_5208; // @[Execute.scala 117:10]
  wire  _GEN_5209; // @[Execute.scala 117:10]
  wire  _GEN_5210; // @[Execute.scala 117:10]
  wire  _GEN_5211; // @[Execute.scala 117:10]
  wire  _GEN_5212; // @[Execute.scala 117:10]
  wire  _GEN_5213; // @[Execute.scala 117:10]
  wire  _GEN_5214; // @[Execute.scala 117:10]
  wire  _GEN_5215; // @[Execute.scala 117:10]
  wire  _GEN_5216; // @[Execute.scala 117:10]
  wire  _GEN_5217; // @[Execute.scala 117:10]
  wire  _GEN_5218; // @[Execute.scala 117:10]
  wire  _GEN_5219; // @[Execute.scala 117:10]
  wire  _GEN_5220; // @[Execute.scala 117:10]
  wire  _GEN_5221; // @[Execute.scala 117:10]
  wire  _GEN_5222; // @[Execute.scala 117:10]
  wire  _GEN_5223; // @[Execute.scala 117:10]
  wire  _GEN_5224; // @[Execute.scala 117:10]
  wire  _GEN_5225; // @[Execute.scala 117:10]
  wire  _GEN_5226; // @[Execute.scala 117:10]
  wire  _GEN_5227; // @[Execute.scala 117:10]
  wire  _GEN_5228; // @[Execute.scala 117:10]
  wire  _GEN_5229; // @[Execute.scala 117:10]
  wire  _GEN_5230; // @[Execute.scala 117:10]
  wire  _GEN_5231; // @[Execute.scala 117:10]
  wire  _GEN_5232; // @[Execute.scala 117:10]
  wire  _GEN_5233; // @[Execute.scala 117:10]
  wire  _GEN_5234; // @[Execute.scala 117:10]
  wire  _GEN_5235; // @[Execute.scala 117:10]
  wire  _GEN_5236; // @[Execute.scala 117:10]
  wire  _GEN_5237; // @[Execute.scala 117:10]
  wire  _GEN_5238; // @[Execute.scala 117:10]
  wire  _GEN_5239; // @[Execute.scala 117:10]
  wire  _GEN_5240; // @[Execute.scala 117:10]
  wire  _GEN_5241; // @[Execute.scala 117:10]
  wire  _GEN_5242; // @[Execute.scala 117:10]
  wire  _GEN_5243; // @[Execute.scala 117:10]
  wire  _GEN_5244; // @[Execute.scala 117:10]
  wire  _GEN_5245; // @[Execute.scala 117:10]
  wire  _GEN_5246; // @[Execute.scala 117:10]
  wire  _GEN_5247; // @[Execute.scala 117:10]
  wire  _GEN_5248; // @[Execute.scala 117:10]
  wire  _GEN_5249; // @[Execute.scala 117:10]
  wire  _T_491; // @[Execute.scala 117:10]
  wire  _T_492; // @[Execute.scala 117:15]
  wire [5:0] _T_494; // @[Execute.scala 117:37]
  wire [5:0] _T_498; // @[Execute.scala 117:60]
  wire  _GEN_5251; // @[Execute.scala 117:10]
  wire  _GEN_5252; // @[Execute.scala 117:10]
  wire  _GEN_5253; // @[Execute.scala 117:10]
  wire  _GEN_5254; // @[Execute.scala 117:10]
  wire  _GEN_5255; // @[Execute.scala 117:10]
  wire  _GEN_5256; // @[Execute.scala 117:10]
  wire  _GEN_5257; // @[Execute.scala 117:10]
  wire  _GEN_5258; // @[Execute.scala 117:10]
  wire  _GEN_5259; // @[Execute.scala 117:10]
  wire  _GEN_5260; // @[Execute.scala 117:10]
  wire  _GEN_5261; // @[Execute.scala 117:10]
  wire  _GEN_5262; // @[Execute.scala 117:10]
  wire  _GEN_5263; // @[Execute.scala 117:10]
  wire  _GEN_5264; // @[Execute.scala 117:10]
  wire  _GEN_5265; // @[Execute.scala 117:10]
  wire  _GEN_5266; // @[Execute.scala 117:10]
  wire  _GEN_5267; // @[Execute.scala 117:10]
  wire  _GEN_5268; // @[Execute.scala 117:10]
  wire  _GEN_5269; // @[Execute.scala 117:10]
  wire  _GEN_5270; // @[Execute.scala 117:10]
  wire  _GEN_5271; // @[Execute.scala 117:10]
  wire  _GEN_5272; // @[Execute.scala 117:10]
  wire  _GEN_5273; // @[Execute.scala 117:10]
  wire  _GEN_5274; // @[Execute.scala 117:10]
  wire  _GEN_5275; // @[Execute.scala 117:10]
  wire  _GEN_5276; // @[Execute.scala 117:10]
  wire  _GEN_5277; // @[Execute.scala 117:10]
  wire  _GEN_5278; // @[Execute.scala 117:10]
  wire  _GEN_5279; // @[Execute.scala 117:10]
  wire  _GEN_5280; // @[Execute.scala 117:10]
  wire  _GEN_5281; // @[Execute.scala 117:10]
  wire  _GEN_5282; // @[Execute.scala 117:10]
  wire  _GEN_5283; // @[Execute.scala 117:10]
  wire  _GEN_5284; // @[Execute.scala 117:10]
  wire  _GEN_5285; // @[Execute.scala 117:10]
  wire  _GEN_5286; // @[Execute.scala 117:10]
  wire  _GEN_5287; // @[Execute.scala 117:10]
  wire  _GEN_5288; // @[Execute.scala 117:10]
  wire  _GEN_5289; // @[Execute.scala 117:10]
  wire  _GEN_5290; // @[Execute.scala 117:10]
  wire  _GEN_5291; // @[Execute.scala 117:10]
  wire  _GEN_5292; // @[Execute.scala 117:10]
  wire  _GEN_5293; // @[Execute.scala 117:10]
  wire  _GEN_5294; // @[Execute.scala 117:10]
  wire  _GEN_5295; // @[Execute.scala 117:10]
  wire  _GEN_5296; // @[Execute.scala 117:10]
  wire  _GEN_5297; // @[Execute.scala 117:10]
  wire  _GEN_5298; // @[Execute.scala 117:10]
  wire  _GEN_5299; // @[Execute.scala 117:10]
  wire  _GEN_5300; // @[Execute.scala 117:10]
  wire  _GEN_5301; // @[Execute.scala 117:10]
  wire  _GEN_5302; // @[Execute.scala 117:10]
  wire  _GEN_5303; // @[Execute.scala 117:10]
  wire  _GEN_5304; // @[Execute.scala 117:10]
  wire  _GEN_5305; // @[Execute.scala 117:10]
  wire  _GEN_5306; // @[Execute.scala 117:10]
  wire  _GEN_5307; // @[Execute.scala 117:10]
  wire  _GEN_5308; // @[Execute.scala 117:10]
  wire  _GEN_5309; // @[Execute.scala 117:10]
  wire  _GEN_5310; // @[Execute.scala 117:10]
  wire  _GEN_5311; // @[Execute.scala 117:10]
  wire  _GEN_5312; // @[Execute.scala 117:10]
  wire  _GEN_5313; // @[Execute.scala 117:10]
  wire  _GEN_5315; // @[Execute.scala 117:10]
  wire  _GEN_5316; // @[Execute.scala 117:10]
  wire  _GEN_5317; // @[Execute.scala 117:10]
  wire  _GEN_5318; // @[Execute.scala 117:10]
  wire  _GEN_5319; // @[Execute.scala 117:10]
  wire  _GEN_5320; // @[Execute.scala 117:10]
  wire  _GEN_5321; // @[Execute.scala 117:10]
  wire  _GEN_5322; // @[Execute.scala 117:10]
  wire  _GEN_5323; // @[Execute.scala 117:10]
  wire  _GEN_5324; // @[Execute.scala 117:10]
  wire  _GEN_5325; // @[Execute.scala 117:10]
  wire  _GEN_5326; // @[Execute.scala 117:10]
  wire  _GEN_5327; // @[Execute.scala 117:10]
  wire  _GEN_5328; // @[Execute.scala 117:10]
  wire  _GEN_5329; // @[Execute.scala 117:10]
  wire  _GEN_5330; // @[Execute.scala 117:10]
  wire  _GEN_5331; // @[Execute.scala 117:10]
  wire  _GEN_5332; // @[Execute.scala 117:10]
  wire  _GEN_5333; // @[Execute.scala 117:10]
  wire  _GEN_5334; // @[Execute.scala 117:10]
  wire  _GEN_5335; // @[Execute.scala 117:10]
  wire  _GEN_5336; // @[Execute.scala 117:10]
  wire  _GEN_5337; // @[Execute.scala 117:10]
  wire  _GEN_5338; // @[Execute.scala 117:10]
  wire  _GEN_5339; // @[Execute.scala 117:10]
  wire  _GEN_5340; // @[Execute.scala 117:10]
  wire  _GEN_5341; // @[Execute.scala 117:10]
  wire  _GEN_5342; // @[Execute.scala 117:10]
  wire  _GEN_5343; // @[Execute.scala 117:10]
  wire  _GEN_5344; // @[Execute.scala 117:10]
  wire  _GEN_5345; // @[Execute.scala 117:10]
  wire  _GEN_5346; // @[Execute.scala 117:10]
  wire  _GEN_5347; // @[Execute.scala 117:10]
  wire  _GEN_5348; // @[Execute.scala 117:10]
  wire  _GEN_5349; // @[Execute.scala 117:10]
  wire  _GEN_5350; // @[Execute.scala 117:10]
  wire  _GEN_5351; // @[Execute.scala 117:10]
  wire  _GEN_5352; // @[Execute.scala 117:10]
  wire  _GEN_5353; // @[Execute.scala 117:10]
  wire  _GEN_5354; // @[Execute.scala 117:10]
  wire  _GEN_5355; // @[Execute.scala 117:10]
  wire  _GEN_5356; // @[Execute.scala 117:10]
  wire  _GEN_5357; // @[Execute.scala 117:10]
  wire  _GEN_5358; // @[Execute.scala 117:10]
  wire  _GEN_5359; // @[Execute.scala 117:10]
  wire  _GEN_5360; // @[Execute.scala 117:10]
  wire  _GEN_5361; // @[Execute.scala 117:10]
  wire  _GEN_5362; // @[Execute.scala 117:10]
  wire  _GEN_5363; // @[Execute.scala 117:10]
  wire  _GEN_5364; // @[Execute.scala 117:10]
  wire  _GEN_5365; // @[Execute.scala 117:10]
  wire  _GEN_5366; // @[Execute.scala 117:10]
  wire  _GEN_5367; // @[Execute.scala 117:10]
  wire  _GEN_5368; // @[Execute.scala 117:10]
  wire  _GEN_5369; // @[Execute.scala 117:10]
  wire  _GEN_5370; // @[Execute.scala 117:10]
  wire  _GEN_5371; // @[Execute.scala 117:10]
  wire  _GEN_5372; // @[Execute.scala 117:10]
  wire  _GEN_5373; // @[Execute.scala 117:10]
  wire  _GEN_5374; // @[Execute.scala 117:10]
  wire  _GEN_5375; // @[Execute.scala 117:10]
  wire  _GEN_5376; // @[Execute.scala 117:10]
  wire  _GEN_5377; // @[Execute.scala 117:10]
  wire  _T_501; // @[Execute.scala 117:10]
  wire  _T_502; // @[Execute.scala 117:15]
  wire [5:0] _T_504; // @[Execute.scala 117:37]
  wire [5:0] _T_508; // @[Execute.scala 117:60]
  wire  _GEN_5379; // @[Execute.scala 117:10]
  wire  _GEN_5380; // @[Execute.scala 117:10]
  wire  _GEN_5381; // @[Execute.scala 117:10]
  wire  _GEN_5382; // @[Execute.scala 117:10]
  wire  _GEN_5383; // @[Execute.scala 117:10]
  wire  _GEN_5384; // @[Execute.scala 117:10]
  wire  _GEN_5385; // @[Execute.scala 117:10]
  wire  _GEN_5386; // @[Execute.scala 117:10]
  wire  _GEN_5387; // @[Execute.scala 117:10]
  wire  _GEN_5388; // @[Execute.scala 117:10]
  wire  _GEN_5389; // @[Execute.scala 117:10]
  wire  _GEN_5390; // @[Execute.scala 117:10]
  wire  _GEN_5391; // @[Execute.scala 117:10]
  wire  _GEN_5392; // @[Execute.scala 117:10]
  wire  _GEN_5393; // @[Execute.scala 117:10]
  wire  _GEN_5394; // @[Execute.scala 117:10]
  wire  _GEN_5395; // @[Execute.scala 117:10]
  wire  _GEN_5396; // @[Execute.scala 117:10]
  wire  _GEN_5397; // @[Execute.scala 117:10]
  wire  _GEN_5398; // @[Execute.scala 117:10]
  wire  _GEN_5399; // @[Execute.scala 117:10]
  wire  _GEN_5400; // @[Execute.scala 117:10]
  wire  _GEN_5401; // @[Execute.scala 117:10]
  wire  _GEN_5402; // @[Execute.scala 117:10]
  wire  _GEN_5403; // @[Execute.scala 117:10]
  wire  _GEN_5404; // @[Execute.scala 117:10]
  wire  _GEN_5405; // @[Execute.scala 117:10]
  wire  _GEN_5406; // @[Execute.scala 117:10]
  wire  _GEN_5407; // @[Execute.scala 117:10]
  wire  _GEN_5408; // @[Execute.scala 117:10]
  wire  _GEN_5409; // @[Execute.scala 117:10]
  wire  _GEN_5410; // @[Execute.scala 117:10]
  wire  _GEN_5411; // @[Execute.scala 117:10]
  wire  _GEN_5412; // @[Execute.scala 117:10]
  wire  _GEN_5413; // @[Execute.scala 117:10]
  wire  _GEN_5414; // @[Execute.scala 117:10]
  wire  _GEN_5415; // @[Execute.scala 117:10]
  wire  _GEN_5416; // @[Execute.scala 117:10]
  wire  _GEN_5417; // @[Execute.scala 117:10]
  wire  _GEN_5418; // @[Execute.scala 117:10]
  wire  _GEN_5419; // @[Execute.scala 117:10]
  wire  _GEN_5420; // @[Execute.scala 117:10]
  wire  _GEN_5421; // @[Execute.scala 117:10]
  wire  _GEN_5422; // @[Execute.scala 117:10]
  wire  _GEN_5423; // @[Execute.scala 117:10]
  wire  _GEN_5424; // @[Execute.scala 117:10]
  wire  _GEN_5425; // @[Execute.scala 117:10]
  wire  _GEN_5426; // @[Execute.scala 117:10]
  wire  _GEN_5427; // @[Execute.scala 117:10]
  wire  _GEN_5428; // @[Execute.scala 117:10]
  wire  _GEN_5429; // @[Execute.scala 117:10]
  wire  _GEN_5430; // @[Execute.scala 117:10]
  wire  _GEN_5431; // @[Execute.scala 117:10]
  wire  _GEN_5432; // @[Execute.scala 117:10]
  wire  _GEN_5433; // @[Execute.scala 117:10]
  wire  _GEN_5434; // @[Execute.scala 117:10]
  wire  _GEN_5435; // @[Execute.scala 117:10]
  wire  _GEN_5436; // @[Execute.scala 117:10]
  wire  _GEN_5437; // @[Execute.scala 117:10]
  wire  _GEN_5438; // @[Execute.scala 117:10]
  wire  _GEN_5439; // @[Execute.scala 117:10]
  wire  _GEN_5440; // @[Execute.scala 117:10]
  wire  _GEN_5441; // @[Execute.scala 117:10]
  wire  _GEN_5443; // @[Execute.scala 117:10]
  wire  _GEN_5444; // @[Execute.scala 117:10]
  wire  _GEN_5445; // @[Execute.scala 117:10]
  wire  _GEN_5446; // @[Execute.scala 117:10]
  wire  _GEN_5447; // @[Execute.scala 117:10]
  wire  _GEN_5448; // @[Execute.scala 117:10]
  wire  _GEN_5449; // @[Execute.scala 117:10]
  wire  _GEN_5450; // @[Execute.scala 117:10]
  wire  _GEN_5451; // @[Execute.scala 117:10]
  wire  _GEN_5452; // @[Execute.scala 117:10]
  wire  _GEN_5453; // @[Execute.scala 117:10]
  wire  _GEN_5454; // @[Execute.scala 117:10]
  wire  _GEN_5455; // @[Execute.scala 117:10]
  wire  _GEN_5456; // @[Execute.scala 117:10]
  wire  _GEN_5457; // @[Execute.scala 117:10]
  wire  _GEN_5458; // @[Execute.scala 117:10]
  wire  _GEN_5459; // @[Execute.scala 117:10]
  wire  _GEN_5460; // @[Execute.scala 117:10]
  wire  _GEN_5461; // @[Execute.scala 117:10]
  wire  _GEN_5462; // @[Execute.scala 117:10]
  wire  _GEN_5463; // @[Execute.scala 117:10]
  wire  _GEN_5464; // @[Execute.scala 117:10]
  wire  _GEN_5465; // @[Execute.scala 117:10]
  wire  _GEN_5466; // @[Execute.scala 117:10]
  wire  _GEN_5467; // @[Execute.scala 117:10]
  wire  _GEN_5468; // @[Execute.scala 117:10]
  wire  _GEN_5469; // @[Execute.scala 117:10]
  wire  _GEN_5470; // @[Execute.scala 117:10]
  wire  _GEN_5471; // @[Execute.scala 117:10]
  wire  _GEN_5472; // @[Execute.scala 117:10]
  wire  _GEN_5473; // @[Execute.scala 117:10]
  wire  _GEN_5474; // @[Execute.scala 117:10]
  wire  _GEN_5475; // @[Execute.scala 117:10]
  wire  _GEN_5476; // @[Execute.scala 117:10]
  wire  _GEN_5477; // @[Execute.scala 117:10]
  wire  _GEN_5478; // @[Execute.scala 117:10]
  wire  _GEN_5479; // @[Execute.scala 117:10]
  wire  _GEN_5480; // @[Execute.scala 117:10]
  wire  _GEN_5481; // @[Execute.scala 117:10]
  wire  _GEN_5482; // @[Execute.scala 117:10]
  wire  _GEN_5483; // @[Execute.scala 117:10]
  wire  _GEN_5484; // @[Execute.scala 117:10]
  wire  _GEN_5485; // @[Execute.scala 117:10]
  wire  _GEN_5486; // @[Execute.scala 117:10]
  wire  _GEN_5487; // @[Execute.scala 117:10]
  wire  _GEN_5488; // @[Execute.scala 117:10]
  wire  _GEN_5489; // @[Execute.scala 117:10]
  wire  _GEN_5490; // @[Execute.scala 117:10]
  wire  _GEN_5491; // @[Execute.scala 117:10]
  wire  _GEN_5492; // @[Execute.scala 117:10]
  wire  _GEN_5493; // @[Execute.scala 117:10]
  wire  _GEN_5494; // @[Execute.scala 117:10]
  wire  _GEN_5495; // @[Execute.scala 117:10]
  wire  _GEN_5496; // @[Execute.scala 117:10]
  wire  _GEN_5497; // @[Execute.scala 117:10]
  wire  _GEN_5498; // @[Execute.scala 117:10]
  wire  _GEN_5499; // @[Execute.scala 117:10]
  wire  _GEN_5500; // @[Execute.scala 117:10]
  wire  _GEN_5501; // @[Execute.scala 117:10]
  wire  _GEN_5502; // @[Execute.scala 117:10]
  wire  _GEN_5503; // @[Execute.scala 117:10]
  wire  _GEN_5504; // @[Execute.scala 117:10]
  wire  _GEN_5505; // @[Execute.scala 117:10]
  wire  _T_511; // @[Execute.scala 117:10]
  wire  _T_512; // @[Execute.scala 117:15]
  wire [5:0] _T_514; // @[Execute.scala 117:37]
  wire [5:0] _T_518; // @[Execute.scala 117:60]
  wire  _GEN_5507; // @[Execute.scala 117:10]
  wire  _GEN_5508; // @[Execute.scala 117:10]
  wire  _GEN_5509; // @[Execute.scala 117:10]
  wire  _GEN_5510; // @[Execute.scala 117:10]
  wire  _GEN_5511; // @[Execute.scala 117:10]
  wire  _GEN_5512; // @[Execute.scala 117:10]
  wire  _GEN_5513; // @[Execute.scala 117:10]
  wire  _GEN_5514; // @[Execute.scala 117:10]
  wire  _GEN_5515; // @[Execute.scala 117:10]
  wire  _GEN_5516; // @[Execute.scala 117:10]
  wire  _GEN_5517; // @[Execute.scala 117:10]
  wire  _GEN_5518; // @[Execute.scala 117:10]
  wire  _GEN_5519; // @[Execute.scala 117:10]
  wire  _GEN_5520; // @[Execute.scala 117:10]
  wire  _GEN_5521; // @[Execute.scala 117:10]
  wire  _GEN_5522; // @[Execute.scala 117:10]
  wire  _GEN_5523; // @[Execute.scala 117:10]
  wire  _GEN_5524; // @[Execute.scala 117:10]
  wire  _GEN_5525; // @[Execute.scala 117:10]
  wire  _GEN_5526; // @[Execute.scala 117:10]
  wire  _GEN_5527; // @[Execute.scala 117:10]
  wire  _GEN_5528; // @[Execute.scala 117:10]
  wire  _GEN_5529; // @[Execute.scala 117:10]
  wire  _GEN_5530; // @[Execute.scala 117:10]
  wire  _GEN_5531; // @[Execute.scala 117:10]
  wire  _GEN_5532; // @[Execute.scala 117:10]
  wire  _GEN_5533; // @[Execute.scala 117:10]
  wire  _GEN_5534; // @[Execute.scala 117:10]
  wire  _GEN_5535; // @[Execute.scala 117:10]
  wire  _GEN_5536; // @[Execute.scala 117:10]
  wire  _GEN_5537; // @[Execute.scala 117:10]
  wire  _GEN_5538; // @[Execute.scala 117:10]
  wire  _GEN_5539; // @[Execute.scala 117:10]
  wire  _GEN_5540; // @[Execute.scala 117:10]
  wire  _GEN_5541; // @[Execute.scala 117:10]
  wire  _GEN_5542; // @[Execute.scala 117:10]
  wire  _GEN_5543; // @[Execute.scala 117:10]
  wire  _GEN_5544; // @[Execute.scala 117:10]
  wire  _GEN_5545; // @[Execute.scala 117:10]
  wire  _GEN_5546; // @[Execute.scala 117:10]
  wire  _GEN_5547; // @[Execute.scala 117:10]
  wire  _GEN_5548; // @[Execute.scala 117:10]
  wire  _GEN_5549; // @[Execute.scala 117:10]
  wire  _GEN_5550; // @[Execute.scala 117:10]
  wire  _GEN_5551; // @[Execute.scala 117:10]
  wire  _GEN_5552; // @[Execute.scala 117:10]
  wire  _GEN_5553; // @[Execute.scala 117:10]
  wire  _GEN_5554; // @[Execute.scala 117:10]
  wire  _GEN_5555; // @[Execute.scala 117:10]
  wire  _GEN_5556; // @[Execute.scala 117:10]
  wire  _GEN_5557; // @[Execute.scala 117:10]
  wire  _GEN_5558; // @[Execute.scala 117:10]
  wire  _GEN_5559; // @[Execute.scala 117:10]
  wire  _GEN_5560; // @[Execute.scala 117:10]
  wire  _GEN_5561; // @[Execute.scala 117:10]
  wire  _GEN_5562; // @[Execute.scala 117:10]
  wire  _GEN_5563; // @[Execute.scala 117:10]
  wire  _GEN_5564; // @[Execute.scala 117:10]
  wire  _GEN_5565; // @[Execute.scala 117:10]
  wire  _GEN_5566; // @[Execute.scala 117:10]
  wire  _GEN_5567; // @[Execute.scala 117:10]
  wire  _GEN_5568; // @[Execute.scala 117:10]
  wire  _GEN_5569; // @[Execute.scala 117:10]
  wire  _GEN_5571; // @[Execute.scala 117:10]
  wire  _GEN_5572; // @[Execute.scala 117:10]
  wire  _GEN_5573; // @[Execute.scala 117:10]
  wire  _GEN_5574; // @[Execute.scala 117:10]
  wire  _GEN_5575; // @[Execute.scala 117:10]
  wire  _GEN_5576; // @[Execute.scala 117:10]
  wire  _GEN_5577; // @[Execute.scala 117:10]
  wire  _GEN_5578; // @[Execute.scala 117:10]
  wire  _GEN_5579; // @[Execute.scala 117:10]
  wire  _GEN_5580; // @[Execute.scala 117:10]
  wire  _GEN_5581; // @[Execute.scala 117:10]
  wire  _GEN_5582; // @[Execute.scala 117:10]
  wire  _GEN_5583; // @[Execute.scala 117:10]
  wire  _GEN_5584; // @[Execute.scala 117:10]
  wire  _GEN_5585; // @[Execute.scala 117:10]
  wire  _GEN_5586; // @[Execute.scala 117:10]
  wire  _GEN_5587; // @[Execute.scala 117:10]
  wire  _GEN_5588; // @[Execute.scala 117:10]
  wire  _GEN_5589; // @[Execute.scala 117:10]
  wire  _GEN_5590; // @[Execute.scala 117:10]
  wire  _GEN_5591; // @[Execute.scala 117:10]
  wire  _GEN_5592; // @[Execute.scala 117:10]
  wire  _GEN_5593; // @[Execute.scala 117:10]
  wire  _GEN_5594; // @[Execute.scala 117:10]
  wire  _GEN_5595; // @[Execute.scala 117:10]
  wire  _GEN_5596; // @[Execute.scala 117:10]
  wire  _GEN_5597; // @[Execute.scala 117:10]
  wire  _GEN_5598; // @[Execute.scala 117:10]
  wire  _GEN_5599; // @[Execute.scala 117:10]
  wire  _GEN_5600; // @[Execute.scala 117:10]
  wire  _GEN_5601; // @[Execute.scala 117:10]
  wire  _GEN_5602; // @[Execute.scala 117:10]
  wire  _GEN_5603; // @[Execute.scala 117:10]
  wire  _GEN_5604; // @[Execute.scala 117:10]
  wire  _GEN_5605; // @[Execute.scala 117:10]
  wire  _GEN_5606; // @[Execute.scala 117:10]
  wire  _GEN_5607; // @[Execute.scala 117:10]
  wire  _GEN_5608; // @[Execute.scala 117:10]
  wire  _GEN_5609; // @[Execute.scala 117:10]
  wire  _GEN_5610; // @[Execute.scala 117:10]
  wire  _GEN_5611; // @[Execute.scala 117:10]
  wire  _GEN_5612; // @[Execute.scala 117:10]
  wire  _GEN_5613; // @[Execute.scala 117:10]
  wire  _GEN_5614; // @[Execute.scala 117:10]
  wire  _GEN_5615; // @[Execute.scala 117:10]
  wire  _GEN_5616; // @[Execute.scala 117:10]
  wire  _GEN_5617; // @[Execute.scala 117:10]
  wire  _GEN_5618; // @[Execute.scala 117:10]
  wire  _GEN_5619; // @[Execute.scala 117:10]
  wire  _GEN_5620; // @[Execute.scala 117:10]
  wire  _GEN_5621; // @[Execute.scala 117:10]
  wire  _GEN_5622; // @[Execute.scala 117:10]
  wire  _GEN_5623; // @[Execute.scala 117:10]
  wire  _GEN_5624; // @[Execute.scala 117:10]
  wire  _GEN_5625; // @[Execute.scala 117:10]
  wire  _GEN_5626; // @[Execute.scala 117:10]
  wire  _GEN_5627; // @[Execute.scala 117:10]
  wire  _GEN_5628; // @[Execute.scala 117:10]
  wire  _GEN_5629; // @[Execute.scala 117:10]
  wire  _GEN_5630; // @[Execute.scala 117:10]
  wire  _GEN_5631; // @[Execute.scala 117:10]
  wire  _GEN_5632; // @[Execute.scala 117:10]
  wire  _GEN_5633; // @[Execute.scala 117:10]
  wire  _T_521; // @[Execute.scala 117:10]
  wire  _T_522; // @[Execute.scala 117:15]
  wire [5:0] _T_524; // @[Execute.scala 117:37]
  wire [5:0] _T_528; // @[Execute.scala 117:60]
  wire  _GEN_5635; // @[Execute.scala 117:10]
  wire  _GEN_5636; // @[Execute.scala 117:10]
  wire  _GEN_5637; // @[Execute.scala 117:10]
  wire  _GEN_5638; // @[Execute.scala 117:10]
  wire  _GEN_5639; // @[Execute.scala 117:10]
  wire  _GEN_5640; // @[Execute.scala 117:10]
  wire  _GEN_5641; // @[Execute.scala 117:10]
  wire  _GEN_5642; // @[Execute.scala 117:10]
  wire  _GEN_5643; // @[Execute.scala 117:10]
  wire  _GEN_5644; // @[Execute.scala 117:10]
  wire  _GEN_5645; // @[Execute.scala 117:10]
  wire  _GEN_5646; // @[Execute.scala 117:10]
  wire  _GEN_5647; // @[Execute.scala 117:10]
  wire  _GEN_5648; // @[Execute.scala 117:10]
  wire  _GEN_5649; // @[Execute.scala 117:10]
  wire  _GEN_5650; // @[Execute.scala 117:10]
  wire  _GEN_5651; // @[Execute.scala 117:10]
  wire  _GEN_5652; // @[Execute.scala 117:10]
  wire  _GEN_5653; // @[Execute.scala 117:10]
  wire  _GEN_5654; // @[Execute.scala 117:10]
  wire  _GEN_5655; // @[Execute.scala 117:10]
  wire  _GEN_5656; // @[Execute.scala 117:10]
  wire  _GEN_5657; // @[Execute.scala 117:10]
  wire  _GEN_5658; // @[Execute.scala 117:10]
  wire  _GEN_5659; // @[Execute.scala 117:10]
  wire  _GEN_5660; // @[Execute.scala 117:10]
  wire  _GEN_5661; // @[Execute.scala 117:10]
  wire  _GEN_5662; // @[Execute.scala 117:10]
  wire  _GEN_5663; // @[Execute.scala 117:10]
  wire  _GEN_5664; // @[Execute.scala 117:10]
  wire  _GEN_5665; // @[Execute.scala 117:10]
  wire  _GEN_5666; // @[Execute.scala 117:10]
  wire  _GEN_5667; // @[Execute.scala 117:10]
  wire  _GEN_5668; // @[Execute.scala 117:10]
  wire  _GEN_5669; // @[Execute.scala 117:10]
  wire  _GEN_5670; // @[Execute.scala 117:10]
  wire  _GEN_5671; // @[Execute.scala 117:10]
  wire  _GEN_5672; // @[Execute.scala 117:10]
  wire  _GEN_5673; // @[Execute.scala 117:10]
  wire  _GEN_5674; // @[Execute.scala 117:10]
  wire  _GEN_5675; // @[Execute.scala 117:10]
  wire  _GEN_5676; // @[Execute.scala 117:10]
  wire  _GEN_5677; // @[Execute.scala 117:10]
  wire  _GEN_5678; // @[Execute.scala 117:10]
  wire  _GEN_5679; // @[Execute.scala 117:10]
  wire  _GEN_5680; // @[Execute.scala 117:10]
  wire  _GEN_5681; // @[Execute.scala 117:10]
  wire  _GEN_5682; // @[Execute.scala 117:10]
  wire  _GEN_5683; // @[Execute.scala 117:10]
  wire  _GEN_5684; // @[Execute.scala 117:10]
  wire  _GEN_5685; // @[Execute.scala 117:10]
  wire  _GEN_5686; // @[Execute.scala 117:10]
  wire  _GEN_5687; // @[Execute.scala 117:10]
  wire  _GEN_5688; // @[Execute.scala 117:10]
  wire  _GEN_5689; // @[Execute.scala 117:10]
  wire  _GEN_5690; // @[Execute.scala 117:10]
  wire  _GEN_5691; // @[Execute.scala 117:10]
  wire  _GEN_5692; // @[Execute.scala 117:10]
  wire  _GEN_5693; // @[Execute.scala 117:10]
  wire  _GEN_5694; // @[Execute.scala 117:10]
  wire  _GEN_5695; // @[Execute.scala 117:10]
  wire  _GEN_5696; // @[Execute.scala 117:10]
  wire  _GEN_5697; // @[Execute.scala 117:10]
  wire  _GEN_5699; // @[Execute.scala 117:10]
  wire  _GEN_5700; // @[Execute.scala 117:10]
  wire  _GEN_5701; // @[Execute.scala 117:10]
  wire  _GEN_5702; // @[Execute.scala 117:10]
  wire  _GEN_5703; // @[Execute.scala 117:10]
  wire  _GEN_5704; // @[Execute.scala 117:10]
  wire  _GEN_5705; // @[Execute.scala 117:10]
  wire  _GEN_5706; // @[Execute.scala 117:10]
  wire  _GEN_5707; // @[Execute.scala 117:10]
  wire  _GEN_5708; // @[Execute.scala 117:10]
  wire  _GEN_5709; // @[Execute.scala 117:10]
  wire  _GEN_5710; // @[Execute.scala 117:10]
  wire  _GEN_5711; // @[Execute.scala 117:10]
  wire  _GEN_5712; // @[Execute.scala 117:10]
  wire  _GEN_5713; // @[Execute.scala 117:10]
  wire  _GEN_5714; // @[Execute.scala 117:10]
  wire  _GEN_5715; // @[Execute.scala 117:10]
  wire  _GEN_5716; // @[Execute.scala 117:10]
  wire  _GEN_5717; // @[Execute.scala 117:10]
  wire  _GEN_5718; // @[Execute.scala 117:10]
  wire  _GEN_5719; // @[Execute.scala 117:10]
  wire  _GEN_5720; // @[Execute.scala 117:10]
  wire  _GEN_5721; // @[Execute.scala 117:10]
  wire  _GEN_5722; // @[Execute.scala 117:10]
  wire  _GEN_5723; // @[Execute.scala 117:10]
  wire  _GEN_5724; // @[Execute.scala 117:10]
  wire  _GEN_5725; // @[Execute.scala 117:10]
  wire  _GEN_5726; // @[Execute.scala 117:10]
  wire  _GEN_5727; // @[Execute.scala 117:10]
  wire  _GEN_5728; // @[Execute.scala 117:10]
  wire  _GEN_5729; // @[Execute.scala 117:10]
  wire  _GEN_5730; // @[Execute.scala 117:10]
  wire  _GEN_5731; // @[Execute.scala 117:10]
  wire  _GEN_5732; // @[Execute.scala 117:10]
  wire  _GEN_5733; // @[Execute.scala 117:10]
  wire  _GEN_5734; // @[Execute.scala 117:10]
  wire  _GEN_5735; // @[Execute.scala 117:10]
  wire  _GEN_5736; // @[Execute.scala 117:10]
  wire  _GEN_5737; // @[Execute.scala 117:10]
  wire  _GEN_5738; // @[Execute.scala 117:10]
  wire  _GEN_5739; // @[Execute.scala 117:10]
  wire  _GEN_5740; // @[Execute.scala 117:10]
  wire  _GEN_5741; // @[Execute.scala 117:10]
  wire  _GEN_5742; // @[Execute.scala 117:10]
  wire  _GEN_5743; // @[Execute.scala 117:10]
  wire  _GEN_5744; // @[Execute.scala 117:10]
  wire  _GEN_5745; // @[Execute.scala 117:10]
  wire  _GEN_5746; // @[Execute.scala 117:10]
  wire  _GEN_5747; // @[Execute.scala 117:10]
  wire  _GEN_5748; // @[Execute.scala 117:10]
  wire  _GEN_5749; // @[Execute.scala 117:10]
  wire  _GEN_5750; // @[Execute.scala 117:10]
  wire  _GEN_5751; // @[Execute.scala 117:10]
  wire  _GEN_5752; // @[Execute.scala 117:10]
  wire  _GEN_5753; // @[Execute.scala 117:10]
  wire  _GEN_5754; // @[Execute.scala 117:10]
  wire  _GEN_5755; // @[Execute.scala 117:10]
  wire  _GEN_5756; // @[Execute.scala 117:10]
  wire  _GEN_5757; // @[Execute.scala 117:10]
  wire  _GEN_5758; // @[Execute.scala 117:10]
  wire  _GEN_5759; // @[Execute.scala 117:10]
  wire  _GEN_5760; // @[Execute.scala 117:10]
  wire  _GEN_5761; // @[Execute.scala 117:10]
  wire  _T_531; // @[Execute.scala 117:10]
  wire  _T_532; // @[Execute.scala 117:15]
  wire [5:0] _T_534; // @[Execute.scala 117:37]
  wire [5:0] _T_538; // @[Execute.scala 117:60]
  wire  _GEN_5763; // @[Execute.scala 117:10]
  wire  _GEN_5764; // @[Execute.scala 117:10]
  wire  _GEN_5765; // @[Execute.scala 117:10]
  wire  _GEN_5766; // @[Execute.scala 117:10]
  wire  _GEN_5767; // @[Execute.scala 117:10]
  wire  _GEN_5768; // @[Execute.scala 117:10]
  wire  _GEN_5769; // @[Execute.scala 117:10]
  wire  _GEN_5770; // @[Execute.scala 117:10]
  wire  _GEN_5771; // @[Execute.scala 117:10]
  wire  _GEN_5772; // @[Execute.scala 117:10]
  wire  _GEN_5773; // @[Execute.scala 117:10]
  wire  _GEN_5774; // @[Execute.scala 117:10]
  wire  _GEN_5775; // @[Execute.scala 117:10]
  wire  _GEN_5776; // @[Execute.scala 117:10]
  wire  _GEN_5777; // @[Execute.scala 117:10]
  wire  _GEN_5778; // @[Execute.scala 117:10]
  wire  _GEN_5779; // @[Execute.scala 117:10]
  wire  _GEN_5780; // @[Execute.scala 117:10]
  wire  _GEN_5781; // @[Execute.scala 117:10]
  wire  _GEN_5782; // @[Execute.scala 117:10]
  wire  _GEN_5783; // @[Execute.scala 117:10]
  wire  _GEN_5784; // @[Execute.scala 117:10]
  wire  _GEN_5785; // @[Execute.scala 117:10]
  wire  _GEN_5786; // @[Execute.scala 117:10]
  wire  _GEN_5787; // @[Execute.scala 117:10]
  wire  _GEN_5788; // @[Execute.scala 117:10]
  wire  _GEN_5789; // @[Execute.scala 117:10]
  wire  _GEN_5790; // @[Execute.scala 117:10]
  wire  _GEN_5791; // @[Execute.scala 117:10]
  wire  _GEN_5792; // @[Execute.scala 117:10]
  wire  _GEN_5793; // @[Execute.scala 117:10]
  wire  _GEN_5794; // @[Execute.scala 117:10]
  wire  _GEN_5795; // @[Execute.scala 117:10]
  wire  _GEN_5796; // @[Execute.scala 117:10]
  wire  _GEN_5797; // @[Execute.scala 117:10]
  wire  _GEN_5798; // @[Execute.scala 117:10]
  wire  _GEN_5799; // @[Execute.scala 117:10]
  wire  _GEN_5800; // @[Execute.scala 117:10]
  wire  _GEN_5801; // @[Execute.scala 117:10]
  wire  _GEN_5802; // @[Execute.scala 117:10]
  wire  _GEN_5803; // @[Execute.scala 117:10]
  wire  _GEN_5804; // @[Execute.scala 117:10]
  wire  _GEN_5805; // @[Execute.scala 117:10]
  wire  _GEN_5806; // @[Execute.scala 117:10]
  wire  _GEN_5807; // @[Execute.scala 117:10]
  wire  _GEN_5808; // @[Execute.scala 117:10]
  wire  _GEN_5809; // @[Execute.scala 117:10]
  wire  _GEN_5810; // @[Execute.scala 117:10]
  wire  _GEN_5811; // @[Execute.scala 117:10]
  wire  _GEN_5812; // @[Execute.scala 117:10]
  wire  _GEN_5813; // @[Execute.scala 117:10]
  wire  _GEN_5814; // @[Execute.scala 117:10]
  wire  _GEN_5815; // @[Execute.scala 117:10]
  wire  _GEN_5816; // @[Execute.scala 117:10]
  wire  _GEN_5817; // @[Execute.scala 117:10]
  wire  _GEN_5818; // @[Execute.scala 117:10]
  wire  _GEN_5819; // @[Execute.scala 117:10]
  wire  _GEN_5820; // @[Execute.scala 117:10]
  wire  _GEN_5821; // @[Execute.scala 117:10]
  wire  _GEN_5822; // @[Execute.scala 117:10]
  wire  _GEN_5823; // @[Execute.scala 117:10]
  wire  _GEN_5824; // @[Execute.scala 117:10]
  wire  _GEN_5825; // @[Execute.scala 117:10]
  wire  _GEN_5827; // @[Execute.scala 117:10]
  wire  _GEN_5828; // @[Execute.scala 117:10]
  wire  _GEN_5829; // @[Execute.scala 117:10]
  wire  _GEN_5830; // @[Execute.scala 117:10]
  wire  _GEN_5831; // @[Execute.scala 117:10]
  wire  _GEN_5832; // @[Execute.scala 117:10]
  wire  _GEN_5833; // @[Execute.scala 117:10]
  wire  _GEN_5834; // @[Execute.scala 117:10]
  wire  _GEN_5835; // @[Execute.scala 117:10]
  wire  _GEN_5836; // @[Execute.scala 117:10]
  wire  _GEN_5837; // @[Execute.scala 117:10]
  wire  _GEN_5838; // @[Execute.scala 117:10]
  wire  _GEN_5839; // @[Execute.scala 117:10]
  wire  _GEN_5840; // @[Execute.scala 117:10]
  wire  _GEN_5841; // @[Execute.scala 117:10]
  wire  _GEN_5842; // @[Execute.scala 117:10]
  wire  _GEN_5843; // @[Execute.scala 117:10]
  wire  _GEN_5844; // @[Execute.scala 117:10]
  wire  _GEN_5845; // @[Execute.scala 117:10]
  wire  _GEN_5846; // @[Execute.scala 117:10]
  wire  _GEN_5847; // @[Execute.scala 117:10]
  wire  _GEN_5848; // @[Execute.scala 117:10]
  wire  _GEN_5849; // @[Execute.scala 117:10]
  wire  _GEN_5850; // @[Execute.scala 117:10]
  wire  _GEN_5851; // @[Execute.scala 117:10]
  wire  _GEN_5852; // @[Execute.scala 117:10]
  wire  _GEN_5853; // @[Execute.scala 117:10]
  wire  _GEN_5854; // @[Execute.scala 117:10]
  wire  _GEN_5855; // @[Execute.scala 117:10]
  wire  _GEN_5856; // @[Execute.scala 117:10]
  wire  _GEN_5857; // @[Execute.scala 117:10]
  wire  _GEN_5858; // @[Execute.scala 117:10]
  wire  _GEN_5859; // @[Execute.scala 117:10]
  wire  _GEN_5860; // @[Execute.scala 117:10]
  wire  _GEN_5861; // @[Execute.scala 117:10]
  wire  _GEN_5862; // @[Execute.scala 117:10]
  wire  _GEN_5863; // @[Execute.scala 117:10]
  wire  _GEN_5864; // @[Execute.scala 117:10]
  wire  _GEN_5865; // @[Execute.scala 117:10]
  wire  _GEN_5866; // @[Execute.scala 117:10]
  wire  _GEN_5867; // @[Execute.scala 117:10]
  wire  _GEN_5868; // @[Execute.scala 117:10]
  wire  _GEN_5869; // @[Execute.scala 117:10]
  wire  _GEN_5870; // @[Execute.scala 117:10]
  wire  _GEN_5871; // @[Execute.scala 117:10]
  wire  _GEN_5872; // @[Execute.scala 117:10]
  wire  _GEN_5873; // @[Execute.scala 117:10]
  wire  _GEN_5874; // @[Execute.scala 117:10]
  wire  _GEN_5875; // @[Execute.scala 117:10]
  wire  _GEN_5876; // @[Execute.scala 117:10]
  wire  _GEN_5877; // @[Execute.scala 117:10]
  wire  _GEN_5878; // @[Execute.scala 117:10]
  wire  _GEN_5879; // @[Execute.scala 117:10]
  wire  _GEN_5880; // @[Execute.scala 117:10]
  wire  _GEN_5881; // @[Execute.scala 117:10]
  wire  _GEN_5882; // @[Execute.scala 117:10]
  wire  _GEN_5883; // @[Execute.scala 117:10]
  wire  _GEN_5884; // @[Execute.scala 117:10]
  wire  _GEN_5885; // @[Execute.scala 117:10]
  wire  _GEN_5886; // @[Execute.scala 117:10]
  wire  _GEN_5887; // @[Execute.scala 117:10]
  wire  _GEN_5888; // @[Execute.scala 117:10]
  wire  _GEN_5889; // @[Execute.scala 117:10]
  wire  _T_541; // @[Execute.scala 117:10]
  wire  _T_542; // @[Execute.scala 117:15]
  wire [5:0] _T_544; // @[Execute.scala 117:37]
  wire [5:0] _T_548; // @[Execute.scala 117:60]
  wire  _GEN_5891; // @[Execute.scala 117:10]
  wire  _GEN_5892; // @[Execute.scala 117:10]
  wire  _GEN_5893; // @[Execute.scala 117:10]
  wire  _GEN_5894; // @[Execute.scala 117:10]
  wire  _GEN_5895; // @[Execute.scala 117:10]
  wire  _GEN_5896; // @[Execute.scala 117:10]
  wire  _GEN_5897; // @[Execute.scala 117:10]
  wire  _GEN_5898; // @[Execute.scala 117:10]
  wire  _GEN_5899; // @[Execute.scala 117:10]
  wire  _GEN_5900; // @[Execute.scala 117:10]
  wire  _GEN_5901; // @[Execute.scala 117:10]
  wire  _GEN_5902; // @[Execute.scala 117:10]
  wire  _GEN_5903; // @[Execute.scala 117:10]
  wire  _GEN_5904; // @[Execute.scala 117:10]
  wire  _GEN_5905; // @[Execute.scala 117:10]
  wire  _GEN_5906; // @[Execute.scala 117:10]
  wire  _GEN_5907; // @[Execute.scala 117:10]
  wire  _GEN_5908; // @[Execute.scala 117:10]
  wire  _GEN_5909; // @[Execute.scala 117:10]
  wire  _GEN_5910; // @[Execute.scala 117:10]
  wire  _GEN_5911; // @[Execute.scala 117:10]
  wire  _GEN_5912; // @[Execute.scala 117:10]
  wire  _GEN_5913; // @[Execute.scala 117:10]
  wire  _GEN_5914; // @[Execute.scala 117:10]
  wire  _GEN_5915; // @[Execute.scala 117:10]
  wire  _GEN_5916; // @[Execute.scala 117:10]
  wire  _GEN_5917; // @[Execute.scala 117:10]
  wire  _GEN_5918; // @[Execute.scala 117:10]
  wire  _GEN_5919; // @[Execute.scala 117:10]
  wire  _GEN_5920; // @[Execute.scala 117:10]
  wire  _GEN_5921; // @[Execute.scala 117:10]
  wire  _GEN_5922; // @[Execute.scala 117:10]
  wire  _GEN_5923; // @[Execute.scala 117:10]
  wire  _GEN_5924; // @[Execute.scala 117:10]
  wire  _GEN_5925; // @[Execute.scala 117:10]
  wire  _GEN_5926; // @[Execute.scala 117:10]
  wire  _GEN_5927; // @[Execute.scala 117:10]
  wire  _GEN_5928; // @[Execute.scala 117:10]
  wire  _GEN_5929; // @[Execute.scala 117:10]
  wire  _GEN_5930; // @[Execute.scala 117:10]
  wire  _GEN_5931; // @[Execute.scala 117:10]
  wire  _GEN_5932; // @[Execute.scala 117:10]
  wire  _GEN_5933; // @[Execute.scala 117:10]
  wire  _GEN_5934; // @[Execute.scala 117:10]
  wire  _GEN_5935; // @[Execute.scala 117:10]
  wire  _GEN_5936; // @[Execute.scala 117:10]
  wire  _GEN_5937; // @[Execute.scala 117:10]
  wire  _GEN_5938; // @[Execute.scala 117:10]
  wire  _GEN_5939; // @[Execute.scala 117:10]
  wire  _GEN_5940; // @[Execute.scala 117:10]
  wire  _GEN_5941; // @[Execute.scala 117:10]
  wire  _GEN_5942; // @[Execute.scala 117:10]
  wire  _GEN_5943; // @[Execute.scala 117:10]
  wire  _GEN_5944; // @[Execute.scala 117:10]
  wire  _GEN_5945; // @[Execute.scala 117:10]
  wire  _GEN_5946; // @[Execute.scala 117:10]
  wire  _GEN_5947; // @[Execute.scala 117:10]
  wire  _GEN_5948; // @[Execute.scala 117:10]
  wire  _GEN_5949; // @[Execute.scala 117:10]
  wire  _GEN_5950; // @[Execute.scala 117:10]
  wire  _GEN_5951; // @[Execute.scala 117:10]
  wire  _GEN_5952; // @[Execute.scala 117:10]
  wire  _GEN_5953; // @[Execute.scala 117:10]
  wire  _GEN_5955; // @[Execute.scala 117:10]
  wire  _GEN_5956; // @[Execute.scala 117:10]
  wire  _GEN_5957; // @[Execute.scala 117:10]
  wire  _GEN_5958; // @[Execute.scala 117:10]
  wire  _GEN_5959; // @[Execute.scala 117:10]
  wire  _GEN_5960; // @[Execute.scala 117:10]
  wire  _GEN_5961; // @[Execute.scala 117:10]
  wire  _GEN_5962; // @[Execute.scala 117:10]
  wire  _GEN_5963; // @[Execute.scala 117:10]
  wire  _GEN_5964; // @[Execute.scala 117:10]
  wire  _GEN_5965; // @[Execute.scala 117:10]
  wire  _GEN_5966; // @[Execute.scala 117:10]
  wire  _GEN_5967; // @[Execute.scala 117:10]
  wire  _GEN_5968; // @[Execute.scala 117:10]
  wire  _GEN_5969; // @[Execute.scala 117:10]
  wire  _GEN_5970; // @[Execute.scala 117:10]
  wire  _GEN_5971; // @[Execute.scala 117:10]
  wire  _GEN_5972; // @[Execute.scala 117:10]
  wire  _GEN_5973; // @[Execute.scala 117:10]
  wire  _GEN_5974; // @[Execute.scala 117:10]
  wire  _GEN_5975; // @[Execute.scala 117:10]
  wire  _GEN_5976; // @[Execute.scala 117:10]
  wire  _GEN_5977; // @[Execute.scala 117:10]
  wire  _GEN_5978; // @[Execute.scala 117:10]
  wire  _GEN_5979; // @[Execute.scala 117:10]
  wire  _GEN_5980; // @[Execute.scala 117:10]
  wire  _GEN_5981; // @[Execute.scala 117:10]
  wire  _GEN_5982; // @[Execute.scala 117:10]
  wire  _GEN_5983; // @[Execute.scala 117:10]
  wire  _GEN_5984; // @[Execute.scala 117:10]
  wire  _GEN_5985; // @[Execute.scala 117:10]
  wire  _GEN_5986; // @[Execute.scala 117:10]
  wire  _GEN_5987; // @[Execute.scala 117:10]
  wire  _GEN_5988; // @[Execute.scala 117:10]
  wire  _GEN_5989; // @[Execute.scala 117:10]
  wire  _GEN_5990; // @[Execute.scala 117:10]
  wire  _GEN_5991; // @[Execute.scala 117:10]
  wire  _GEN_5992; // @[Execute.scala 117:10]
  wire  _GEN_5993; // @[Execute.scala 117:10]
  wire  _GEN_5994; // @[Execute.scala 117:10]
  wire  _GEN_5995; // @[Execute.scala 117:10]
  wire  _GEN_5996; // @[Execute.scala 117:10]
  wire  _GEN_5997; // @[Execute.scala 117:10]
  wire  _GEN_5998; // @[Execute.scala 117:10]
  wire  _GEN_5999; // @[Execute.scala 117:10]
  wire  _GEN_6000; // @[Execute.scala 117:10]
  wire  _GEN_6001; // @[Execute.scala 117:10]
  wire  _GEN_6002; // @[Execute.scala 117:10]
  wire  _GEN_6003; // @[Execute.scala 117:10]
  wire  _GEN_6004; // @[Execute.scala 117:10]
  wire  _GEN_6005; // @[Execute.scala 117:10]
  wire  _GEN_6006; // @[Execute.scala 117:10]
  wire  _GEN_6007; // @[Execute.scala 117:10]
  wire  _GEN_6008; // @[Execute.scala 117:10]
  wire  _GEN_6009; // @[Execute.scala 117:10]
  wire  _GEN_6010; // @[Execute.scala 117:10]
  wire  _GEN_6011; // @[Execute.scala 117:10]
  wire  _GEN_6012; // @[Execute.scala 117:10]
  wire  _GEN_6013; // @[Execute.scala 117:10]
  wire  _GEN_6014; // @[Execute.scala 117:10]
  wire  _GEN_6015; // @[Execute.scala 117:10]
  wire  _GEN_6016; // @[Execute.scala 117:10]
  wire  _GEN_6017; // @[Execute.scala 117:10]
  wire  _T_551; // @[Execute.scala 117:10]
  wire  _T_552; // @[Execute.scala 117:15]
  wire [5:0] _T_554; // @[Execute.scala 117:37]
  wire [5:0] _T_558; // @[Execute.scala 117:60]
  wire  _GEN_6019; // @[Execute.scala 117:10]
  wire  _GEN_6020; // @[Execute.scala 117:10]
  wire  _GEN_6021; // @[Execute.scala 117:10]
  wire  _GEN_6022; // @[Execute.scala 117:10]
  wire  _GEN_6023; // @[Execute.scala 117:10]
  wire  _GEN_6024; // @[Execute.scala 117:10]
  wire  _GEN_6025; // @[Execute.scala 117:10]
  wire  _GEN_6026; // @[Execute.scala 117:10]
  wire  _GEN_6027; // @[Execute.scala 117:10]
  wire  _GEN_6028; // @[Execute.scala 117:10]
  wire  _GEN_6029; // @[Execute.scala 117:10]
  wire  _GEN_6030; // @[Execute.scala 117:10]
  wire  _GEN_6031; // @[Execute.scala 117:10]
  wire  _GEN_6032; // @[Execute.scala 117:10]
  wire  _GEN_6033; // @[Execute.scala 117:10]
  wire  _GEN_6034; // @[Execute.scala 117:10]
  wire  _GEN_6035; // @[Execute.scala 117:10]
  wire  _GEN_6036; // @[Execute.scala 117:10]
  wire  _GEN_6037; // @[Execute.scala 117:10]
  wire  _GEN_6038; // @[Execute.scala 117:10]
  wire  _GEN_6039; // @[Execute.scala 117:10]
  wire  _GEN_6040; // @[Execute.scala 117:10]
  wire  _GEN_6041; // @[Execute.scala 117:10]
  wire  _GEN_6042; // @[Execute.scala 117:10]
  wire  _GEN_6043; // @[Execute.scala 117:10]
  wire  _GEN_6044; // @[Execute.scala 117:10]
  wire  _GEN_6045; // @[Execute.scala 117:10]
  wire  _GEN_6046; // @[Execute.scala 117:10]
  wire  _GEN_6047; // @[Execute.scala 117:10]
  wire  _GEN_6048; // @[Execute.scala 117:10]
  wire  _GEN_6049; // @[Execute.scala 117:10]
  wire  _GEN_6050; // @[Execute.scala 117:10]
  wire  _GEN_6051; // @[Execute.scala 117:10]
  wire  _GEN_6052; // @[Execute.scala 117:10]
  wire  _GEN_6053; // @[Execute.scala 117:10]
  wire  _GEN_6054; // @[Execute.scala 117:10]
  wire  _GEN_6055; // @[Execute.scala 117:10]
  wire  _GEN_6056; // @[Execute.scala 117:10]
  wire  _GEN_6057; // @[Execute.scala 117:10]
  wire  _GEN_6058; // @[Execute.scala 117:10]
  wire  _GEN_6059; // @[Execute.scala 117:10]
  wire  _GEN_6060; // @[Execute.scala 117:10]
  wire  _GEN_6061; // @[Execute.scala 117:10]
  wire  _GEN_6062; // @[Execute.scala 117:10]
  wire  _GEN_6063; // @[Execute.scala 117:10]
  wire  _GEN_6064; // @[Execute.scala 117:10]
  wire  _GEN_6065; // @[Execute.scala 117:10]
  wire  _GEN_6066; // @[Execute.scala 117:10]
  wire  _GEN_6067; // @[Execute.scala 117:10]
  wire  _GEN_6068; // @[Execute.scala 117:10]
  wire  _GEN_6069; // @[Execute.scala 117:10]
  wire  _GEN_6070; // @[Execute.scala 117:10]
  wire  _GEN_6071; // @[Execute.scala 117:10]
  wire  _GEN_6072; // @[Execute.scala 117:10]
  wire  _GEN_6073; // @[Execute.scala 117:10]
  wire  _GEN_6074; // @[Execute.scala 117:10]
  wire  _GEN_6075; // @[Execute.scala 117:10]
  wire  _GEN_6076; // @[Execute.scala 117:10]
  wire  _GEN_6077; // @[Execute.scala 117:10]
  wire  _GEN_6078; // @[Execute.scala 117:10]
  wire  _GEN_6079; // @[Execute.scala 117:10]
  wire  _GEN_6080; // @[Execute.scala 117:10]
  wire  _GEN_6081; // @[Execute.scala 117:10]
  wire  _GEN_6083; // @[Execute.scala 117:10]
  wire  _GEN_6084; // @[Execute.scala 117:10]
  wire  _GEN_6085; // @[Execute.scala 117:10]
  wire  _GEN_6086; // @[Execute.scala 117:10]
  wire  _GEN_6087; // @[Execute.scala 117:10]
  wire  _GEN_6088; // @[Execute.scala 117:10]
  wire  _GEN_6089; // @[Execute.scala 117:10]
  wire  _GEN_6090; // @[Execute.scala 117:10]
  wire  _GEN_6091; // @[Execute.scala 117:10]
  wire  _GEN_6092; // @[Execute.scala 117:10]
  wire  _GEN_6093; // @[Execute.scala 117:10]
  wire  _GEN_6094; // @[Execute.scala 117:10]
  wire  _GEN_6095; // @[Execute.scala 117:10]
  wire  _GEN_6096; // @[Execute.scala 117:10]
  wire  _GEN_6097; // @[Execute.scala 117:10]
  wire  _GEN_6098; // @[Execute.scala 117:10]
  wire  _GEN_6099; // @[Execute.scala 117:10]
  wire  _GEN_6100; // @[Execute.scala 117:10]
  wire  _GEN_6101; // @[Execute.scala 117:10]
  wire  _GEN_6102; // @[Execute.scala 117:10]
  wire  _GEN_6103; // @[Execute.scala 117:10]
  wire  _GEN_6104; // @[Execute.scala 117:10]
  wire  _GEN_6105; // @[Execute.scala 117:10]
  wire  _GEN_6106; // @[Execute.scala 117:10]
  wire  _GEN_6107; // @[Execute.scala 117:10]
  wire  _GEN_6108; // @[Execute.scala 117:10]
  wire  _GEN_6109; // @[Execute.scala 117:10]
  wire  _GEN_6110; // @[Execute.scala 117:10]
  wire  _GEN_6111; // @[Execute.scala 117:10]
  wire  _GEN_6112; // @[Execute.scala 117:10]
  wire  _GEN_6113; // @[Execute.scala 117:10]
  wire  _GEN_6114; // @[Execute.scala 117:10]
  wire  _GEN_6115; // @[Execute.scala 117:10]
  wire  _GEN_6116; // @[Execute.scala 117:10]
  wire  _GEN_6117; // @[Execute.scala 117:10]
  wire  _GEN_6118; // @[Execute.scala 117:10]
  wire  _GEN_6119; // @[Execute.scala 117:10]
  wire  _GEN_6120; // @[Execute.scala 117:10]
  wire  _GEN_6121; // @[Execute.scala 117:10]
  wire  _GEN_6122; // @[Execute.scala 117:10]
  wire  _GEN_6123; // @[Execute.scala 117:10]
  wire  _GEN_6124; // @[Execute.scala 117:10]
  wire  _GEN_6125; // @[Execute.scala 117:10]
  wire  _GEN_6126; // @[Execute.scala 117:10]
  wire  _GEN_6127; // @[Execute.scala 117:10]
  wire  _GEN_6128; // @[Execute.scala 117:10]
  wire  _GEN_6129; // @[Execute.scala 117:10]
  wire  _GEN_6130; // @[Execute.scala 117:10]
  wire  _GEN_6131; // @[Execute.scala 117:10]
  wire  _GEN_6132; // @[Execute.scala 117:10]
  wire  _GEN_6133; // @[Execute.scala 117:10]
  wire  _GEN_6134; // @[Execute.scala 117:10]
  wire  _GEN_6135; // @[Execute.scala 117:10]
  wire  _GEN_6136; // @[Execute.scala 117:10]
  wire  _GEN_6137; // @[Execute.scala 117:10]
  wire  _GEN_6138; // @[Execute.scala 117:10]
  wire  _GEN_6139; // @[Execute.scala 117:10]
  wire  _GEN_6140; // @[Execute.scala 117:10]
  wire  _GEN_6141; // @[Execute.scala 117:10]
  wire  _GEN_6142; // @[Execute.scala 117:10]
  wire  _GEN_6143; // @[Execute.scala 117:10]
  wire  _GEN_6144; // @[Execute.scala 117:10]
  wire  _GEN_6145; // @[Execute.scala 117:10]
  wire  _T_561; // @[Execute.scala 117:10]
  wire  _T_562; // @[Execute.scala 117:15]
  wire [5:0] _T_564; // @[Execute.scala 117:37]
  wire [5:0] _T_568; // @[Execute.scala 117:60]
  wire  _GEN_6147; // @[Execute.scala 117:10]
  wire  _GEN_6148; // @[Execute.scala 117:10]
  wire  _GEN_6149; // @[Execute.scala 117:10]
  wire  _GEN_6150; // @[Execute.scala 117:10]
  wire  _GEN_6151; // @[Execute.scala 117:10]
  wire  _GEN_6152; // @[Execute.scala 117:10]
  wire  _GEN_6153; // @[Execute.scala 117:10]
  wire  _GEN_6154; // @[Execute.scala 117:10]
  wire  _GEN_6155; // @[Execute.scala 117:10]
  wire  _GEN_6156; // @[Execute.scala 117:10]
  wire  _GEN_6157; // @[Execute.scala 117:10]
  wire  _GEN_6158; // @[Execute.scala 117:10]
  wire  _GEN_6159; // @[Execute.scala 117:10]
  wire  _GEN_6160; // @[Execute.scala 117:10]
  wire  _GEN_6161; // @[Execute.scala 117:10]
  wire  _GEN_6162; // @[Execute.scala 117:10]
  wire  _GEN_6163; // @[Execute.scala 117:10]
  wire  _GEN_6164; // @[Execute.scala 117:10]
  wire  _GEN_6165; // @[Execute.scala 117:10]
  wire  _GEN_6166; // @[Execute.scala 117:10]
  wire  _GEN_6167; // @[Execute.scala 117:10]
  wire  _GEN_6168; // @[Execute.scala 117:10]
  wire  _GEN_6169; // @[Execute.scala 117:10]
  wire  _GEN_6170; // @[Execute.scala 117:10]
  wire  _GEN_6171; // @[Execute.scala 117:10]
  wire  _GEN_6172; // @[Execute.scala 117:10]
  wire  _GEN_6173; // @[Execute.scala 117:10]
  wire  _GEN_6174; // @[Execute.scala 117:10]
  wire  _GEN_6175; // @[Execute.scala 117:10]
  wire  _GEN_6176; // @[Execute.scala 117:10]
  wire  _GEN_6177; // @[Execute.scala 117:10]
  wire  _GEN_6178; // @[Execute.scala 117:10]
  wire  _GEN_6179; // @[Execute.scala 117:10]
  wire  _GEN_6180; // @[Execute.scala 117:10]
  wire  _GEN_6181; // @[Execute.scala 117:10]
  wire  _GEN_6182; // @[Execute.scala 117:10]
  wire  _GEN_6183; // @[Execute.scala 117:10]
  wire  _GEN_6184; // @[Execute.scala 117:10]
  wire  _GEN_6185; // @[Execute.scala 117:10]
  wire  _GEN_6186; // @[Execute.scala 117:10]
  wire  _GEN_6187; // @[Execute.scala 117:10]
  wire  _GEN_6188; // @[Execute.scala 117:10]
  wire  _GEN_6189; // @[Execute.scala 117:10]
  wire  _GEN_6190; // @[Execute.scala 117:10]
  wire  _GEN_6191; // @[Execute.scala 117:10]
  wire  _GEN_6192; // @[Execute.scala 117:10]
  wire  _GEN_6193; // @[Execute.scala 117:10]
  wire  _GEN_6194; // @[Execute.scala 117:10]
  wire  _GEN_6195; // @[Execute.scala 117:10]
  wire  _GEN_6196; // @[Execute.scala 117:10]
  wire  _GEN_6197; // @[Execute.scala 117:10]
  wire  _GEN_6198; // @[Execute.scala 117:10]
  wire  _GEN_6199; // @[Execute.scala 117:10]
  wire  _GEN_6200; // @[Execute.scala 117:10]
  wire  _GEN_6201; // @[Execute.scala 117:10]
  wire  _GEN_6202; // @[Execute.scala 117:10]
  wire  _GEN_6203; // @[Execute.scala 117:10]
  wire  _GEN_6204; // @[Execute.scala 117:10]
  wire  _GEN_6205; // @[Execute.scala 117:10]
  wire  _GEN_6206; // @[Execute.scala 117:10]
  wire  _GEN_6207; // @[Execute.scala 117:10]
  wire  _GEN_6208; // @[Execute.scala 117:10]
  wire  _GEN_6209; // @[Execute.scala 117:10]
  wire  _GEN_6211; // @[Execute.scala 117:10]
  wire  _GEN_6212; // @[Execute.scala 117:10]
  wire  _GEN_6213; // @[Execute.scala 117:10]
  wire  _GEN_6214; // @[Execute.scala 117:10]
  wire  _GEN_6215; // @[Execute.scala 117:10]
  wire  _GEN_6216; // @[Execute.scala 117:10]
  wire  _GEN_6217; // @[Execute.scala 117:10]
  wire  _GEN_6218; // @[Execute.scala 117:10]
  wire  _GEN_6219; // @[Execute.scala 117:10]
  wire  _GEN_6220; // @[Execute.scala 117:10]
  wire  _GEN_6221; // @[Execute.scala 117:10]
  wire  _GEN_6222; // @[Execute.scala 117:10]
  wire  _GEN_6223; // @[Execute.scala 117:10]
  wire  _GEN_6224; // @[Execute.scala 117:10]
  wire  _GEN_6225; // @[Execute.scala 117:10]
  wire  _GEN_6226; // @[Execute.scala 117:10]
  wire  _GEN_6227; // @[Execute.scala 117:10]
  wire  _GEN_6228; // @[Execute.scala 117:10]
  wire  _GEN_6229; // @[Execute.scala 117:10]
  wire  _GEN_6230; // @[Execute.scala 117:10]
  wire  _GEN_6231; // @[Execute.scala 117:10]
  wire  _GEN_6232; // @[Execute.scala 117:10]
  wire  _GEN_6233; // @[Execute.scala 117:10]
  wire  _GEN_6234; // @[Execute.scala 117:10]
  wire  _GEN_6235; // @[Execute.scala 117:10]
  wire  _GEN_6236; // @[Execute.scala 117:10]
  wire  _GEN_6237; // @[Execute.scala 117:10]
  wire  _GEN_6238; // @[Execute.scala 117:10]
  wire  _GEN_6239; // @[Execute.scala 117:10]
  wire  _GEN_6240; // @[Execute.scala 117:10]
  wire  _GEN_6241; // @[Execute.scala 117:10]
  wire  _GEN_6242; // @[Execute.scala 117:10]
  wire  _GEN_6243; // @[Execute.scala 117:10]
  wire  _GEN_6244; // @[Execute.scala 117:10]
  wire  _GEN_6245; // @[Execute.scala 117:10]
  wire  _GEN_6246; // @[Execute.scala 117:10]
  wire  _GEN_6247; // @[Execute.scala 117:10]
  wire  _GEN_6248; // @[Execute.scala 117:10]
  wire  _GEN_6249; // @[Execute.scala 117:10]
  wire  _GEN_6250; // @[Execute.scala 117:10]
  wire  _GEN_6251; // @[Execute.scala 117:10]
  wire  _GEN_6252; // @[Execute.scala 117:10]
  wire  _GEN_6253; // @[Execute.scala 117:10]
  wire  _GEN_6254; // @[Execute.scala 117:10]
  wire  _GEN_6255; // @[Execute.scala 117:10]
  wire  _GEN_6256; // @[Execute.scala 117:10]
  wire  _GEN_6257; // @[Execute.scala 117:10]
  wire  _GEN_6258; // @[Execute.scala 117:10]
  wire  _GEN_6259; // @[Execute.scala 117:10]
  wire  _GEN_6260; // @[Execute.scala 117:10]
  wire  _GEN_6261; // @[Execute.scala 117:10]
  wire  _GEN_6262; // @[Execute.scala 117:10]
  wire  _GEN_6263; // @[Execute.scala 117:10]
  wire  _GEN_6264; // @[Execute.scala 117:10]
  wire  _GEN_6265; // @[Execute.scala 117:10]
  wire  _GEN_6266; // @[Execute.scala 117:10]
  wire  _GEN_6267; // @[Execute.scala 117:10]
  wire  _GEN_6268; // @[Execute.scala 117:10]
  wire  _GEN_6269; // @[Execute.scala 117:10]
  wire  _GEN_6270; // @[Execute.scala 117:10]
  wire  _GEN_6271; // @[Execute.scala 117:10]
  wire  _GEN_6272; // @[Execute.scala 117:10]
  wire  _GEN_6273; // @[Execute.scala 117:10]
  wire  _T_571; // @[Execute.scala 117:10]
  wire  _T_572; // @[Execute.scala 117:15]
  wire [5:0] _T_574; // @[Execute.scala 117:37]
  wire [5:0] _T_578; // @[Execute.scala 117:60]
  wire  _GEN_6275; // @[Execute.scala 117:10]
  wire  _GEN_6276; // @[Execute.scala 117:10]
  wire  _GEN_6277; // @[Execute.scala 117:10]
  wire  _GEN_6278; // @[Execute.scala 117:10]
  wire  _GEN_6279; // @[Execute.scala 117:10]
  wire  _GEN_6280; // @[Execute.scala 117:10]
  wire  _GEN_6281; // @[Execute.scala 117:10]
  wire  _GEN_6282; // @[Execute.scala 117:10]
  wire  _GEN_6283; // @[Execute.scala 117:10]
  wire  _GEN_6284; // @[Execute.scala 117:10]
  wire  _GEN_6285; // @[Execute.scala 117:10]
  wire  _GEN_6286; // @[Execute.scala 117:10]
  wire  _GEN_6287; // @[Execute.scala 117:10]
  wire  _GEN_6288; // @[Execute.scala 117:10]
  wire  _GEN_6289; // @[Execute.scala 117:10]
  wire  _GEN_6290; // @[Execute.scala 117:10]
  wire  _GEN_6291; // @[Execute.scala 117:10]
  wire  _GEN_6292; // @[Execute.scala 117:10]
  wire  _GEN_6293; // @[Execute.scala 117:10]
  wire  _GEN_6294; // @[Execute.scala 117:10]
  wire  _GEN_6295; // @[Execute.scala 117:10]
  wire  _GEN_6296; // @[Execute.scala 117:10]
  wire  _GEN_6297; // @[Execute.scala 117:10]
  wire  _GEN_6298; // @[Execute.scala 117:10]
  wire  _GEN_6299; // @[Execute.scala 117:10]
  wire  _GEN_6300; // @[Execute.scala 117:10]
  wire  _GEN_6301; // @[Execute.scala 117:10]
  wire  _GEN_6302; // @[Execute.scala 117:10]
  wire  _GEN_6303; // @[Execute.scala 117:10]
  wire  _GEN_6304; // @[Execute.scala 117:10]
  wire  _GEN_6305; // @[Execute.scala 117:10]
  wire  _GEN_6306; // @[Execute.scala 117:10]
  wire  _GEN_6307; // @[Execute.scala 117:10]
  wire  _GEN_6308; // @[Execute.scala 117:10]
  wire  _GEN_6309; // @[Execute.scala 117:10]
  wire  _GEN_6310; // @[Execute.scala 117:10]
  wire  _GEN_6311; // @[Execute.scala 117:10]
  wire  _GEN_6312; // @[Execute.scala 117:10]
  wire  _GEN_6313; // @[Execute.scala 117:10]
  wire  _GEN_6314; // @[Execute.scala 117:10]
  wire  _GEN_6315; // @[Execute.scala 117:10]
  wire  _GEN_6316; // @[Execute.scala 117:10]
  wire  _GEN_6317; // @[Execute.scala 117:10]
  wire  _GEN_6318; // @[Execute.scala 117:10]
  wire  _GEN_6319; // @[Execute.scala 117:10]
  wire  _GEN_6320; // @[Execute.scala 117:10]
  wire  _GEN_6321; // @[Execute.scala 117:10]
  wire  _GEN_6322; // @[Execute.scala 117:10]
  wire  _GEN_6323; // @[Execute.scala 117:10]
  wire  _GEN_6324; // @[Execute.scala 117:10]
  wire  _GEN_6325; // @[Execute.scala 117:10]
  wire  _GEN_6326; // @[Execute.scala 117:10]
  wire  _GEN_6327; // @[Execute.scala 117:10]
  wire  _GEN_6328; // @[Execute.scala 117:10]
  wire  _GEN_6329; // @[Execute.scala 117:10]
  wire  _GEN_6330; // @[Execute.scala 117:10]
  wire  _GEN_6331; // @[Execute.scala 117:10]
  wire  _GEN_6332; // @[Execute.scala 117:10]
  wire  _GEN_6333; // @[Execute.scala 117:10]
  wire  _GEN_6334; // @[Execute.scala 117:10]
  wire  _GEN_6335; // @[Execute.scala 117:10]
  wire  _GEN_6336; // @[Execute.scala 117:10]
  wire  _GEN_6337; // @[Execute.scala 117:10]
  wire  _GEN_6339; // @[Execute.scala 117:10]
  wire  _GEN_6340; // @[Execute.scala 117:10]
  wire  _GEN_6341; // @[Execute.scala 117:10]
  wire  _GEN_6342; // @[Execute.scala 117:10]
  wire  _GEN_6343; // @[Execute.scala 117:10]
  wire  _GEN_6344; // @[Execute.scala 117:10]
  wire  _GEN_6345; // @[Execute.scala 117:10]
  wire  _GEN_6346; // @[Execute.scala 117:10]
  wire  _GEN_6347; // @[Execute.scala 117:10]
  wire  _GEN_6348; // @[Execute.scala 117:10]
  wire  _GEN_6349; // @[Execute.scala 117:10]
  wire  _GEN_6350; // @[Execute.scala 117:10]
  wire  _GEN_6351; // @[Execute.scala 117:10]
  wire  _GEN_6352; // @[Execute.scala 117:10]
  wire  _GEN_6353; // @[Execute.scala 117:10]
  wire  _GEN_6354; // @[Execute.scala 117:10]
  wire  _GEN_6355; // @[Execute.scala 117:10]
  wire  _GEN_6356; // @[Execute.scala 117:10]
  wire  _GEN_6357; // @[Execute.scala 117:10]
  wire  _GEN_6358; // @[Execute.scala 117:10]
  wire  _GEN_6359; // @[Execute.scala 117:10]
  wire  _GEN_6360; // @[Execute.scala 117:10]
  wire  _GEN_6361; // @[Execute.scala 117:10]
  wire  _GEN_6362; // @[Execute.scala 117:10]
  wire  _GEN_6363; // @[Execute.scala 117:10]
  wire  _GEN_6364; // @[Execute.scala 117:10]
  wire  _GEN_6365; // @[Execute.scala 117:10]
  wire  _GEN_6366; // @[Execute.scala 117:10]
  wire  _GEN_6367; // @[Execute.scala 117:10]
  wire  _GEN_6368; // @[Execute.scala 117:10]
  wire  _GEN_6369; // @[Execute.scala 117:10]
  wire  _GEN_6370; // @[Execute.scala 117:10]
  wire  _GEN_6371; // @[Execute.scala 117:10]
  wire  _GEN_6372; // @[Execute.scala 117:10]
  wire  _GEN_6373; // @[Execute.scala 117:10]
  wire  _GEN_6374; // @[Execute.scala 117:10]
  wire  _GEN_6375; // @[Execute.scala 117:10]
  wire  _GEN_6376; // @[Execute.scala 117:10]
  wire  _GEN_6377; // @[Execute.scala 117:10]
  wire  _GEN_6378; // @[Execute.scala 117:10]
  wire  _GEN_6379; // @[Execute.scala 117:10]
  wire  _GEN_6380; // @[Execute.scala 117:10]
  wire  _GEN_6381; // @[Execute.scala 117:10]
  wire  _GEN_6382; // @[Execute.scala 117:10]
  wire  _GEN_6383; // @[Execute.scala 117:10]
  wire  _GEN_6384; // @[Execute.scala 117:10]
  wire  _GEN_6385; // @[Execute.scala 117:10]
  wire  _GEN_6386; // @[Execute.scala 117:10]
  wire  _GEN_6387; // @[Execute.scala 117:10]
  wire  _GEN_6388; // @[Execute.scala 117:10]
  wire  _GEN_6389; // @[Execute.scala 117:10]
  wire  _GEN_6390; // @[Execute.scala 117:10]
  wire  _GEN_6391; // @[Execute.scala 117:10]
  wire  _GEN_6392; // @[Execute.scala 117:10]
  wire  _GEN_6393; // @[Execute.scala 117:10]
  wire  _GEN_6394; // @[Execute.scala 117:10]
  wire  _GEN_6395; // @[Execute.scala 117:10]
  wire  _GEN_6396; // @[Execute.scala 117:10]
  wire  _GEN_6397; // @[Execute.scala 117:10]
  wire  _GEN_6398; // @[Execute.scala 117:10]
  wire  _GEN_6399; // @[Execute.scala 117:10]
  wire  _GEN_6400; // @[Execute.scala 117:10]
  wire  _GEN_6401; // @[Execute.scala 117:10]
  wire  _T_581; // @[Execute.scala 117:10]
  wire  _T_582; // @[Execute.scala 117:15]
  wire [5:0] _T_584; // @[Execute.scala 117:37]
  wire [5:0] _T_588; // @[Execute.scala 117:60]
  wire  _GEN_6403; // @[Execute.scala 117:10]
  wire  _GEN_6404; // @[Execute.scala 117:10]
  wire  _GEN_6405; // @[Execute.scala 117:10]
  wire  _GEN_6406; // @[Execute.scala 117:10]
  wire  _GEN_6407; // @[Execute.scala 117:10]
  wire  _GEN_6408; // @[Execute.scala 117:10]
  wire  _GEN_6409; // @[Execute.scala 117:10]
  wire  _GEN_6410; // @[Execute.scala 117:10]
  wire  _GEN_6411; // @[Execute.scala 117:10]
  wire  _GEN_6412; // @[Execute.scala 117:10]
  wire  _GEN_6413; // @[Execute.scala 117:10]
  wire  _GEN_6414; // @[Execute.scala 117:10]
  wire  _GEN_6415; // @[Execute.scala 117:10]
  wire  _GEN_6416; // @[Execute.scala 117:10]
  wire  _GEN_6417; // @[Execute.scala 117:10]
  wire  _GEN_6418; // @[Execute.scala 117:10]
  wire  _GEN_6419; // @[Execute.scala 117:10]
  wire  _GEN_6420; // @[Execute.scala 117:10]
  wire  _GEN_6421; // @[Execute.scala 117:10]
  wire  _GEN_6422; // @[Execute.scala 117:10]
  wire  _GEN_6423; // @[Execute.scala 117:10]
  wire  _GEN_6424; // @[Execute.scala 117:10]
  wire  _GEN_6425; // @[Execute.scala 117:10]
  wire  _GEN_6426; // @[Execute.scala 117:10]
  wire  _GEN_6427; // @[Execute.scala 117:10]
  wire  _GEN_6428; // @[Execute.scala 117:10]
  wire  _GEN_6429; // @[Execute.scala 117:10]
  wire  _GEN_6430; // @[Execute.scala 117:10]
  wire  _GEN_6431; // @[Execute.scala 117:10]
  wire  _GEN_6432; // @[Execute.scala 117:10]
  wire  _GEN_6433; // @[Execute.scala 117:10]
  wire  _GEN_6434; // @[Execute.scala 117:10]
  wire  _GEN_6435; // @[Execute.scala 117:10]
  wire  _GEN_6436; // @[Execute.scala 117:10]
  wire  _GEN_6437; // @[Execute.scala 117:10]
  wire  _GEN_6438; // @[Execute.scala 117:10]
  wire  _GEN_6439; // @[Execute.scala 117:10]
  wire  _GEN_6440; // @[Execute.scala 117:10]
  wire  _GEN_6441; // @[Execute.scala 117:10]
  wire  _GEN_6442; // @[Execute.scala 117:10]
  wire  _GEN_6443; // @[Execute.scala 117:10]
  wire  _GEN_6444; // @[Execute.scala 117:10]
  wire  _GEN_6445; // @[Execute.scala 117:10]
  wire  _GEN_6446; // @[Execute.scala 117:10]
  wire  _GEN_6447; // @[Execute.scala 117:10]
  wire  _GEN_6448; // @[Execute.scala 117:10]
  wire  _GEN_6449; // @[Execute.scala 117:10]
  wire  _GEN_6450; // @[Execute.scala 117:10]
  wire  _GEN_6451; // @[Execute.scala 117:10]
  wire  _GEN_6452; // @[Execute.scala 117:10]
  wire  _GEN_6453; // @[Execute.scala 117:10]
  wire  _GEN_6454; // @[Execute.scala 117:10]
  wire  _GEN_6455; // @[Execute.scala 117:10]
  wire  _GEN_6456; // @[Execute.scala 117:10]
  wire  _GEN_6457; // @[Execute.scala 117:10]
  wire  _GEN_6458; // @[Execute.scala 117:10]
  wire  _GEN_6459; // @[Execute.scala 117:10]
  wire  _GEN_6460; // @[Execute.scala 117:10]
  wire  _GEN_6461; // @[Execute.scala 117:10]
  wire  _GEN_6462; // @[Execute.scala 117:10]
  wire  _GEN_6463; // @[Execute.scala 117:10]
  wire  _GEN_6464; // @[Execute.scala 117:10]
  wire  _GEN_6465; // @[Execute.scala 117:10]
  wire  _GEN_6467; // @[Execute.scala 117:10]
  wire  _GEN_6468; // @[Execute.scala 117:10]
  wire  _GEN_6469; // @[Execute.scala 117:10]
  wire  _GEN_6470; // @[Execute.scala 117:10]
  wire  _GEN_6471; // @[Execute.scala 117:10]
  wire  _GEN_6472; // @[Execute.scala 117:10]
  wire  _GEN_6473; // @[Execute.scala 117:10]
  wire  _GEN_6474; // @[Execute.scala 117:10]
  wire  _GEN_6475; // @[Execute.scala 117:10]
  wire  _GEN_6476; // @[Execute.scala 117:10]
  wire  _GEN_6477; // @[Execute.scala 117:10]
  wire  _GEN_6478; // @[Execute.scala 117:10]
  wire  _GEN_6479; // @[Execute.scala 117:10]
  wire  _GEN_6480; // @[Execute.scala 117:10]
  wire  _GEN_6481; // @[Execute.scala 117:10]
  wire  _GEN_6482; // @[Execute.scala 117:10]
  wire  _GEN_6483; // @[Execute.scala 117:10]
  wire  _GEN_6484; // @[Execute.scala 117:10]
  wire  _GEN_6485; // @[Execute.scala 117:10]
  wire  _GEN_6486; // @[Execute.scala 117:10]
  wire  _GEN_6487; // @[Execute.scala 117:10]
  wire  _GEN_6488; // @[Execute.scala 117:10]
  wire  _GEN_6489; // @[Execute.scala 117:10]
  wire  _GEN_6490; // @[Execute.scala 117:10]
  wire  _GEN_6491; // @[Execute.scala 117:10]
  wire  _GEN_6492; // @[Execute.scala 117:10]
  wire  _GEN_6493; // @[Execute.scala 117:10]
  wire  _GEN_6494; // @[Execute.scala 117:10]
  wire  _GEN_6495; // @[Execute.scala 117:10]
  wire  _GEN_6496; // @[Execute.scala 117:10]
  wire  _GEN_6497; // @[Execute.scala 117:10]
  wire  _GEN_6498; // @[Execute.scala 117:10]
  wire  _GEN_6499; // @[Execute.scala 117:10]
  wire  _GEN_6500; // @[Execute.scala 117:10]
  wire  _GEN_6501; // @[Execute.scala 117:10]
  wire  _GEN_6502; // @[Execute.scala 117:10]
  wire  _GEN_6503; // @[Execute.scala 117:10]
  wire  _GEN_6504; // @[Execute.scala 117:10]
  wire  _GEN_6505; // @[Execute.scala 117:10]
  wire  _GEN_6506; // @[Execute.scala 117:10]
  wire  _GEN_6507; // @[Execute.scala 117:10]
  wire  _GEN_6508; // @[Execute.scala 117:10]
  wire  _GEN_6509; // @[Execute.scala 117:10]
  wire  _GEN_6510; // @[Execute.scala 117:10]
  wire  _GEN_6511; // @[Execute.scala 117:10]
  wire  _GEN_6512; // @[Execute.scala 117:10]
  wire  _GEN_6513; // @[Execute.scala 117:10]
  wire  _GEN_6514; // @[Execute.scala 117:10]
  wire  _GEN_6515; // @[Execute.scala 117:10]
  wire  _GEN_6516; // @[Execute.scala 117:10]
  wire  _GEN_6517; // @[Execute.scala 117:10]
  wire  _GEN_6518; // @[Execute.scala 117:10]
  wire  _GEN_6519; // @[Execute.scala 117:10]
  wire  _GEN_6520; // @[Execute.scala 117:10]
  wire  _GEN_6521; // @[Execute.scala 117:10]
  wire  _GEN_6522; // @[Execute.scala 117:10]
  wire  _GEN_6523; // @[Execute.scala 117:10]
  wire  _GEN_6524; // @[Execute.scala 117:10]
  wire  _GEN_6525; // @[Execute.scala 117:10]
  wire  _GEN_6526; // @[Execute.scala 117:10]
  wire  _GEN_6527; // @[Execute.scala 117:10]
  wire  _GEN_6528; // @[Execute.scala 117:10]
  wire  _GEN_6529; // @[Execute.scala 117:10]
  wire  _T_591; // @[Execute.scala 117:10]
  wire  _T_592; // @[Execute.scala 117:15]
  wire [5:0] _T_594; // @[Execute.scala 117:37]
  wire [5:0] _T_598; // @[Execute.scala 117:60]
  wire  _GEN_6531; // @[Execute.scala 117:10]
  wire  _GEN_6532; // @[Execute.scala 117:10]
  wire  _GEN_6533; // @[Execute.scala 117:10]
  wire  _GEN_6534; // @[Execute.scala 117:10]
  wire  _GEN_6535; // @[Execute.scala 117:10]
  wire  _GEN_6536; // @[Execute.scala 117:10]
  wire  _GEN_6537; // @[Execute.scala 117:10]
  wire  _GEN_6538; // @[Execute.scala 117:10]
  wire  _GEN_6539; // @[Execute.scala 117:10]
  wire  _GEN_6540; // @[Execute.scala 117:10]
  wire  _GEN_6541; // @[Execute.scala 117:10]
  wire  _GEN_6542; // @[Execute.scala 117:10]
  wire  _GEN_6543; // @[Execute.scala 117:10]
  wire  _GEN_6544; // @[Execute.scala 117:10]
  wire  _GEN_6545; // @[Execute.scala 117:10]
  wire  _GEN_6546; // @[Execute.scala 117:10]
  wire  _GEN_6547; // @[Execute.scala 117:10]
  wire  _GEN_6548; // @[Execute.scala 117:10]
  wire  _GEN_6549; // @[Execute.scala 117:10]
  wire  _GEN_6550; // @[Execute.scala 117:10]
  wire  _GEN_6551; // @[Execute.scala 117:10]
  wire  _GEN_6552; // @[Execute.scala 117:10]
  wire  _GEN_6553; // @[Execute.scala 117:10]
  wire  _GEN_6554; // @[Execute.scala 117:10]
  wire  _GEN_6555; // @[Execute.scala 117:10]
  wire  _GEN_6556; // @[Execute.scala 117:10]
  wire  _GEN_6557; // @[Execute.scala 117:10]
  wire  _GEN_6558; // @[Execute.scala 117:10]
  wire  _GEN_6559; // @[Execute.scala 117:10]
  wire  _GEN_6560; // @[Execute.scala 117:10]
  wire  _GEN_6561; // @[Execute.scala 117:10]
  wire  _GEN_6562; // @[Execute.scala 117:10]
  wire  _GEN_6563; // @[Execute.scala 117:10]
  wire  _GEN_6564; // @[Execute.scala 117:10]
  wire  _GEN_6565; // @[Execute.scala 117:10]
  wire  _GEN_6566; // @[Execute.scala 117:10]
  wire  _GEN_6567; // @[Execute.scala 117:10]
  wire  _GEN_6568; // @[Execute.scala 117:10]
  wire  _GEN_6569; // @[Execute.scala 117:10]
  wire  _GEN_6570; // @[Execute.scala 117:10]
  wire  _GEN_6571; // @[Execute.scala 117:10]
  wire  _GEN_6572; // @[Execute.scala 117:10]
  wire  _GEN_6573; // @[Execute.scala 117:10]
  wire  _GEN_6574; // @[Execute.scala 117:10]
  wire  _GEN_6575; // @[Execute.scala 117:10]
  wire  _GEN_6576; // @[Execute.scala 117:10]
  wire  _GEN_6577; // @[Execute.scala 117:10]
  wire  _GEN_6578; // @[Execute.scala 117:10]
  wire  _GEN_6579; // @[Execute.scala 117:10]
  wire  _GEN_6580; // @[Execute.scala 117:10]
  wire  _GEN_6581; // @[Execute.scala 117:10]
  wire  _GEN_6582; // @[Execute.scala 117:10]
  wire  _GEN_6583; // @[Execute.scala 117:10]
  wire  _GEN_6584; // @[Execute.scala 117:10]
  wire  _GEN_6585; // @[Execute.scala 117:10]
  wire  _GEN_6586; // @[Execute.scala 117:10]
  wire  _GEN_6587; // @[Execute.scala 117:10]
  wire  _GEN_6588; // @[Execute.scala 117:10]
  wire  _GEN_6589; // @[Execute.scala 117:10]
  wire  _GEN_6590; // @[Execute.scala 117:10]
  wire  _GEN_6591; // @[Execute.scala 117:10]
  wire  _GEN_6592; // @[Execute.scala 117:10]
  wire  _GEN_6593; // @[Execute.scala 117:10]
  wire  _GEN_6595; // @[Execute.scala 117:10]
  wire  _GEN_6596; // @[Execute.scala 117:10]
  wire  _GEN_6597; // @[Execute.scala 117:10]
  wire  _GEN_6598; // @[Execute.scala 117:10]
  wire  _GEN_6599; // @[Execute.scala 117:10]
  wire  _GEN_6600; // @[Execute.scala 117:10]
  wire  _GEN_6601; // @[Execute.scala 117:10]
  wire  _GEN_6602; // @[Execute.scala 117:10]
  wire  _GEN_6603; // @[Execute.scala 117:10]
  wire  _GEN_6604; // @[Execute.scala 117:10]
  wire  _GEN_6605; // @[Execute.scala 117:10]
  wire  _GEN_6606; // @[Execute.scala 117:10]
  wire  _GEN_6607; // @[Execute.scala 117:10]
  wire  _GEN_6608; // @[Execute.scala 117:10]
  wire  _GEN_6609; // @[Execute.scala 117:10]
  wire  _GEN_6610; // @[Execute.scala 117:10]
  wire  _GEN_6611; // @[Execute.scala 117:10]
  wire  _GEN_6612; // @[Execute.scala 117:10]
  wire  _GEN_6613; // @[Execute.scala 117:10]
  wire  _GEN_6614; // @[Execute.scala 117:10]
  wire  _GEN_6615; // @[Execute.scala 117:10]
  wire  _GEN_6616; // @[Execute.scala 117:10]
  wire  _GEN_6617; // @[Execute.scala 117:10]
  wire  _GEN_6618; // @[Execute.scala 117:10]
  wire  _GEN_6619; // @[Execute.scala 117:10]
  wire  _GEN_6620; // @[Execute.scala 117:10]
  wire  _GEN_6621; // @[Execute.scala 117:10]
  wire  _GEN_6622; // @[Execute.scala 117:10]
  wire  _GEN_6623; // @[Execute.scala 117:10]
  wire  _GEN_6624; // @[Execute.scala 117:10]
  wire  _GEN_6625; // @[Execute.scala 117:10]
  wire  _GEN_6626; // @[Execute.scala 117:10]
  wire  _GEN_6627; // @[Execute.scala 117:10]
  wire  _GEN_6628; // @[Execute.scala 117:10]
  wire  _GEN_6629; // @[Execute.scala 117:10]
  wire  _GEN_6630; // @[Execute.scala 117:10]
  wire  _GEN_6631; // @[Execute.scala 117:10]
  wire  _GEN_6632; // @[Execute.scala 117:10]
  wire  _GEN_6633; // @[Execute.scala 117:10]
  wire  _GEN_6634; // @[Execute.scala 117:10]
  wire  _GEN_6635; // @[Execute.scala 117:10]
  wire  _GEN_6636; // @[Execute.scala 117:10]
  wire  _GEN_6637; // @[Execute.scala 117:10]
  wire  _GEN_6638; // @[Execute.scala 117:10]
  wire  _GEN_6639; // @[Execute.scala 117:10]
  wire  _GEN_6640; // @[Execute.scala 117:10]
  wire  _GEN_6641; // @[Execute.scala 117:10]
  wire  _GEN_6642; // @[Execute.scala 117:10]
  wire  _GEN_6643; // @[Execute.scala 117:10]
  wire  _GEN_6644; // @[Execute.scala 117:10]
  wire  _GEN_6645; // @[Execute.scala 117:10]
  wire  _GEN_6646; // @[Execute.scala 117:10]
  wire  _GEN_6647; // @[Execute.scala 117:10]
  wire  _GEN_6648; // @[Execute.scala 117:10]
  wire  _GEN_6649; // @[Execute.scala 117:10]
  wire  _GEN_6650; // @[Execute.scala 117:10]
  wire  _GEN_6651; // @[Execute.scala 117:10]
  wire  _GEN_6652; // @[Execute.scala 117:10]
  wire  _GEN_6653; // @[Execute.scala 117:10]
  wire  _GEN_6654; // @[Execute.scala 117:10]
  wire  _GEN_6655; // @[Execute.scala 117:10]
  wire  _GEN_6656; // @[Execute.scala 117:10]
  wire  _GEN_6657; // @[Execute.scala 117:10]
  wire  _T_601; // @[Execute.scala 117:10]
  wire  _T_602; // @[Execute.scala 117:15]
  wire [5:0] _T_604; // @[Execute.scala 117:37]
  wire [5:0] _T_608; // @[Execute.scala 117:60]
  wire  _GEN_6659; // @[Execute.scala 117:10]
  wire  _GEN_6660; // @[Execute.scala 117:10]
  wire  _GEN_6661; // @[Execute.scala 117:10]
  wire  _GEN_6662; // @[Execute.scala 117:10]
  wire  _GEN_6663; // @[Execute.scala 117:10]
  wire  _GEN_6664; // @[Execute.scala 117:10]
  wire  _GEN_6665; // @[Execute.scala 117:10]
  wire  _GEN_6666; // @[Execute.scala 117:10]
  wire  _GEN_6667; // @[Execute.scala 117:10]
  wire  _GEN_6668; // @[Execute.scala 117:10]
  wire  _GEN_6669; // @[Execute.scala 117:10]
  wire  _GEN_6670; // @[Execute.scala 117:10]
  wire  _GEN_6671; // @[Execute.scala 117:10]
  wire  _GEN_6672; // @[Execute.scala 117:10]
  wire  _GEN_6673; // @[Execute.scala 117:10]
  wire  _GEN_6674; // @[Execute.scala 117:10]
  wire  _GEN_6675; // @[Execute.scala 117:10]
  wire  _GEN_6676; // @[Execute.scala 117:10]
  wire  _GEN_6677; // @[Execute.scala 117:10]
  wire  _GEN_6678; // @[Execute.scala 117:10]
  wire  _GEN_6679; // @[Execute.scala 117:10]
  wire  _GEN_6680; // @[Execute.scala 117:10]
  wire  _GEN_6681; // @[Execute.scala 117:10]
  wire  _GEN_6682; // @[Execute.scala 117:10]
  wire  _GEN_6683; // @[Execute.scala 117:10]
  wire  _GEN_6684; // @[Execute.scala 117:10]
  wire  _GEN_6685; // @[Execute.scala 117:10]
  wire  _GEN_6686; // @[Execute.scala 117:10]
  wire  _GEN_6687; // @[Execute.scala 117:10]
  wire  _GEN_6688; // @[Execute.scala 117:10]
  wire  _GEN_6689; // @[Execute.scala 117:10]
  wire  _GEN_6690; // @[Execute.scala 117:10]
  wire  _GEN_6691; // @[Execute.scala 117:10]
  wire  _GEN_6692; // @[Execute.scala 117:10]
  wire  _GEN_6693; // @[Execute.scala 117:10]
  wire  _GEN_6694; // @[Execute.scala 117:10]
  wire  _GEN_6695; // @[Execute.scala 117:10]
  wire  _GEN_6696; // @[Execute.scala 117:10]
  wire  _GEN_6697; // @[Execute.scala 117:10]
  wire  _GEN_6698; // @[Execute.scala 117:10]
  wire  _GEN_6699; // @[Execute.scala 117:10]
  wire  _GEN_6700; // @[Execute.scala 117:10]
  wire  _GEN_6701; // @[Execute.scala 117:10]
  wire  _GEN_6702; // @[Execute.scala 117:10]
  wire  _GEN_6703; // @[Execute.scala 117:10]
  wire  _GEN_6704; // @[Execute.scala 117:10]
  wire  _GEN_6705; // @[Execute.scala 117:10]
  wire  _GEN_6706; // @[Execute.scala 117:10]
  wire  _GEN_6707; // @[Execute.scala 117:10]
  wire  _GEN_6708; // @[Execute.scala 117:10]
  wire  _GEN_6709; // @[Execute.scala 117:10]
  wire  _GEN_6710; // @[Execute.scala 117:10]
  wire  _GEN_6711; // @[Execute.scala 117:10]
  wire  _GEN_6712; // @[Execute.scala 117:10]
  wire  _GEN_6713; // @[Execute.scala 117:10]
  wire  _GEN_6714; // @[Execute.scala 117:10]
  wire  _GEN_6715; // @[Execute.scala 117:10]
  wire  _GEN_6716; // @[Execute.scala 117:10]
  wire  _GEN_6717; // @[Execute.scala 117:10]
  wire  _GEN_6718; // @[Execute.scala 117:10]
  wire  _GEN_6719; // @[Execute.scala 117:10]
  wire  _GEN_6720; // @[Execute.scala 117:10]
  wire  _GEN_6721; // @[Execute.scala 117:10]
  wire  _GEN_6723; // @[Execute.scala 117:10]
  wire  _GEN_6724; // @[Execute.scala 117:10]
  wire  _GEN_6725; // @[Execute.scala 117:10]
  wire  _GEN_6726; // @[Execute.scala 117:10]
  wire  _GEN_6727; // @[Execute.scala 117:10]
  wire  _GEN_6728; // @[Execute.scala 117:10]
  wire  _GEN_6729; // @[Execute.scala 117:10]
  wire  _GEN_6730; // @[Execute.scala 117:10]
  wire  _GEN_6731; // @[Execute.scala 117:10]
  wire  _GEN_6732; // @[Execute.scala 117:10]
  wire  _GEN_6733; // @[Execute.scala 117:10]
  wire  _GEN_6734; // @[Execute.scala 117:10]
  wire  _GEN_6735; // @[Execute.scala 117:10]
  wire  _GEN_6736; // @[Execute.scala 117:10]
  wire  _GEN_6737; // @[Execute.scala 117:10]
  wire  _GEN_6738; // @[Execute.scala 117:10]
  wire  _GEN_6739; // @[Execute.scala 117:10]
  wire  _GEN_6740; // @[Execute.scala 117:10]
  wire  _GEN_6741; // @[Execute.scala 117:10]
  wire  _GEN_6742; // @[Execute.scala 117:10]
  wire  _GEN_6743; // @[Execute.scala 117:10]
  wire  _GEN_6744; // @[Execute.scala 117:10]
  wire  _GEN_6745; // @[Execute.scala 117:10]
  wire  _GEN_6746; // @[Execute.scala 117:10]
  wire  _GEN_6747; // @[Execute.scala 117:10]
  wire  _GEN_6748; // @[Execute.scala 117:10]
  wire  _GEN_6749; // @[Execute.scala 117:10]
  wire  _GEN_6750; // @[Execute.scala 117:10]
  wire  _GEN_6751; // @[Execute.scala 117:10]
  wire  _GEN_6752; // @[Execute.scala 117:10]
  wire  _GEN_6753; // @[Execute.scala 117:10]
  wire  _GEN_6754; // @[Execute.scala 117:10]
  wire  _GEN_6755; // @[Execute.scala 117:10]
  wire  _GEN_6756; // @[Execute.scala 117:10]
  wire  _GEN_6757; // @[Execute.scala 117:10]
  wire  _GEN_6758; // @[Execute.scala 117:10]
  wire  _GEN_6759; // @[Execute.scala 117:10]
  wire  _GEN_6760; // @[Execute.scala 117:10]
  wire  _GEN_6761; // @[Execute.scala 117:10]
  wire  _GEN_6762; // @[Execute.scala 117:10]
  wire  _GEN_6763; // @[Execute.scala 117:10]
  wire  _GEN_6764; // @[Execute.scala 117:10]
  wire  _GEN_6765; // @[Execute.scala 117:10]
  wire  _GEN_6766; // @[Execute.scala 117:10]
  wire  _GEN_6767; // @[Execute.scala 117:10]
  wire  _GEN_6768; // @[Execute.scala 117:10]
  wire  _GEN_6769; // @[Execute.scala 117:10]
  wire  _GEN_6770; // @[Execute.scala 117:10]
  wire  _GEN_6771; // @[Execute.scala 117:10]
  wire  _GEN_6772; // @[Execute.scala 117:10]
  wire  _GEN_6773; // @[Execute.scala 117:10]
  wire  _GEN_6774; // @[Execute.scala 117:10]
  wire  _GEN_6775; // @[Execute.scala 117:10]
  wire  _GEN_6776; // @[Execute.scala 117:10]
  wire  _GEN_6777; // @[Execute.scala 117:10]
  wire  _GEN_6778; // @[Execute.scala 117:10]
  wire  _GEN_6779; // @[Execute.scala 117:10]
  wire  _GEN_6780; // @[Execute.scala 117:10]
  wire  _GEN_6781; // @[Execute.scala 117:10]
  wire  _GEN_6782; // @[Execute.scala 117:10]
  wire  _GEN_6783; // @[Execute.scala 117:10]
  wire  _GEN_6784; // @[Execute.scala 117:10]
  wire  _GEN_6785; // @[Execute.scala 117:10]
  wire  _T_611; // @[Execute.scala 117:10]
  wire  _T_612; // @[Execute.scala 117:15]
  wire [5:0] _T_614; // @[Execute.scala 117:37]
  wire [5:0] _T_618; // @[Execute.scala 117:60]
  wire  _GEN_6787; // @[Execute.scala 117:10]
  wire  _GEN_6788; // @[Execute.scala 117:10]
  wire  _GEN_6789; // @[Execute.scala 117:10]
  wire  _GEN_6790; // @[Execute.scala 117:10]
  wire  _GEN_6791; // @[Execute.scala 117:10]
  wire  _GEN_6792; // @[Execute.scala 117:10]
  wire  _GEN_6793; // @[Execute.scala 117:10]
  wire  _GEN_6794; // @[Execute.scala 117:10]
  wire  _GEN_6795; // @[Execute.scala 117:10]
  wire  _GEN_6796; // @[Execute.scala 117:10]
  wire  _GEN_6797; // @[Execute.scala 117:10]
  wire  _GEN_6798; // @[Execute.scala 117:10]
  wire  _GEN_6799; // @[Execute.scala 117:10]
  wire  _GEN_6800; // @[Execute.scala 117:10]
  wire  _GEN_6801; // @[Execute.scala 117:10]
  wire  _GEN_6802; // @[Execute.scala 117:10]
  wire  _GEN_6803; // @[Execute.scala 117:10]
  wire  _GEN_6804; // @[Execute.scala 117:10]
  wire  _GEN_6805; // @[Execute.scala 117:10]
  wire  _GEN_6806; // @[Execute.scala 117:10]
  wire  _GEN_6807; // @[Execute.scala 117:10]
  wire  _GEN_6808; // @[Execute.scala 117:10]
  wire  _GEN_6809; // @[Execute.scala 117:10]
  wire  _GEN_6810; // @[Execute.scala 117:10]
  wire  _GEN_6811; // @[Execute.scala 117:10]
  wire  _GEN_6812; // @[Execute.scala 117:10]
  wire  _GEN_6813; // @[Execute.scala 117:10]
  wire  _GEN_6814; // @[Execute.scala 117:10]
  wire  _GEN_6815; // @[Execute.scala 117:10]
  wire  _GEN_6816; // @[Execute.scala 117:10]
  wire  _GEN_6817; // @[Execute.scala 117:10]
  wire  _GEN_6818; // @[Execute.scala 117:10]
  wire  _GEN_6819; // @[Execute.scala 117:10]
  wire  _GEN_6820; // @[Execute.scala 117:10]
  wire  _GEN_6821; // @[Execute.scala 117:10]
  wire  _GEN_6822; // @[Execute.scala 117:10]
  wire  _GEN_6823; // @[Execute.scala 117:10]
  wire  _GEN_6824; // @[Execute.scala 117:10]
  wire  _GEN_6825; // @[Execute.scala 117:10]
  wire  _GEN_6826; // @[Execute.scala 117:10]
  wire  _GEN_6827; // @[Execute.scala 117:10]
  wire  _GEN_6828; // @[Execute.scala 117:10]
  wire  _GEN_6829; // @[Execute.scala 117:10]
  wire  _GEN_6830; // @[Execute.scala 117:10]
  wire  _GEN_6831; // @[Execute.scala 117:10]
  wire  _GEN_6832; // @[Execute.scala 117:10]
  wire  _GEN_6833; // @[Execute.scala 117:10]
  wire  _GEN_6834; // @[Execute.scala 117:10]
  wire  _GEN_6835; // @[Execute.scala 117:10]
  wire  _GEN_6836; // @[Execute.scala 117:10]
  wire  _GEN_6837; // @[Execute.scala 117:10]
  wire  _GEN_6838; // @[Execute.scala 117:10]
  wire  _GEN_6839; // @[Execute.scala 117:10]
  wire  _GEN_6840; // @[Execute.scala 117:10]
  wire  _GEN_6841; // @[Execute.scala 117:10]
  wire  _GEN_6842; // @[Execute.scala 117:10]
  wire  _GEN_6843; // @[Execute.scala 117:10]
  wire  _GEN_6844; // @[Execute.scala 117:10]
  wire  _GEN_6845; // @[Execute.scala 117:10]
  wire  _GEN_6846; // @[Execute.scala 117:10]
  wire  _GEN_6847; // @[Execute.scala 117:10]
  wire  _GEN_6848; // @[Execute.scala 117:10]
  wire  _GEN_6849; // @[Execute.scala 117:10]
  wire  _GEN_6851; // @[Execute.scala 117:10]
  wire  _GEN_6852; // @[Execute.scala 117:10]
  wire  _GEN_6853; // @[Execute.scala 117:10]
  wire  _GEN_6854; // @[Execute.scala 117:10]
  wire  _GEN_6855; // @[Execute.scala 117:10]
  wire  _GEN_6856; // @[Execute.scala 117:10]
  wire  _GEN_6857; // @[Execute.scala 117:10]
  wire  _GEN_6858; // @[Execute.scala 117:10]
  wire  _GEN_6859; // @[Execute.scala 117:10]
  wire  _GEN_6860; // @[Execute.scala 117:10]
  wire  _GEN_6861; // @[Execute.scala 117:10]
  wire  _GEN_6862; // @[Execute.scala 117:10]
  wire  _GEN_6863; // @[Execute.scala 117:10]
  wire  _GEN_6864; // @[Execute.scala 117:10]
  wire  _GEN_6865; // @[Execute.scala 117:10]
  wire  _GEN_6866; // @[Execute.scala 117:10]
  wire  _GEN_6867; // @[Execute.scala 117:10]
  wire  _GEN_6868; // @[Execute.scala 117:10]
  wire  _GEN_6869; // @[Execute.scala 117:10]
  wire  _GEN_6870; // @[Execute.scala 117:10]
  wire  _GEN_6871; // @[Execute.scala 117:10]
  wire  _GEN_6872; // @[Execute.scala 117:10]
  wire  _GEN_6873; // @[Execute.scala 117:10]
  wire  _GEN_6874; // @[Execute.scala 117:10]
  wire  _GEN_6875; // @[Execute.scala 117:10]
  wire  _GEN_6876; // @[Execute.scala 117:10]
  wire  _GEN_6877; // @[Execute.scala 117:10]
  wire  _GEN_6878; // @[Execute.scala 117:10]
  wire  _GEN_6879; // @[Execute.scala 117:10]
  wire  _GEN_6880; // @[Execute.scala 117:10]
  wire  _GEN_6881; // @[Execute.scala 117:10]
  wire  _GEN_6882; // @[Execute.scala 117:10]
  wire  _GEN_6883; // @[Execute.scala 117:10]
  wire  _GEN_6884; // @[Execute.scala 117:10]
  wire  _GEN_6885; // @[Execute.scala 117:10]
  wire  _GEN_6886; // @[Execute.scala 117:10]
  wire  _GEN_6887; // @[Execute.scala 117:10]
  wire  _GEN_6888; // @[Execute.scala 117:10]
  wire  _GEN_6889; // @[Execute.scala 117:10]
  wire  _GEN_6890; // @[Execute.scala 117:10]
  wire  _GEN_6891; // @[Execute.scala 117:10]
  wire  _GEN_6892; // @[Execute.scala 117:10]
  wire  _GEN_6893; // @[Execute.scala 117:10]
  wire  _GEN_6894; // @[Execute.scala 117:10]
  wire  _GEN_6895; // @[Execute.scala 117:10]
  wire  _GEN_6896; // @[Execute.scala 117:10]
  wire  _GEN_6897; // @[Execute.scala 117:10]
  wire  _GEN_6898; // @[Execute.scala 117:10]
  wire  _GEN_6899; // @[Execute.scala 117:10]
  wire  _GEN_6900; // @[Execute.scala 117:10]
  wire  _GEN_6901; // @[Execute.scala 117:10]
  wire  _GEN_6902; // @[Execute.scala 117:10]
  wire  _GEN_6903; // @[Execute.scala 117:10]
  wire  _GEN_6904; // @[Execute.scala 117:10]
  wire  _GEN_6905; // @[Execute.scala 117:10]
  wire  _GEN_6906; // @[Execute.scala 117:10]
  wire  _GEN_6907; // @[Execute.scala 117:10]
  wire  _GEN_6908; // @[Execute.scala 117:10]
  wire  _GEN_6909; // @[Execute.scala 117:10]
  wire  _GEN_6910; // @[Execute.scala 117:10]
  wire  _GEN_6911; // @[Execute.scala 117:10]
  wire  _GEN_6912; // @[Execute.scala 117:10]
  wire  _GEN_6913; // @[Execute.scala 117:10]
  wire  _T_621; // @[Execute.scala 117:10]
  wire  _T_622; // @[Execute.scala 117:15]
  wire [5:0] _T_624; // @[Execute.scala 117:37]
  wire [5:0] _T_628; // @[Execute.scala 117:60]
  wire  _GEN_6915; // @[Execute.scala 117:10]
  wire  _GEN_6916; // @[Execute.scala 117:10]
  wire  _GEN_6917; // @[Execute.scala 117:10]
  wire  _GEN_6918; // @[Execute.scala 117:10]
  wire  _GEN_6919; // @[Execute.scala 117:10]
  wire  _GEN_6920; // @[Execute.scala 117:10]
  wire  _GEN_6921; // @[Execute.scala 117:10]
  wire  _GEN_6922; // @[Execute.scala 117:10]
  wire  _GEN_6923; // @[Execute.scala 117:10]
  wire  _GEN_6924; // @[Execute.scala 117:10]
  wire  _GEN_6925; // @[Execute.scala 117:10]
  wire  _GEN_6926; // @[Execute.scala 117:10]
  wire  _GEN_6927; // @[Execute.scala 117:10]
  wire  _GEN_6928; // @[Execute.scala 117:10]
  wire  _GEN_6929; // @[Execute.scala 117:10]
  wire  _GEN_6930; // @[Execute.scala 117:10]
  wire  _GEN_6931; // @[Execute.scala 117:10]
  wire  _GEN_6932; // @[Execute.scala 117:10]
  wire  _GEN_6933; // @[Execute.scala 117:10]
  wire  _GEN_6934; // @[Execute.scala 117:10]
  wire  _GEN_6935; // @[Execute.scala 117:10]
  wire  _GEN_6936; // @[Execute.scala 117:10]
  wire  _GEN_6937; // @[Execute.scala 117:10]
  wire  _GEN_6938; // @[Execute.scala 117:10]
  wire  _GEN_6939; // @[Execute.scala 117:10]
  wire  _GEN_6940; // @[Execute.scala 117:10]
  wire  _GEN_6941; // @[Execute.scala 117:10]
  wire  _GEN_6942; // @[Execute.scala 117:10]
  wire  _GEN_6943; // @[Execute.scala 117:10]
  wire  _GEN_6944; // @[Execute.scala 117:10]
  wire  _GEN_6945; // @[Execute.scala 117:10]
  wire  _GEN_6946; // @[Execute.scala 117:10]
  wire  _GEN_6947; // @[Execute.scala 117:10]
  wire  _GEN_6948; // @[Execute.scala 117:10]
  wire  _GEN_6949; // @[Execute.scala 117:10]
  wire  _GEN_6950; // @[Execute.scala 117:10]
  wire  _GEN_6951; // @[Execute.scala 117:10]
  wire  _GEN_6952; // @[Execute.scala 117:10]
  wire  _GEN_6953; // @[Execute.scala 117:10]
  wire  _GEN_6954; // @[Execute.scala 117:10]
  wire  _GEN_6955; // @[Execute.scala 117:10]
  wire  _GEN_6956; // @[Execute.scala 117:10]
  wire  _GEN_6957; // @[Execute.scala 117:10]
  wire  _GEN_6958; // @[Execute.scala 117:10]
  wire  _GEN_6959; // @[Execute.scala 117:10]
  wire  _GEN_6960; // @[Execute.scala 117:10]
  wire  _GEN_6961; // @[Execute.scala 117:10]
  wire  _GEN_6962; // @[Execute.scala 117:10]
  wire  _GEN_6963; // @[Execute.scala 117:10]
  wire  _GEN_6964; // @[Execute.scala 117:10]
  wire  _GEN_6965; // @[Execute.scala 117:10]
  wire  _GEN_6966; // @[Execute.scala 117:10]
  wire  _GEN_6967; // @[Execute.scala 117:10]
  wire  _GEN_6968; // @[Execute.scala 117:10]
  wire  _GEN_6969; // @[Execute.scala 117:10]
  wire  _GEN_6970; // @[Execute.scala 117:10]
  wire  _GEN_6971; // @[Execute.scala 117:10]
  wire  _GEN_6972; // @[Execute.scala 117:10]
  wire  _GEN_6973; // @[Execute.scala 117:10]
  wire  _GEN_6974; // @[Execute.scala 117:10]
  wire  _GEN_6975; // @[Execute.scala 117:10]
  wire  _GEN_6976; // @[Execute.scala 117:10]
  wire  _GEN_6977; // @[Execute.scala 117:10]
  wire  _GEN_6979; // @[Execute.scala 117:10]
  wire  _GEN_6980; // @[Execute.scala 117:10]
  wire  _GEN_6981; // @[Execute.scala 117:10]
  wire  _GEN_6982; // @[Execute.scala 117:10]
  wire  _GEN_6983; // @[Execute.scala 117:10]
  wire  _GEN_6984; // @[Execute.scala 117:10]
  wire  _GEN_6985; // @[Execute.scala 117:10]
  wire  _GEN_6986; // @[Execute.scala 117:10]
  wire  _GEN_6987; // @[Execute.scala 117:10]
  wire  _GEN_6988; // @[Execute.scala 117:10]
  wire  _GEN_6989; // @[Execute.scala 117:10]
  wire  _GEN_6990; // @[Execute.scala 117:10]
  wire  _GEN_6991; // @[Execute.scala 117:10]
  wire  _GEN_6992; // @[Execute.scala 117:10]
  wire  _GEN_6993; // @[Execute.scala 117:10]
  wire  _GEN_6994; // @[Execute.scala 117:10]
  wire  _GEN_6995; // @[Execute.scala 117:10]
  wire  _GEN_6996; // @[Execute.scala 117:10]
  wire  _GEN_6997; // @[Execute.scala 117:10]
  wire  _GEN_6998; // @[Execute.scala 117:10]
  wire  _GEN_6999; // @[Execute.scala 117:10]
  wire  _GEN_7000; // @[Execute.scala 117:10]
  wire  _GEN_7001; // @[Execute.scala 117:10]
  wire  _GEN_7002; // @[Execute.scala 117:10]
  wire  _GEN_7003; // @[Execute.scala 117:10]
  wire  _GEN_7004; // @[Execute.scala 117:10]
  wire  _GEN_7005; // @[Execute.scala 117:10]
  wire  _GEN_7006; // @[Execute.scala 117:10]
  wire  _GEN_7007; // @[Execute.scala 117:10]
  wire  _GEN_7008; // @[Execute.scala 117:10]
  wire  _GEN_7009; // @[Execute.scala 117:10]
  wire  _GEN_7010; // @[Execute.scala 117:10]
  wire  _GEN_7011; // @[Execute.scala 117:10]
  wire  _GEN_7012; // @[Execute.scala 117:10]
  wire  _GEN_7013; // @[Execute.scala 117:10]
  wire  _GEN_7014; // @[Execute.scala 117:10]
  wire  _GEN_7015; // @[Execute.scala 117:10]
  wire  _GEN_7016; // @[Execute.scala 117:10]
  wire  _GEN_7017; // @[Execute.scala 117:10]
  wire  _GEN_7018; // @[Execute.scala 117:10]
  wire  _GEN_7019; // @[Execute.scala 117:10]
  wire  _GEN_7020; // @[Execute.scala 117:10]
  wire  _GEN_7021; // @[Execute.scala 117:10]
  wire  _GEN_7022; // @[Execute.scala 117:10]
  wire  _GEN_7023; // @[Execute.scala 117:10]
  wire  _GEN_7024; // @[Execute.scala 117:10]
  wire  _GEN_7025; // @[Execute.scala 117:10]
  wire  _GEN_7026; // @[Execute.scala 117:10]
  wire  _GEN_7027; // @[Execute.scala 117:10]
  wire  _GEN_7028; // @[Execute.scala 117:10]
  wire  _GEN_7029; // @[Execute.scala 117:10]
  wire  _GEN_7030; // @[Execute.scala 117:10]
  wire  _GEN_7031; // @[Execute.scala 117:10]
  wire  _GEN_7032; // @[Execute.scala 117:10]
  wire  _GEN_7033; // @[Execute.scala 117:10]
  wire  _GEN_7034; // @[Execute.scala 117:10]
  wire  _GEN_7035; // @[Execute.scala 117:10]
  wire  _GEN_7036; // @[Execute.scala 117:10]
  wire  _GEN_7037; // @[Execute.scala 117:10]
  wire  _GEN_7038; // @[Execute.scala 117:10]
  wire  _GEN_7039; // @[Execute.scala 117:10]
  wire  _GEN_7040; // @[Execute.scala 117:10]
  wire  _GEN_7041; // @[Execute.scala 117:10]
  wire  _T_631; // @[Execute.scala 117:10]
  wire  _T_632; // @[Execute.scala 117:15]
  wire [5:0] _T_634; // @[Execute.scala 117:37]
  wire [5:0] _T_638; // @[Execute.scala 117:60]
  wire  _GEN_7043; // @[Execute.scala 117:10]
  wire  _GEN_7044; // @[Execute.scala 117:10]
  wire  _GEN_7045; // @[Execute.scala 117:10]
  wire  _GEN_7046; // @[Execute.scala 117:10]
  wire  _GEN_7047; // @[Execute.scala 117:10]
  wire  _GEN_7048; // @[Execute.scala 117:10]
  wire  _GEN_7049; // @[Execute.scala 117:10]
  wire  _GEN_7050; // @[Execute.scala 117:10]
  wire  _GEN_7051; // @[Execute.scala 117:10]
  wire  _GEN_7052; // @[Execute.scala 117:10]
  wire  _GEN_7053; // @[Execute.scala 117:10]
  wire  _GEN_7054; // @[Execute.scala 117:10]
  wire  _GEN_7055; // @[Execute.scala 117:10]
  wire  _GEN_7056; // @[Execute.scala 117:10]
  wire  _GEN_7057; // @[Execute.scala 117:10]
  wire  _GEN_7058; // @[Execute.scala 117:10]
  wire  _GEN_7059; // @[Execute.scala 117:10]
  wire  _GEN_7060; // @[Execute.scala 117:10]
  wire  _GEN_7061; // @[Execute.scala 117:10]
  wire  _GEN_7062; // @[Execute.scala 117:10]
  wire  _GEN_7063; // @[Execute.scala 117:10]
  wire  _GEN_7064; // @[Execute.scala 117:10]
  wire  _GEN_7065; // @[Execute.scala 117:10]
  wire  _GEN_7066; // @[Execute.scala 117:10]
  wire  _GEN_7067; // @[Execute.scala 117:10]
  wire  _GEN_7068; // @[Execute.scala 117:10]
  wire  _GEN_7069; // @[Execute.scala 117:10]
  wire  _GEN_7070; // @[Execute.scala 117:10]
  wire  _GEN_7071; // @[Execute.scala 117:10]
  wire  _GEN_7072; // @[Execute.scala 117:10]
  wire  _GEN_7073; // @[Execute.scala 117:10]
  wire  _GEN_7074; // @[Execute.scala 117:10]
  wire  _GEN_7075; // @[Execute.scala 117:10]
  wire  _GEN_7076; // @[Execute.scala 117:10]
  wire  _GEN_7077; // @[Execute.scala 117:10]
  wire  _GEN_7078; // @[Execute.scala 117:10]
  wire  _GEN_7079; // @[Execute.scala 117:10]
  wire  _GEN_7080; // @[Execute.scala 117:10]
  wire  _GEN_7081; // @[Execute.scala 117:10]
  wire  _GEN_7082; // @[Execute.scala 117:10]
  wire  _GEN_7083; // @[Execute.scala 117:10]
  wire  _GEN_7084; // @[Execute.scala 117:10]
  wire  _GEN_7085; // @[Execute.scala 117:10]
  wire  _GEN_7086; // @[Execute.scala 117:10]
  wire  _GEN_7087; // @[Execute.scala 117:10]
  wire  _GEN_7088; // @[Execute.scala 117:10]
  wire  _GEN_7089; // @[Execute.scala 117:10]
  wire  _GEN_7090; // @[Execute.scala 117:10]
  wire  _GEN_7091; // @[Execute.scala 117:10]
  wire  _GEN_7092; // @[Execute.scala 117:10]
  wire  _GEN_7093; // @[Execute.scala 117:10]
  wire  _GEN_7094; // @[Execute.scala 117:10]
  wire  _GEN_7095; // @[Execute.scala 117:10]
  wire  _GEN_7096; // @[Execute.scala 117:10]
  wire  _GEN_7097; // @[Execute.scala 117:10]
  wire  _GEN_7098; // @[Execute.scala 117:10]
  wire  _GEN_7099; // @[Execute.scala 117:10]
  wire  _GEN_7100; // @[Execute.scala 117:10]
  wire  _GEN_7101; // @[Execute.scala 117:10]
  wire  _GEN_7102; // @[Execute.scala 117:10]
  wire  _GEN_7103; // @[Execute.scala 117:10]
  wire  _GEN_7104; // @[Execute.scala 117:10]
  wire  _GEN_7105; // @[Execute.scala 117:10]
  wire  _GEN_7107; // @[Execute.scala 117:10]
  wire  _GEN_7108; // @[Execute.scala 117:10]
  wire  _GEN_7109; // @[Execute.scala 117:10]
  wire  _GEN_7110; // @[Execute.scala 117:10]
  wire  _GEN_7111; // @[Execute.scala 117:10]
  wire  _GEN_7112; // @[Execute.scala 117:10]
  wire  _GEN_7113; // @[Execute.scala 117:10]
  wire  _GEN_7114; // @[Execute.scala 117:10]
  wire  _GEN_7115; // @[Execute.scala 117:10]
  wire  _GEN_7116; // @[Execute.scala 117:10]
  wire  _GEN_7117; // @[Execute.scala 117:10]
  wire  _GEN_7118; // @[Execute.scala 117:10]
  wire  _GEN_7119; // @[Execute.scala 117:10]
  wire  _GEN_7120; // @[Execute.scala 117:10]
  wire  _GEN_7121; // @[Execute.scala 117:10]
  wire  _GEN_7122; // @[Execute.scala 117:10]
  wire  _GEN_7123; // @[Execute.scala 117:10]
  wire  _GEN_7124; // @[Execute.scala 117:10]
  wire  _GEN_7125; // @[Execute.scala 117:10]
  wire  _GEN_7126; // @[Execute.scala 117:10]
  wire  _GEN_7127; // @[Execute.scala 117:10]
  wire  _GEN_7128; // @[Execute.scala 117:10]
  wire  _GEN_7129; // @[Execute.scala 117:10]
  wire  _GEN_7130; // @[Execute.scala 117:10]
  wire  _GEN_7131; // @[Execute.scala 117:10]
  wire  _GEN_7132; // @[Execute.scala 117:10]
  wire  _GEN_7133; // @[Execute.scala 117:10]
  wire  _GEN_7134; // @[Execute.scala 117:10]
  wire  _GEN_7135; // @[Execute.scala 117:10]
  wire  _GEN_7136; // @[Execute.scala 117:10]
  wire  _GEN_7137; // @[Execute.scala 117:10]
  wire  _GEN_7138; // @[Execute.scala 117:10]
  wire  _GEN_7139; // @[Execute.scala 117:10]
  wire  _GEN_7140; // @[Execute.scala 117:10]
  wire  _GEN_7141; // @[Execute.scala 117:10]
  wire  _GEN_7142; // @[Execute.scala 117:10]
  wire  _GEN_7143; // @[Execute.scala 117:10]
  wire  _GEN_7144; // @[Execute.scala 117:10]
  wire  _GEN_7145; // @[Execute.scala 117:10]
  wire  _GEN_7146; // @[Execute.scala 117:10]
  wire  _GEN_7147; // @[Execute.scala 117:10]
  wire  _GEN_7148; // @[Execute.scala 117:10]
  wire  _GEN_7149; // @[Execute.scala 117:10]
  wire  _GEN_7150; // @[Execute.scala 117:10]
  wire  _GEN_7151; // @[Execute.scala 117:10]
  wire  _GEN_7152; // @[Execute.scala 117:10]
  wire  _GEN_7153; // @[Execute.scala 117:10]
  wire  _GEN_7154; // @[Execute.scala 117:10]
  wire  _GEN_7155; // @[Execute.scala 117:10]
  wire  _GEN_7156; // @[Execute.scala 117:10]
  wire  _GEN_7157; // @[Execute.scala 117:10]
  wire  _GEN_7158; // @[Execute.scala 117:10]
  wire  _GEN_7159; // @[Execute.scala 117:10]
  wire  _GEN_7160; // @[Execute.scala 117:10]
  wire  _GEN_7161; // @[Execute.scala 117:10]
  wire  _GEN_7162; // @[Execute.scala 117:10]
  wire  _GEN_7163; // @[Execute.scala 117:10]
  wire  _GEN_7164; // @[Execute.scala 117:10]
  wire  _GEN_7165; // @[Execute.scala 117:10]
  wire  _GEN_7166; // @[Execute.scala 117:10]
  wire  _GEN_7167; // @[Execute.scala 117:10]
  wire  _GEN_7168; // @[Execute.scala 117:10]
  wire  _GEN_7169; // @[Execute.scala 117:10]
  wire  _T_641; // @[Execute.scala 117:10]
  wire  _T_642; // @[Execute.scala 117:15]
  wire [5:0] _T_644; // @[Execute.scala 117:37]
  wire [5:0] _T_648; // @[Execute.scala 117:60]
  wire  _GEN_7171; // @[Execute.scala 117:10]
  wire  _GEN_7172; // @[Execute.scala 117:10]
  wire  _GEN_7173; // @[Execute.scala 117:10]
  wire  _GEN_7174; // @[Execute.scala 117:10]
  wire  _GEN_7175; // @[Execute.scala 117:10]
  wire  _GEN_7176; // @[Execute.scala 117:10]
  wire  _GEN_7177; // @[Execute.scala 117:10]
  wire  _GEN_7178; // @[Execute.scala 117:10]
  wire  _GEN_7179; // @[Execute.scala 117:10]
  wire  _GEN_7180; // @[Execute.scala 117:10]
  wire  _GEN_7181; // @[Execute.scala 117:10]
  wire  _GEN_7182; // @[Execute.scala 117:10]
  wire  _GEN_7183; // @[Execute.scala 117:10]
  wire  _GEN_7184; // @[Execute.scala 117:10]
  wire  _GEN_7185; // @[Execute.scala 117:10]
  wire  _GEN_7186; // @[Execute.scala 117:10]
  wire  _GEN_7187; // @[Execute.scala 117:10]
  wire  _GEN_7188; // @[Execute.scala 117:10]
  wire  _GEN_7189; // @[Execute.scala 117:10]
  wire  _GEN_7190; // @[Execute.scala 117:10]
  wire  _GEN_7191; // @[Execute.scala 117:10]
  wire  _GEN_7192; // @[Execute.scala 117:10]
  wire  _GEN_7193; // @[Execute.scala 117:10]
  wire  _GEN_7194; // @[Execute.scala 117:10]
  wire  _GEN_7195; // @[Execute.scala 117:10]
  wire  _GEN_7196; // @[Execute.scala 117:10]
  wire  _GEN_7197; // @[Execute.scala 117:10]
  wire  _GEN_7198; // @[Execute.scala 117:10]
  wire  _GEN_7199; // @[Execute.scala 117:10]
  wire  _GEN_7200; // @[Execute.scala 117:10]
  wire  _GEN_7201; // @[Execute.scala 117:10]
  wire  _GEN_7202; // @[Execute.scala 117:10]
  wire  _GEN_7203; // @[Execute.scala 117:10]
  wire  _GEN_7204; // @[Execute.scala 117:10]
  wire  _GEN_7205; // @[Execute.scala 117:10]
  wire  _GEN_7206; // @[Execute.scala 117:10]
  wire  _GEN_7207; // @[Execute.scala 117:10]
  wire  _GEN_7208; // @[Execute.scala 117:10]
  wire  _GEN_7209; // @[Execute.scala 117:10]
  wire  _GEN_7210; // @[Execute.scala 117:10]
  wire  _GEN_7211; // @[Execute.scala 117:10]
  wire  _GEN_7212; // @[Execute.scala 117:10]
  wire  _GEN_7213; // @[Execute.scala 117:10]
  wire  _GEN_7214; // @[Execute.scala 117:10]
  wire  _GEN_7215; // @[Execute.scala 117:10]
  wire  _GEN_7216; // @[Execute.scala 117:10]
  wire  _GEN_7217; // @[Execute.scala 117:10]
  wire  _GEN_7218; // @[Execute.scala 117:10]
  wire  _GEN_7219; // @[Execute.scala 117:10]
  wire  _GEN_7220; // @[Execute.scala 117:10]
  wire  _GEN_7221; // @[Execute.scala 117:10]
  wire  _GEN_7222; // @[Execute.scala 117:10]
  wire  _GEN_7223; // @[Execute.scala 117:10]
  wire  _GEN_7224; // @[Execute.scala 117:10]
  wire  _GEN_7225; // @[Execute.scala 117:10]
  wire  _GEN_7226; // @[Execute.scala 117:10]
  wire  _GEN_7227; // @[Execute.scala 117:10]
  wire  _GEN_7228; // @[Execute.scala 117:10]
  wire  _GEN_7229; // @[Execute.scala 117:10]
  wire  _GEN_7230; // @[Execute.scala 117:10]
  wire  _GEN_7231; // @[Execute.scala 117:10]
  wire  _GEN_7232; // @[Execute.scala 117:10]
  wire  _GEN_7233; // @[Execute.scala 117:10]
  wire  _GEN_7235; // @[Execute.scala 117:10]
  wire  _GEN_7236; // @[Execute.scala 117:10]
  wire  _GEN_7237; // @[Execute.scala 117:10]
  wire  _GEN_7238; // @[Execute.scala 117:10]
  wire  _GEN_7239; // @[Execute.scala 117:10]
  wire  _GEN_7240; // @[Execute.scala 117:10]
  wire  _GEN_7241; // @[Execute.scala 117:10]
  wire  _GEN_7242; // @[Execute.scala 117:10]
  wire  _GEN_7243; // @[Execute.scala 117:10]
  wire  _GEN_7244; // @[Execute.scala 117:10]
  wire  _GEN_7245; // @[Execute.scala 117:10]
  wire  _GEN_7246; // @[Execute.scala 117:10]
  wire  _GEN_7247; // @[Execute.scala 117:10]
  wire  _GEN_7248; // @[Execute.scala 117:10]
  wire  _GEN_7249; // @[Execute.scala 117:10]
  wire  _GEN_7250; // @[Execute.scala 117:10]
  wire  _GEN_7251; // @[Execute.scala 117:10]
  wire  _GEN_7252; // @[Execute.scala 117:10]
  wire  _GEN_7253; // @[Execute.scala 117:10]
  wire  _GEN_7254; // @[Execute.scala 117:10]
  wire  _GEN_7255; // @[Execute.scala 117:10]
  wire  _GEN_7256; // @[Execute.scala 117:10]
  wire  _GEN_7257; // @[Execute.scala 117:10]
  wire  _GEN_7258; // @[Execute.scala 117:10]
  wire  _GEN_7259; // @[Execute.scala 117:10]
  wire  _GEN_7260; // @[Execute.scala 117:10]
  wire  _GEN_7261; // @[Execute.scala 117:10]
  wire  _GEN_7262; // @[Execute.scala 117:10]
  wire  _GEN_7263; // @[Execute.scala 117:10]
  wire  _GEN_7264; // @[Execute.scala 117:10]
  wire  _GEN_7265; // @[Execute.scala 117:10]
  wire  _GEN_7266; // @[Execute.scala 117:10]
  wire  _GEN_7267; // @[Execute.scala 117:10]
  wire  _GEN_7268; // @[Execute.scala 117:10]
  wire  _GEN_7269; // @[Execute.scala 117:10]
  wire  _GEN_7270; // @[Execute.scala 117:10]
  wire  _GEN_7271; // @[Execute.scala 117:10]
  wire  _GEN_7272; // @[Execute.scala 117:10]
  wire  _GEN_7273; // @[Execute.scala 117:10]
  wire  _GEN_7274; // @[Execute.scala 117:10]
  wire  _GEN_7275; // @[Execute.scala 117:10]
  wire  _GEN_7276; // @[Execute.scala 117:10]
  wire  _GEN_7277; // @[Execute.scala 117:10]
  wire  _GEN_7278; // @[Execute.scala 117:10]
  wire  _GEN_7279; // @[Execute.scala 117:10]
  wire  _GEN_7280; // @[Execute.scala 117:10]
  wire  _GEN_7281; // @[Execute.scala 117:10]
  wire  _GEN_7282; // @[Execute.scala 117:10]
  wire  _GEN_7283; // @[Execute.scala 117:10]
  wire  _GEN_7284; // @[Execute.scala 117:10]
  wire  _GEN_7285; // @[Execute.scala 117:10]
  wire  _GEN_7286; // @[Execute.scala 117:10]
  wire  _GEN_7287; // @[Execute.scala 117:10]
  wire  _GEN_7288; // @[Execute.scala 117:10]
  wire  _GEN_7289; // @[Execute.scala 117:10]
  wire  _GEN_7290; // @[Execute.scala 117:10]
  wire  _GEN_7291; // @[Execute.scala 117:10]
  wire  _GEN_7292; // @[Execute.scala 117:10]
  wire  _GEN_7293; // @[Execute.scala 117:10]
  wire  _GEN_7294; // @[Execute.scala 117:10]
  wire  _GEN_7295; // @[Execute.scala 117:10]
  wire  _GEN_7296; // @[Execute.scala 117:10]
  wire  _GEN_7297; // @[Execute.scala 117:10]
  wire  _T_651; // @[Execute.scala 117:10]
  wire  _T_652; // @[Execute.scala 117:15]
  wire [5:0] _T_654; // @[Execute.scala 117:37]
  wire [5:0] _T_658; // @[Execute.scala 117:60]
  wire  _GEN_7299; // @[Execute.scala 117:10]
  wire  _GEN_7300; // @[Execute.scala 117:10]
  wire  _GEN_7301; // @[Execute.scala 117:10]
  wire  _GEN_7302; // @[Execute.scala 117:10]
  wire  _GEN_7303; // @[Execute.scala 117:10]
  wire  _GEN_7304; // @[Execute.scala 117:10]
  wire  _GEN_7305; // @[Execute.scala 117:10]
  wire  _GEN_7306; // @[Execute.scala 117:10]
  wire  _GEN_7307; // @[Execute.scala 117:10]
  wire  _GEN_7308; // @[Execute.scala 117:10]
  wire  _GEN_7309; // @[Execute.scala 117:10]
  wire  _GEN_7310; // @[Execute.scala 117:10]
  wire  _GEN_7311; // @[Execute.scala 117:10]
  wire  _GEN_7312; // @[Execute.scala 117:10]
  wire  _GEN_7313; // @[Execute.scala 117:10]
  wire  _GEN_7314; // @[Execute.scala 117:10]
  wire  _GEN_7315; // @[Execute.scala 117:10]
  wire  _GEN_7316; // @[Execute.scala 117:10]
  wire  _GEN_7317; // @[Execute.scala 117:10]
  wire  _GEN_7318; // @[Execute.scala 117:10]
  wire  _GEN_7319; // @[Execute.scala 117:10]
  wire  _GEN_7320; // @[Execute.scala 117:10]
  wire  _GEN_7321; // @[Execute.scala 117:10]
  wire  _GEN_7322; // @[Execute.scala 117:10]
  wire  _GEN_7323; // @[Execute.scala 117:10]
  wire  _GEN_7324; // @[Execute.scala 117:10]
  wire  _GEN_7325; // @[Execute.scala 117:10]
  wire  _GEN_7326; // @[Execute.scala 117:10]
  wire  _GEN_7327; // @[Execute.scala 117:10]
  wire  _GEN_7328; // @[Execute.scala 117:10]
  wire  _GEN_7329; // @[Execute.scala 117:10]
  wire  _GEN_7330; // @[Execute.scala 117:10]
  wire  _GEN_7331; // @[Execute.scala 117:10]
  wire  _GEN_7332; // @[Execute.scala 117:10]
  wire  _GEN_7333; // @[Execute.scala 117:10]
  wire  _GEN_7334; // @[Execute.scala 117:10]
  wire  _GEN_7335; // @[Execute.scala 117:10]
  wire  _GEN_7336; // @[Execute.scala 117:10]
  wire  _GEN_7337; // @[Execute.scala 117:10]
  wire  _GEN_7338; // @[Execute.scala 117:10]
  wire  _GEN_7339; // @[Execute.scala 117:10]
  wire  _GEN_7340; // @[Execute.scala 117:10]
  wire  _GEN_7341; // @[Execute.scala 117:10]
  wire  _GEN_7342; // @[Execute.scala 117:10]
  wire  _GEN_7343; // @[Execute.scala 117:10]
  wire  _GEN_7344; // @[Execute.scala 117:10]
  wire  _GEN_7345; // @[Execute.scala 117:10]
  wire  _GEN_7346; // @[Execute.scala 117:10]
  wire  _GEN_7347; // @[Execute.scala 117:10]
  wire  _GEN_7348; // @[Execute.scala 117:10]
  wire  _GEN_7349; // @[Execute.scala 117:10]
  wire  _GEN_7350; // @[Execute.scala 117:10]
  wire  _GEN_7351; // @[Execute.scala 117:10]
  wire  _GEN_7352; // @[Execute.scala 117:10]
  wire  _GEN_7353; // @[Execute.scala 117:10]
  wire  _GEN_7354; // @[Execute.scala 117:10]
  wire  _GEN_7355; // @[Execute.scala 117:10]
  wire  _GEN_7356; // @[Execute.scala 117:10]
  wire  _GEN_7357; // @[Execute.scala 117:10]
  wire  _GEN_7358; // @[Execute.scala 117:10]
  wire  _GEN_7359; // @[Execute.scala 117:10]
  wire  _GEN_7360; // @[Execute.scala 117:10]
  wire  _GEN_7361; // @[Execute.scala 117:10]
  wire  _GEN_7363; // @[Execute.scala 117:10]
  wire  _GEN_7364; // @[Execute.scala 117:10]
  wire  _GEN_7365; // @[Execute.scala 117:10]
  wire  _GEN_7366; // @[Execute.scala 117:10]
  wire  _GEN_7367; // @[Execute.scala 117:10]
  wire  _GEN_7368; // @[Execute.scala 117:10]
  wire  _GEN_7369; // @[Execute.scala 117:10]
  wire  _GEN_7370; // @[Execute.scala 117:10]
  wire  _GEN_7371; // @[Execute.scala 117:10]
  wire  _GEN_7372; // @[Execute.scala 117:10]
  wire  _GEN_7373; // @[Execute.scala 117:10]
  wire  _GEN_7374; // @[Execute.scala 117:10]
  wire  _GEN_7375; // @[Execute.scala 117:10]
  wire  _GEN_7376; // @[Execute.scala 117:10]
  wire  _GEN_7377; // @[Execute.scala 117:10]
  wire  _GEN_7378; // @[Execute.scala 117:10]
  wire  _GEN_7379; // @[Execute.scala 117:10]
  wire  _GEN_7380; // @[Execute.scala 117:10]
  wire  _GEN_7381; // @[Execute.scala 117:10]
  wire  _GEN_7382; // @[Execute.scala 117:10]
  wire  _GEN_7383; // @[Execute.scala 117:10]
  wire  _GEN_7384; // @[Execute.scala 117:10]
  wire  _GEN_7385; // @[Execute.scala 117:10]
  wire  _GEN_7386; // @[Execute.scala 117:10]
  wire  _GEN_7387; // @[Execute.scala 117:10]
  wire  _GEN_7388; // @[Execute.scala 117:10]
  wire  _GEN_7389; // @[Execute.scala 117:10]
  wire  _GEN_7390; // @[Execute.scala 117:10]
  wire  _GEN_7391; // @[Execute.scala 117:10]
  wire  _GEN_7392; // @[Execute.scala 117:10]
  wire  _GEN_7393; // @[Execute.scala 117:10]
  wire  _GEN_7394; // @[Execute.scala 117:10]
  wire  _GEN_7395; // @[Execute.scala 117:10]
  wire  _GEN_7396; // @[Execute.scala 117:10]
  wire  _GEN_7397; // @[Execute.scala 117:10]
  wire  _GEN_7398; // @[Execute.scala 117:10]
  wire  _GEN_7399; // @[Execute.scala 117:10]
  wire  _GEN_7400; // @[Execute.scala 117:10]
  wire  _GEN_7401; // @[Execute.scala 117:10]
  wire  _GEN_7402; // @[Execute.scala 117:10]
  wire  _GEN_7403; // @[Execute.scala 117:10]
  wire  _GEN_7404; // @[Execute.scala 117:10]
  wire  _GEN_7405; // @[Execute.scala 117:10]
  wire  _GEN_7406; // @[Execute.scala 117:10]
  wire  _GEN_7407; // @[Execute.scala 117:10]
  wire  _GEN_7408; // @[Execute.scala 117:10]
  wire  _GEN_7409; // @[Execute.scala 117:10]
  wire  _GEN_7410; // @[Execute.scala 117:10]
  wire  _GEN_7411; // @[Execute.scala 117:10]
  wire  _GEN_7412; // @[Execute.scala 117:10]
  wire  _GEN_7413; // @[Execute.scala 117:10]
  wire  _GEN_7414; // @[Execute.scala 117:10]
  wire  _GEN_7415; // @[Execute.scala 117:10]
  wire  _GEN_7416; // @[Execute.scala 117:10]
  wire  _GEN_7417; // @[Execute.scala 117:10]
  wire  _GEN_7418; // @[Execute.scala 117:10]
  wire  _GEN_7419; // @[Execute.scala 117:10]
  wire  _GEN_7420; // @[Execute.scala 117:10]
  wire  _GEN_7421; // @[Execute.scala 117:10]
  wire  _GEN_7422; // @[Execute.scala 117:10]
  wire  _GEN_7423; // @[Execute.scala 117:10]
  wire  _GEN_7424; // @[Execute.scala 117:10]
  wire  _GEN_7425; // @[Execute.scala 117:10]
  wire  _T_661; // @[Execute.scala 117:10]
  wire  _T_662; // @[Execute.scala 117:15]
  wire [5:0] _T_664; // @[Execute.scala 117:37]
  wire [5:0] _T_668; // @[Execute.scala 117:60]
  wire  _GEN_7427; // @[Execute.scala 117:10]
  wire  _GEN_7428; // @[Execute.scala 117:10]
  wire  _GEN_7429; // @[Execute.scala 117:10]
  wire  _GEN_7430; // @[Execute.scala 117:10]
  wire  _GEN_7431; // @[Execute.scala 117:10]
  wire  _GEN_7432; // @[Execute.scala 117:10]
  wire  _GEN_7433; // @[Execute.scala 117:10]
  wire  _GEN_7434; // @[Execute.scala 117:10]
  wire  _GEN_7435; // @[Execute.scala 117:10]
  wire  _GEN_7436; // @[Execute.scala 117:10]
  wire  _GEN_7437; // @[Execute.scala 117:10]
  wire  _GEN_7438; // @[Execute.scala 117:10]
  wire  _GEN_7439; // @[Execute.scala 117:10]
  wire  _GEN_7440; // @[Execute.scala 117:10]
  wire  _GEN_7441; // @[Execute.scala 117:10]
  wire  _GEN_7442; // @[Execute.scala 117:10]
  wire  _GEN_7443; // @[Execute.scala 117:10]
  wire  _GEN_7444; // @[Execute.scala 117:10]
  wire  _GEN_7445; // @[Execute.scala 117:10]
  wire  _GEN_7446; // @[Execute.scala 117:10]
  wire  _GEN_7447; // @[Execute.scala 117:10]
  wire  _GEN_7448; // @[Execute.scala 117:10]
  wire  _GEN_7449; // @[Execute.scala 117:10]
  wire  _GEN_7450; // @[Execute.scala 117:10]
  wire  _GEN_7451; // @[Execute.scala 117:10]
  wire  _GEN_7452; // @[Execute.scala 117:10]
  wire  _GEN_7453; // @[Execute.scala 117:10]
  wire  _GEN_7454; // @[Execute.scala 117:10]
  wire  _GEN_7455; // @[Execute.scala 117:10]
  wire  _GEN_7456; // @[Execute.scala 117:10]
  wire  _GEN_7457; // @[Execute.scala 117:10]
  wire  _GEN_7458; // @[Execute.scala 117:10]
  wire  _GEN_7459; // @[Execute.scala 117:10]
  wire  _GEN_7460; // @[Execute.scala 117:10]
  wire  _GEN_7461; // @[Execute.scala 117:10]
  wire  _GEN_7462; // @[Execute.scala 117:10]
  wire  _GEN_7463; // @[Execute.scala 117:10]
  wire  _GEN_7464; // @[Execute.scala 117:10]
  wire  _GEN_7465; // @[Execute.scala 117:10]
  wire  _GEN_7466; // @[Execute.scala 117:10]
  wire  _GEN_7467; // @[Execute.scala 117:10]
  wire  _GEN_7468; // @[Execute.scala 117:10]
  wire  _GEN_7469; // @[Execute.scala 117:10]
  wire  _GEN_7470; // @[Execute.scala 117:10]
  wire  _GEN_7471; // @[Execute.scala 117:10]
  wire  _GEN_7472; // @[Execute.scala 117:10]
  wire  _GEN_7473; // @[Execute.scala 117:10]
  wire  _GEN_7474; // @[Execute.scala 117:10]
  wire  _GEN_7475; // @[Execute.scala 117:10]
  wire  _GEN_7476; // @[Execute.scala 117:10]
  wire  _GEN_7477; // @[Execute.scala 117:10]
  wire  _GEN_7478; // @[Execute.scala 117:10]
  wire  _GEN_7479; // @[Execute.scala 117:10]
  wire  _GEN_7480; // @[Execute.scala 117:10]
  wire  _GEN_7481; // @[Execute.scala 117:10]
  wire  _GEN_7482; // @[Execute.scala 117:10]
  wire  _GEN_7483; // @[Execute.scala 117:10]
  wire  _GEN_7484; // @[Execute.scala 117:10]
  wire  _GEN_7485; // @[Execute.scala 117:10]
  wire  _GEN_7486; // @[Execute.scala 117:10]
  wire  _GEN_7487; // @[Execute.scala 117:10]
  wire  _GEN_7488; // @[Execute.scala 117:10]
  wire  _GEN_7489; // @[Execute.scala 117:10]
  wire  _GEN_7491; // @[Execute.scala 117:10]
  wire  _GEN_7492; // @[Execute.scala 117:10]
  wire  _GEN_7493; // @[Execute.scala 117:10]
  wire  _GEN_7494; // @[Execute.scala 117:10]
  wire  _GEN_7495; // @[Execute.scala 117:10]
  wire  _GEN_7496; // @[Execute.scala 117:10]
  wire  _GEN_7497; // @[Execute.scala 117:10]
  wire  _GEN_7498; // @[Execute.scala 117:10]
  wire  _GEN_7499; // @[Execute.scala 117:10]
  wire  _GEN_7500; // @[Execute.scala 117:10]
  wire  _GEN_7501; // @[Execute.scala 117:10]
  wire  _GEN_7502; // @[Execute.scala 117:10]
  wire  _GEN_7503; // @[Execute.scala 117:10]
  wire  _GEN_7504; // @[Execute.scala 117:10]
  wire  _GEN_7505; // @[Execute.scala 117:10]
  wire  _GEN_7506; // @[Execute.scala 117:10]
  wire  _GEN_7507; // @[Execute.scala 117:10]
  wire  _GEN_7508; // @[Execute.scala 117:10]
  wire  _GEN_7509; // @[Execute.scala 117:10]
  wire  _GEN_7510; // @[Execute.scala 117:10]
  wire  _GEN_7511; // @[Execute.scala 117:10]
  wire  _GEN_7512; // @[Execute.scala 117:10]
  wire  _GEN_7513; // @[Execute.scala 117:10]
  wire  _GEN_7514; // @[Execute.scala 117:10]
  wire  _GEN_7515; // @[Execute.scala 117:10]
  wire  _GEN_7516; // @[Execute.scala 117:10]
  wire  _GEN_7517; // @[Execute.scala 117:10]
  wire  _GEN_7518; // @[Execute.scala 117:10]
  wire  _GEN_7519; // @[Execute.scala 117:10]
  wire  _GEN_7520; // @[Execute.scala 117:10]
  wire  _GEN_7521; // @[Execute.scala 117:10]
  wire  _GEN_7522; // @[Execute.scala 117:10]
  wire  _GEN_7523; // @[Execute.scala 117:10]
  wire  _GEN_7524; // @[Execute.scala 117:10]
  wire  _GEN_7525; // @[Execute.scala 117:10]
  wire  _GEN_7526; // @[Execute.scala 117:10]
  wire  _GEN_7527; // @[Execute.scala 117:10]
  wire  _GEN_7528; // @[Execute.scala 117:10]
  wire  _GEN_7529; // @[Execute.scala 117:10]
  wire  _GEN_7530; // @[Execute.scala 117:10]
  wire  _GEN_7531; // @[Execute.scala 117:10]
  wire  _GEN_7532; // @[Execute.scala 117:10]
  wire  _GEN_7533; // @[Execute.scala 117:10]
  wire  _GEN_7534; // @[Execute.scala 117:10]
  wire  _GEN_7535; // @[Execute.scala 117:10]
  wire  _GEN_7536; // @[Execute.scala 117:10]
  wire  _GEN_7537; // @[Execute.scala 117:10]
  wire  _GEN_7538; // @[Execute.scala 117:10]
  wire  _GEN_7539; // @[Execute.scala 117:10]
  wire  _GEN_7540; // @[Execute.scala 117:10]
  wire  _GEN_7541; // @[Execute.scala 117:10]
  wire  _GEN_7542; // @[Execute.scala 117:10]
  wire  _GEN_7543; // @[Execute.scala 117:10]
  wire  _GEN_7544; // @[Execute.scala 117:10]
  wire  _GEN_7545; // @[Execute.scala 117:10]
  wire  _GEN_7546; // @[Execute.scala 117:10]
  wire  _GEN_7547; // @[Execute.scala 117:10]
  wire  _GEN_7548; // @[Execute.scala 117:10]
  wire  _GEN_7549; // @[Execute.scala 117:10]
  wire  _GEN_7550; // @[Execute.scala 117:10]
  wire  _GEN_7551; // @[Execute.scala 117:10]
  wire  _GEN_7552; // @[Execute.scala 117:10]
  wire  _GEN_7553; // @[Execute.scala 117:10]
  wire  _T_671; // @[Execute.scala 117:10]
  wire  _T_672; // @[Execute.scala 117:15]
  wire [5:0] _T_674; // @[Execute.scala 117:37]
  wire [5:0] _T_678; // @[Execute.scala 117:60]
  wire  _GEN_7555; // @[Execute.scala 117:10]
  wire  _GEN_7556; // @[Execute.scala 117:10]
  wire  _GEN_7557; // @[Execute.scala 117:10]
  wire  _GEN_7558; // @[Execute.scala 117:10]
  wire  _GEN_7559; // @[Execute.scala 117:10]
  wire  _GEN_7560; // @[Execute.scala 117:10]
  wire  _GEN_7561; // @[Execute.scala 117:10]
  wire  _GEN_7562; // @[Execute.scala 117:10]
  wire  _GEN_7563; // @[Execute.scala 117:10]
  wire  _GEN_7564; // @[Execute.scala 117:10]
  wire  _GEN_7565; // @[Execute.scala 117:10]
  wire  _GEN_7566; // @[Execute.scala 117:10]
  wire  _GEN_7567; // @[Execute.scala 117:10]
  wire  _GEN_7568; // @[Execute.scala 117:10]
  wire  _GEN_7569; // @[Execute.scala 117:10]
  wire  _GEN_7570; // @[Execute.scala 117:10]
  wire  _GEN_7571; // @[Execute.scala 117:10]
  wire  _GEN_7572; // @[Execute.scala 117:10]
  wire  _GEN_7573; // @[Execute.scala 117:10]
  wire  _GEN_7574; // @[Execute.scala 117:10]
  wire  _GEN_7575; // @[Execute.scala 117:10]
  wire  _GEN_7576; // @[Execute.scala 117:10]
  wire  _GEN_7577; // @[Execute.scala 117:10]
  wire  _GEN_7578; // @[Execute.scala 117:10]
  wire  _GEN_7579; // @[Execute.scala 117:10]
  wire  _GEN_7580; // @[Execute.scala 117:10]
  wire  _GEN_7581; // @[Execute.scala 117:10]
  wire  _GEN_7582; // @[Execute.scala 117:10]
  wire  _GEN_7583; // @[Execute.scala 117:10]
  wire  _GEN_7584; // @[Execute.scala 117:10]
  wire  _GEN_7585; // @[Execute.scala 117:10]
  wire  _GEN_7586; // @[Execute.scala 117:10]
  wire  _GEN_7587; // @[Execute.scala 117:10]
  wire  _GEN_7588; // @[Execute.scala 117:10]
  wire  _GEN_7589; // @[Execute.scala 117:10]
  wire  _GEN_7590; // @[Execute.scala 117:10]
  wire  _GEN_7591; // @[Execute.scala 117:10]
  wire  _GEN_7592; // @[Execute.scala 117:10]
  wire  _GEN_7593; // @[Execute.scala 117:10]
  wire  _GEN_7594; // @[Execute.scala 117:10]
  wire  _GEN_7595; // @[Execute.scala 117:10]
  wire  _GEN_7596; // @[Execute.scala 117:10]
  wire  _GEN_7597; // @[Execute.scala 117:10]
  wire  _GEN_7598; // @[Execute.scala 117:10]
  wire  _GEN_7599; // @[Execute.scala 117:10]
  wire  _GEN_7600; // @[Execute.scala 117:10]
  wire  _GEN_7601; // @[Execute.scala 117:10]
  wire  _GEN_7602; // @[Execute.scala 117:10]
  wire  _GEN_7603; // @[Execute.scala 117:10]
  wire  _GEN_7604; // @[Execute.scala 117:10]
  wire  _GEN_7605; // @[Execute.scala 117:10]
  wire  _GEN_7606; // @[Execute.scala 117:10]
  wire  _GEN_7607; // @[Execute.scala 117:10]
  wire  _GEN_7608; // @[Execute.scala 117:10]
  wire  _GEN_7609; // @[Execute.scala 117:10]
  wire  _GEN_7610; // @[Execute.scala 117:10]
  wire  _GEN_7611; // @[Execute.scala 117:10]
  wire  _GEN_7612; // @[Execute.scala 117:10]
  wire  _GEN_7613; // @[Execute.scala 117:10]
  wire  _GEN_7614; // @[Execute.scala 117:10]
  wire  _GEN_7615; // @[Execute.scala 117:10]
  wire  _GEN_7616; // @[Execute.scala 117:10]
  wire  _GEN_7617; // @[Execute.scala 117:10]
  wire  _GEN_7619; // @[Execute.scala 117:10]
  wire  _GEN_7620; // @[Execute.scala 117:10]
  wire  _GEN_7621; // @[Execute.scala 117:10]
  wire  _GEN_7622; // @[Execute.scala 117:10]
  wire  _GEN_7623; // @[Execute.scala 117:10]
  wire  _GEN_7624; // @[Execute.scala 117:10]
  wire  _GEN_7625; // @[Execute.scala 117:10]
  wire  _GEN_7626; // @[Execute.scala 117:10]
  wire  _GEN_7627; // @[Execute.scala 117:10]
  wire  _GEN_7628; // @[Execute.scala 117:10]
  wire  _GEN_7629; // @[Execute.scala 117:10]
  wire  _GEN_7630; // @[Execute.scala 117:10]
  wire  _GEN_7631; // @[Execute.scala 117:10]
  wire  _GEN_7632; // @[Execute.scala 117:10]
  wire  _GEN_7633; // @[Execute.scala 117:10]
  wire  _GEN_7634; // @[Execute.scala 117:10]
  wire  _GEN_7635; // @[Execute.scala 117:10]
  wire  _GEN_7636; // @[Execute.scala 117:10]
  wire  _GEN_7637; // @[Execute.scala 117:10]
  wire  _GEN_7638; // @[Execute.scala 117:10]
  wire  _GEN_7639; // @[Execute.scala 117:10]
  wire  _GEN_7640; // @[Execute.scala 117:10]
  wire  _GEN_7641; // @[Execute.scala 117:10]
  wire  _GEN_7642; // @[Execute.scala 117:10]
  wire  _GEN_7643; // @[Execute.scala 117:10]
  wire  _GEN_7644; // @[Execute.scala 117:10]
  wire  _GEN_7645; // @[Execute.scala 117:10]
  wire  _GEN_7646; // @[Execute.scala 117:10]
  wire  _GEN_7647; // @[Execute.scala 117:10]
  wire  _GEN_7648; // @[Execute.scala 117:10]
  wire  _GEN_7649; // @[Execute.scala 117:10]
  wire  _GEN_7650; // @[Execute.scala 117:10]
  wire  _GEN_7651; // @[Execute.scala 117:10]
  wire  _GEN_7652; // @[Execute.scala 117:10]
  wire  _GEN_7653; // @[Execute.scala 117:10]
  wire  _GEN_7654; // @[Execute.scala 117:10]
  wire  _GEN_7655; // @[Execute.scala 117:10]
  wire  _GEN_7656; // @[Execute.scala 117:10]
  wire  _GEN_7657; // @[Execute.scala 117:10]
  wire  _GEN_7658; // @[Execute.scala 117:10]
  wire  _GEN_7659; // @[Execute.scala 117:10]
  wire  _GEN_7660; // @[Execute.scala 117:10]
  wire  _GEN_7661; // @[Execute.scala 117:10]
  wire  _GEN_7662; // @[Execute.scala 117:10]
  wire  _GEN_7663; // @[Execute.scala 117:10]
  wire  _GEN_7664; // @[Execute.scala 117:10]
  wire  _GEN_7665; // @[Execute.scala 117:10]
  wire  _GEN_7666; // @[Execute.scala 117:10]
  wire  _GEN_7667; // @[Execute.scala 117:10]
  wire  _GEN_7668; // @[Execute.scala 117:10]
  wire  _GEN_7669; // @[Execute.scala 117:10]
  wire  _GEN_7670; // @[Execute.scala 117:10]
  wire  _GEN_7671; // @[Execute.scala 117:10]
  wire  _GEN_7672; // @[Execute.scala 117:10]
  wire  _GEN_7673; // @[Execute.scala 117:10]
  wire  _GEN_7674; // @[Execute.scala 117:10]
  wire  _GEN_7675; // @[Execute.scala 117:10]
  wire  _GEN_7676; // @[Execute.scala 117:10]
  wire  _GEN_7677; // @[Execute.scala 117:10]
  wire  _GEN_7678; // @[Execute.scala 117:10]
  wire  _GEN_7679; // @[Execute.scala 117:10]
  wire  _GEN_7680; // @[Execute.scala 117:10]
  wire  _GEN_7681; // @[Execute.scala 117:10]
  wire  _T_681; // @[Execute.scala 117:10]
  wire  _T_682; // @[Execute.scala 117:15]
  wire [5:0] _T_684; // @[Execute.scala 117:37]
  wire [5:0] _T_688; // @[Execute.scala 117:60]
  wire  _GEN_7683; // @[Execute.scala 117:10]
  wire  _GEN_7684; // @[Execute.scala 117:10]
  wire  _GEN_7685; // @[Execute.scala 117:10]
  wire  _GEN_7686; // @[Execute.scala 117:10]
  wire  _GEN_7687; // @[Execute.scala 117:10]
  wire  _GEN_7688; // @[Execute.scala 117:10]
  wire  _GEN_7689; // @[Execute.scala 117:10]
  wire  _GEN_7690; // @[Execute.scala 117:10]
  wire  _GEN_7691; // @[Execute.scala 117:10]
  wire  _GEN_7692; // @[Execute.scala 117:10]
  wire  _GEN_7693; // @[Execute.scala 117:10]
  wire  _GEN_7694; // @[Execute.scala 117:10]
  wire  _GEN_7695; // @[Execute.scala 117:10]
  wire  _GEN_7696; // @[Execute.scala 117:10]
  wire  _GEN_7697; // @[Execute.scala 117:10]
  wire  _GEN_7698; // @[Execute.scala 117:10]
  wire  _GEN_7699; // @[Execute.scala 117:10]
  wire  _GEN_7700; // @[Execute.scala 117:10]
  wire  _GEN_7701; // @[Execute.scala 117:10]
  wire  _GEN_7702; // @[Execute.scala 117:10]
  wire  _GEN_7703; // @[Execute.scala 117:10]
  wire  _GEN_7704; // @[Execute.scala 117:10]
  wire  _GEN_7705; // @[Execute.scala 117:10]
  wire  _GEN_7706; // @[Execute.scala 117:10]
  wire  _GEN_7707; // @[Execute.scala 117:10]
  wire  _GEN_7708; // @[Execute.scala 117:10]
  wire  _GEN_7709; // @[Execute.scala 117:10]
  wire  _GEN_7710; // @[Execute.scala 117:10]
  wire  _GEN_7711; // @[Execute.scala 117:10]
  wire  _GEN_7712; // @[Execute.scala 117:10]
  wire  _GEN_7713; // @[Execute.scala 117:10]
  wire  _GEN_7714; // @[Execute.scala 117:10]
  wire  _GEN_7715; // @[Execute.scala 117:10]
  wire  _GEN_7716; // @[Execute.scala 117:10]
  wire  _GEN_7717; // @[Execute.scala 117:10]
  wire  _GEN_7718; // @[Execute.scala 117:10]
  wire  _GEN_7719; // @[Execute.scala 117:10]
  wire  _GEN_7720; // @[Execute.scala 117:10]
  wire  _GEN_7721; // @[Execute.scala 117:10]
  wire  _GEN_7722; // @[Execute.scala 117:10]
  wire  _GEN_7723; // @[Execute.scala 117:10]
  wire  _GEN_7724; // @[Execute.scala 117:10]
  wire  _GEN_7725; // @[Execute.scala 117:10]
  wire  _GEN_7726; // @[Execute.scala 117:10]
  wire  _GEN_7727; // @[Execute.scala 117:10]
  wire  _GEN_7728; // @[Execute.scala 117:10]
  wire  _GEN_7729; // @[Execute.scala 117:10]
  wire  _GEN_7730; // @[Execute.scala 117:10]
  wire  _GEN_7731; // @[Execute.scala 117:10]
  wire  _GEN_7732; // @[Execute.scala 117:10]
  wire  _GEN_7733; // @[Execute.scala 117:10]
  wire  _GEN_7734; // @[Execute.scala 117:10]
  wire  _GEN_7735; // @[Execute.scala 117:10]
  wire  _GEN_7736; // @[Execute.scala 117:10]
  wire  _GEN_7737; // @[Execute.scala 117:10]
  wire  _GEN_7738; // @[Execute.scala 117:10]
  wire  _GEN_7739; // @[Execute.scala 117:10]
  wire  _GEN_7740; // @[Execute.scala 117:10]
  wire  _GEN_7741; // @[Execute.scala 117:10]
  wire  _GEN_7742; // @[Execute.scala 117:10]
  wire  _GEN_7743; // @[Execute.scala 117:10]
  wire  _GEN_7744; // @[Execute.scala 117:10]
  wire  _GEN_7745; // @[Execute.scala 117:10]
  wire  _GEN_7747; // @[Execute.scala 117:10]
  wire  _GEN_7748; // @[Execute.scala 117:10]
  wire  _GEN_7749; // @[Execute.scala 117:10]
  wire  _GEN_7750; // @[Execute.scala 117:10]
  wire  _GEN_7751; // @[Execute.scala 117:10]
  wire  _GEN_7752; // @[Execute.scala 117:10]
  wire  _GEN_7753; // @[Execute.scala 117:10]
  wire  _GEN_7754; // @[Execute.scala 117:10]
  wire  _GEN_7755; // @[Execute.scala 117:10]
  wire  _GEN_7756; // @[Execute.scala 117:10]
  wire  _GEN_7757; // @[Execute.scala 117:10]
  wire  _GEN_7758; // @[Execute.scala 117:10]
  wire  _GEN_7759; // @[Execute.scala 117:10]
  wire  _GEN_7760; // @[Execute.scala 117:10]
  wire  _GEN_7761; // @[Execute.scala 117:10]
  wire  _GEN_7762; // @[Execute.scala 117:10]
  wire  _GEN_7763; // @[Execute.scala 117:10]
  wire  _GEN_7764; // @[Execute.scala 117:10]
  wire  _GEN_7765; // @[Execute.scala 117:10]
  wire  _GEN_7766; // @[Execute.scala 117:10]
  wire  _GEN_7767; // @[Execute.scala 117:10]
  wire  _GEN_7768; // @[Execute.scala 117:10]
  wire  _GEN_7769; // @[Execute.scala 117:10]
  wire  _GEN_7770; // @[Execute.scala 117:10]
  wire  _GEN_7771; // @[Execute.scala 117:10]
  wire  _GEN_7772; // @[Execute.scala 117:10]
  wire  _GEN_7773; // @[Execute.scala 117:10]
  wire  _GEN_7774; // @[Execute.scala 117:10]
  wire  _GEN_7775; // @[Execute.scala 117:10]
  wire  _GEN_7776; // @[Execute.scala 117:10]
  wire  _GEN_7777; // @[Execute.scala 117:10]
  wire  _GEN_7778; // @[Execute.scala 117:10]
  wire  _GEN_7779; // @[Execute.scala 117:10]
  wire  _GEN_7780; // @[Execute.scala 117:10]
  wire  _GEN_7781; // @[Execute.scala 117:10]
  wire  _GEN_7782; // @[Execute.scala 117:10]
  wire  _GEN_7783; // @[Execute.scala 117:10]
  wire  _GEN_7784; // @[Execute.scala 117:10]
  wire  _GEN_7785; // @[Execute.scala 117:10]
  wire  _GEN_7786; // @[Execute.scala 117:10]
  wire  _GEN_7787; // @[Execute.scala 117:10]
  wire  _GEN_7788; // @[Execute.scala 117:10]
  wire  _GEN_7789; // @[Execute.scala 117:10]
  wire  _GEN_7790; // @[Execute.scala 117:10]
  wire  _GEN_7791; // @[Execute.scala 117:10]
  wire  _GEN_7792; // @[Execute.scala 117:10]
  wire  _GEN_7793; // @[Execute.scala 117:10]
  wire  _GEN_7794; // @[Execute.scala 117:10]
  wire  _GEN_7795; // @[Execute.scala 117:10]
  wire  _GEN_7796; // @[Execute.scala 117:10]
  wire  _GEN_7797; // @[Execute.scala 117:10]
  wire  _GEN_7798; // @[Execute.scala 117:10]
  wire  _GEN_7799; // @[Execute.scala 117:10]
  wire  _GEN_7800; // @[Execute.scala 117:10]
  wire  _GEN_7801; // @[Execute.scala 117:10]
  wire  _GEN_7802; // @[Execute.scala 117:10]
  wire  _GEN_7803; // @[Execute.scala 117:10]
  wire  _GEN_7804; // @[Execute.scala 117:10]
  wire  _GEN_7805; // @[Execute.scala 117:10]
  wire  _GEN_7806; // @[Execute.scala 117:10]
  wire  _GEN_7807; // @[Execute.scala 117:10]
  wire  _GEN_7808; // @[Execute.scala 117:10]
  wire  _GEN_7809; // @[Execute.scala 117:10]
  wire  _T_691; // @[Execute.scala 117:10]
  wire  _T_692; // @[Execute.scala 117:15]
  wire [5:0] _T_694; // @[Execute.scala 117:37]
  wire [5:0] _T_698; // @[Execute.scala 117:60]
  wire  _GEN_7811; // @[Execute.scala 117:10]
  wire  _GEN_7812; // @[Execute.scala 117:10]
  wire  _GEN_7813; // @[Execute.scala 117:10]
  wire  _GEN_7814; // @[Execute.scala 117:10]
  wire  _GEN_7815; // @[Execute.scala 117:10]
  wire  _GEN_7816; // @[Execute.scala 117:10]
  wire  _GEN_7817; // @[Execute.scala 117:10]
  wire  _GEN_7818; // @[Execute.scala 117:10]
  wire  _GEN_7819; // @[Execute.scala 117:10]
  wire  _GEN_7820; // @[Execute.scala 117:10]
  wire  _GEN_7821; // @[Execute.scala 117:10]
  wire  _GEN_7822; // @[Execute.scala 117:10]
  wire  _GEN_7823; // @[Execute.scala 117:10]
  wire  _GEN_7824; // @[Execute.scala 117:10]
  wire  _GEN_7825; // @[Execute.scala 117:10]
  wire  _GEN_7826; // @[Execute.scala 117:10]
  wire  _GEN_7827; // @[Execute.scala 117:10]
  wire  _GEN_7828; // @[Execute.scala 117:10]
  wire  _GEN_7829; // @[Execute.scala 117:10]
  wire  _GEN_7830; // @[Execute.scala 117:10]
  wire  _GEN_7831; // @[Execute.scala 117:10]
  wire  _GEN_7832; // @[Execute.scala 117:10]
  wire  _GEN_7833; // @[Execute.scala 117:10]
  wire  _GEN_7834; // @[Execute.scala 117:10]
  wire  _GEN_7835; // @[Execute.scala 117:10]
  wire  _GEN_7836; // @[Execute.scala 117:10]
  wire  _GEN_7837; // @[Execute.scala 117:10]
  wire  _GEN_7838; // @[Execute.scala 117:10]
  wire  _GEN_7839; // @[Execute.scala 117:10]
  wire  _GEN_7840; // @[Execute.scala 117:10]
  wire  _GEN_7841; // @[Execute.scala 117:10]
  wire  _GEN_7842; // @[Execute.scala 117:10]
  wire  _GEN_7843; // @[Execute.scala 117:10]
  wire  _GEN_7844; // @[Execute.scala 117:10]
  wire  _GEN_7845; // @[Execute.scala 117:10]
  wire  _GEN_7846; // @[Execute.scala 117:10]
  wire  _GEN_7847; // @[Execute.scala 117:10]
  wire  _GEN_7848; // @[Execute.scala 117:10]
  wire  _GEN_7849; // @[Execute.scala 117:10]
  wire  _GEN_7850; // @[Execute.scala 117:10]
  wire  _GEN_7851; // @[Execute.scala 117:10]
  wire  _GEN_7852; // @[Execute.scala 117:10]
  wire  _GEN_7853; // @[Execute.scala 117:10]
  wire  _GEN_7854; // @[Execute.scala 117:10]
  wire  _GEN_7855; // @[Execute.scala 117:10]
  wire  _GEN_7856; // @[Execute.scala 117:10]
  wire  _GEN_7857; // @[Execute.scala 117:10]
  wire  _GEN_7858; // @[Execute.scala 117:10]
  wire  _GEN_7859; // @[Execute.scala 117:10]
  wire  _GEN_7860; // @[Execute.scala 117:10]
  wire  _GEN_7861; // @[Execute.scala 117:10]
  wire  _GEN_7862; // @[Execute.scala 117:10]
  wire  _GEN_7863; // @[Execute.scala 117:10]
  wire  _GEN_7864; // @[Execute.scala 117:10]
  wire  _GEN_7865; // @[Execute.scala 117:10]
  wire  _GEN_7866; // @[Execute.scala 117:10]
  wire  _GEN_7867; // @[Execute.scala 117:10]
  wire  _GEN_7868; // @[Execute.scala 117:10]
  wire  _GEN_7869; // @[Execute.scala 117:10]
  wire  _GEN_7870; // @[Execute.scala 117:10]
  wire  _GEN_7871; // @[Execute.scala 117:10]
  wire  _GEN_7872; // @[Execute.scala 117:10]
  wire  _GEN_7873; // @[Execute.scala 117:10]
  wire  _GEN_7875; // @[Execute.scala 117:10]
  wire  _GEN_7876; // @[Execute.scala 117:10]
  wire  _GEN_7877; // @[Execute.scala 117:10]
  wire  _GEN_7878; // @[Execute.scala 117:10]
  wire  _GEN_7879; // @[Execute.scala 117:10]
  wire  _GEN_7880; // @[Execute.scala 117:10]
  wire  _GEN_7881; // @[Execute.scala 117:10]
  wire  _GEN_7882; // @[Execute.scala 117:10]
  wire  _GEN_7883; // @[Execute.scala 117:10]
  wire  _GEN_7884; // @[Execute.scala 117:10]
  wire  _GEN_7885; // @[Execute.scala 117:10]
  wire  _GEN_7886; // @[Execute.scala 117:10]
  wire  _GEN_7887; // @[Execute.scala 117:10]
  wire  _GEN_7888; // @[Execute.scala 117:10]
  wire  _GEN_7889; // @[Execute.scala 117:10]
  wire  _GEN_7890; // @[Execute.scala 117:10]
  wire  _GEN_7891; // @[Execute.scala 117:10]
  wire  _GEN_7892; // @[Execute.scala 117:10]
  wire  _GEN_7893; // @[Execute.scala 117:10]
  wire  _GEN_7894; // @[Execute.scala 117:10]
  wire  _GEN_7895; // @[Execute.scala 117:10]
  wire  _GEN_7896; // @[Execute.scala 117:10]
  wire  _GEN_7897; // @[Execute.scala 117:10]
  wire  _GEN_7898; // @[Execute.scala 117:10]
  wire  _GEN_7899; // @[Execute.scala 117:10]
  wire  _GEN_7900; // @[Execute.scala 117:10]
  wire  _GEN_7901; // @[Execute.scala 117:10]
  wire  _GEN_7902; // @[Execute.scala 117:10]
  wire  _GEN_7903; // @[Execute.scala 117:10]
  wire  _GEN_7904; // @[Execute.scala 117:10]
  wire  _GEN_7905; // @[Execute.scala 117:10]
  wire  _GEN_7906; // @[Execute.scala 117:10]
  wire  _GEN_7907; // @[Execute.scala 117:10]
  wire  _GEN_7908; // @[Execute.scala 117:10]
  wire  _GEN_7909; // @[Execute.scala 117:10]
  wire  _GEN_7910; // @[Execute.scala 117:10]
  wire  _GEN_7911; // @[Execute.scala 117:10]
  wire  _GEN_7912; // @[Execute.scala 117:10]
  wire  _GEN_7913; // @[Execute.scala 117:10]
  wire  _GEN_7914; // @[Execute.scala 117:10]
  wire  _GEN_7915; // @[Execute.scala 117:10]
  wire  _GEN_7916; // @[Execute.scala 117:10]
  wire  _GEN_7917; // @[Execute.scala 117:10]
  wire  _GEN_7918; // @[Execute.scala 117:10]
  wire  _GEN_7919; // @[Execute.scala 117:10]
  wire  _GEN_7920; // @[Execute.scala 117:10]
  wire  _GEN_7921; // @[Execute.scala 117:10]
  wire  _GEN_7922; // @[Execute.scala 117:10]
  wire  _GEN_7923; // @[Execute.scala 117:10]
  wire  _GEN_7924; // @[Execute.scala 117:10]
  wire  _GEN_7925; // @[Execute.scala 117:10]
  wire  _GEN_7926; // @[Execute.scala 117:10]
  wire  _GEN_7927; // @[Execute.scala 117:10]
  wire  _GEN_7928; // @[Execute.scala 117:10]
  wire  _GEN_7929; // @[Execute.scala 117:10]
  wire  _GEN_7930; // @[Execute.scala 117:10]
  wire  _GEN_7931; // @[Execute.scala 117:10]
  wire  _GEN_7932; // @[Execute.scala 117:10]
  wire  _GEN_7933; // @[Execute.scala 117:10]
  wire  _GEN_7934; // @[Execute.scala 117:10]
  wire  _GEN_7935; // @[Execute.scala 117:10]
  wire  _GEN_7936; // @[Execute.scala 117:10]
  wire  _GEN_7937; // @[Execute.scala 117:10]
  wire  _T_701; // @[Execute.scala 117:10]
  wire  _T_702; // @[Execute.scala 117:15]
  wire [5:0] _T_704; // @[Execute.scala 117:37]
  wire [5:0] _T_708; // @[Execute.scala 117:60]
  wire  _GEN_7939; // @[Execute.scala 117:10]
  wire  _GEN_7940; // @[Execute.scala 117:10]
  wire  _GEN_7941; // @[Execute.scala 117:10]
  wire  _GEN_7942; // @[Execute.scala 117:10]
  wire  _GEN_7943; // @[Execute.scala 117:10]
  wire  _GEN_7944; // @[Execute.scala 117:10]
  wire  _GEN_7945; // @[Execute.scala 117:10]
  wire  _GEN_7946; // @[Execute.scala 117:10]
  wire  _GEN_7947; // @[Execute.scala 117:10]
  wire  _GEN_7948; // @[Execute.scala 117:10]
  wire  _GEN_7949; // @[Execute.scala 117:10]
  wire  _GEN_7950; // @[Execute.scala 117:10]
  wire  _GEN_7951; // @[Execute.scala 117:10]
  wire  _GEN_7952; // @[Execute.scala 117:10]
  wire  _GEN_7953; // @[Execute.scala 117:10]
  wire  _GEN_7954; // @[Execute.scala 117:10]
  wire  _GEN_7955; // @[Execute.scala 117:10]
  wire  _GEN_7956; // @[Execute.scala 117:10]
  wire  _GEN_7957; // @[Execute.scala 117:10]
  wire  _GEN_7958; // @[Execute.scala 117:10]
  wire  _GEN_7959; // @[Execute.scala 117:10]
  wire  _GEN_7960; // @[Execute.scala 117:10]
  wire  _GEN_7961; // @[Execute.scala 117:10]
  wire  _GEN_7962; // @[Execute.scala 117:10]
  wire  _GEN_7963; // @[Execute.scala 117:10]
  wire  _GEN_7964; // @[Execute.scala 117:10]
  wire  _GEN_7965; // @[Execute.scala 117:10]
  wire  _GEN_7966; // @[Execute.scala 117:10]
  wire  _GEN_7967; // @[Execute.scala 117:10]
  wire  _GEN_7968; // @[Execute.scala 117:10]
  wire  _GEN_7969; // @[Execute.scala 117:10]
  wire  _GEN_7970; // @[Execute.scala 117:10]
  wire  _GEN_7971; // @[Execute.scala 117:10]
  wire  _GEN_7972; // @[Execute.scala 117:10]
  wire  _GEN_7973; // @[Execute.scala 117:10]
  wire  _GEN_7974; // @[Execute.scala 117:10]
  wire  _GEN_7975; // @[Execute.scala 117:10]
  wire  _GEN_7976; // @[Execute.scala 117:10]
  wire  _GEN_7977; // @[Execute.scala 117:10]
  wire  _GEN_7978; // @[Execute.scala 117:10]
  wire  _GEN_7979; // @[Execute.scala 117:10]
  wire  _GEN_7980; // @[Execute.scala 117:10]
  wire  _GEN_7981; // @[Execute.scala 117:10]
  wire  _GEN_7982; // @[Execute.scala 117:10]
  wire  _GEN_7983; // @[Execute.scala 117:10]
  wire  _GEN_7984; // @[Execute.scala 117:10]
  wire  _GEN_7985; // @[Execute.scala 117:10]
  wire  _GEN_7986; // @[Execute.scala 117:10]
  wire  _GEN_7987; // @[Execute.scala 117:10]
  wire  _GEN_7988; // @[Execute.scala 117:10]
  wire  _GEN_7989; // @[Execute.scala 117:10]
  wire  _GEN_7990; // @[Execute.scala 117:10]
  wire  _GEN_7991; // @[Execute.scala 117:10]
  wire  _GEN_7992; // @[Execute.scala 117:10]
  wire  _GEN_7993; // @[Execute.scala 117:10]
  wire  _GEN_7994; // @[Execute.scala 117:10]
  wire  _GEN_7995; // @[Execute.scala 117:10]
  wire  _GEN_7996; // @[Execute.scala 117:10]
  wire  _GEN_7997; // @[Execute.scala 117:10]
  wire  _GEN_7998; // @[Execute.scala 117:10]
  wire  _GEN_7999; // @[Execute.scala 117:10]
  wire  _GEN_8000; // @[Execute.scala 117:10]
  wire  _GEN_8001; // @[Execute.scala 117:10]
  wire  _GEN_8003; // @[Execute.scala 117:10]
  wire  _GEN_8004; // @[Execute.scala 117:10]
  wire  _GEN_8005; // @[Execute.scala 117:10]
  wire  _GEN_8006; // @[Execute.scala 117:10]
  wire  _GEN_8007; // @[Execute.scala 117:10]
  wire  _GEN_8008; // @[Execute.scala 117:10]
  wire  _GEN_8009; // @[Execute.scala 117:10]
  wire  _GEN_8010; // @[Execute.scala 117:10]
  wire  _GEN_8011; // @[Execute.scala 117:10]
  wire  _GEN_8012; // @[Execute.scala 117:10]
  wire  _GEN_8013; // @[Execute.scala 117:10]
  wire  _GEN_8014; // @[Execute.scala 117:10]
  wire  _GEN_8015; // @[Execute.scala 117:10]
  wire  _GEN_8016; // @[Execute.scala 117:10]
  wire  _GEN_8017; // @[Execute.scala 117:10]
  wire  _GEN_8018; // @[Execute.scala 117:10]
  wire  _GEN_8019; // @[Execute.scala 117:10]
  wire  _GEN_8020; // @[Execute.scala 117:10]
  wire  _GEN_8021; // @[Execute.scala 117:10]
  wire  _GEN_8022; // @[Execute.scala 117:10]
  wire  _GEN_8023; // @[Execute.scala 117:10]
  wire  _GEN_8024; // @[Execute.scala 117:10]
  wire  _GEN_8025; // @[Execute.scala 117:10]
  wire  _GEN_8026; // @[Execute.scala 117:10]
  wire  _GEN_8027; // @[Execute.scala 117:10]
  wire  _GEN_8028; // @[Execute.scala 117:10]
  wire  _GEN_8029; // @[Execute.scala 117:10]
  wire  _GEN_8030; // @[Execute.scala 117:10]
  wire  _GEN_8031; // @[Execute.scala 117:10]
  wire  _GEN_8032; // @[Execute.scala 117:10]
  wire  _GEN_8033; // @[Execute.scala 117:10]
  wire  _GEN_8034; // @[Execute.scala 117:10]
  wire  _GEN_8035; // @[Execute.scala 117:10]
  wire  _GEN_8036; // @[Execute.scala 117:10]
  wire  _GEN_8037; // @[Execute.scala 117:10]
  wire  _GEN_8038; // @[Execute.scala 117:10]
  wire  _GEN_8039; // @[Execute.scala 117:10]
  wire  _GEN_8040; // @[Execute.scala 117:10]
  wire  _GEN_8041; // @[Execute.scala 117:10]
  wire  _GEN_8042; // @[Execute.scala 117:10]
  wire  _GEN_8043; // @[Execute.scala 117:10]
  wire  _GEN_8044; // @[Execute.scala 117:10]
  wire  _GEN_8045; // @[Execute.scala 117:10]
  wire  _GEN_8046; // @[Execute.scala 117:10]
  wire  _GEN_8047; // @[Execute.scala 117:10]
  wire  _GEN_8048; // @[Execute.scala 117:10]
  wire  _GEN_8049; // @[Execute.scala 117:10]
  wire  _GEN_8050; // @[Execute.scala 117:10]
  wire  _GEN_8051; // @[Execute.scala 117:10]
  wire  _GEN_8052; // @[Execute.scala 117:10]
  wire  _GEN_8053; // @[Execute.scala 117:10]
  wire  _GEN_8054; // @[Execute.scala 117:10]
  wire  _GEN_8055; // @[Execute.scala 117:10]
  wire  _GEN_8056; // @[Execute.scala 117:10]
  wire  _GEN_8057; // @[Execute.scala 117:10]
  wire  _GEN_8058; // @[Execute.scala 117:10]
  wire  _GEN_8059; // @[Execute.scala 117:10]
  wire  _GEN_8060; // @[Execute.scala 117:10]
  wire  _GEN_8061; // @[Execute.scala 117:10]
  wire  _GEN_8062; // @[Execute.scala 117:10]
  wire  _GEN_8063; // @[Execute.scala 117:10]
  wire  _GEN_8064; // @[Execute.scala 117:10]
  wire  _GEN_8065; // @[Execute.scala 117:10]
  wire  _T_711; // @[Execute.scala 117:10]
  wire  _T_712; // @[Execute.scala 117:15]
  wire [5:0] _T_714; // @[Execute.scala 117:37]
  wire [5:0] _T_718; // @[Execute.scala 117:60]
  wire  _GEN_8067; // @[Execute.scala 117:10]
  wire  _GEN_8068; // @[Execute.scala 117:10]
  wire  _GEN_8069; // @[Execute.scala 117:10]
  wire  _GEN_8070; // @[Execute.scala 117:10]
  wire  _GEN_8071; // @[Execute.scala 117:10]
  wire  _GEN_8072; // @[Execute.scala 117:10]
  wire  _GEN_8073; // @[Execute.scala 117:10]
  wire  _GEN_8074; // @[Execute.scala 117:10]
  wire  _GEN_8075; // @[Execute.scala 117:10]
  wire  _GEN_8076; // @[Execute.scala 117:10]
  wire  _GEN_8077; // @[Execute.scala 117:10]
  wire  _GEN_8078; // @[Execute.scala 117:10]
  wire  _GEN_8079; // @[Execute.scala 117:10]
  wire  _GEN_8080; // @[Execute.scala 117:10]
  wire  _GEN_8081; // @[Execute.scala 117:10]
  wire  _GEN_8082; // @[Execute.scala 117:10]
  wire  _GEN_8083; // @[Execute.scala 117:10]
  wire  _GEN_8084; // @[Execute.scala 117:10]
  wire  _GEN_8085; // @[Execute.scala 117:10]
  wire  _GEN_8086; // @[Execute.scala 117:10]
  wire  _GEN_8087; // @[Execute.scala 117:10]
  wire  _GEN_8088; // @[Execute.scala 117:10]
  wire  _GEN_8089; // @[Execute.scala 117:10]
  wire  _GEN_8090; // @[Execute.scala 117:10]
  wire  _GEN_8091; // @[Execute.scala 117:10]
  wire  _GEN_8092; // @[Execute.scala 117:10]
  wire  _GEN_8093; // @[Execute.scala 117:10]
  wire  _GEN_8094; // @[Execute.scala 117:10]
  wire  _GEN_8095; // @[Execute.scala 117:10]
  wire  _GEN_8096; // @[Execute.scala 117:10]
  wire  _GEN_8097; // @[Execute.scala 117:10]
  wire  _GEN_8098; // @[Execute.scala 117:10]
  wire  _GEN_8099; // @[Execute.scala 117:10]
  wire  _GEN_8100; // @[Execute.scala 117:10]
  wire  _GEN_8101; // @[Execute.scala 117:10]
  wire  _GEN_8102; // @[Execute.scala 117:10]
  wire  _GEN_8103; // @[Execute.scala 117:10]
  wire  _GEN_8104; // @[Execute.scala 117:10]
  wire  _GEN_8105; // @[Execute.scala 117:10]
  wire  _GEN_8106; // @[Execute.scala 117:10]
  wire  _GEN_8107; // @[Execute.scala 117:10]
  wire  _GEN_8108; // @[Execute.scala 117:10]
  wire  _GEN_8109; // @[Execute.scala 117:10]
  wire  _GEN_8110; // @[Execute.scala 117:10]
  wire  _GEN_8111; // @[Execute.scala 117:10]
  wire  _GEN_8112; // @[Execute.scala 117:10]
  wire  _GEN_8113; // @[Execute.scala 117:10]
  wire  _GEN_8114; // @[Execute.scala 117:10]
  wire  _GEN_8115; // @[Execute.scala 117:10]
  wire  _GEN_8116; // @[Execute.scala 117:10]
  wire  _GEN_8117; // @[Execute.scala 117:10]
  wire  _GEN_8118; // @[Execute.scala 117:10]
  wire  _GEN_8119; // @[Execute.scala 117:10]
  wire  _GEN_8120; // @[Execute.scala 117:10]
  wire  _GEN_8121; // @[Execute.scala 117:10]
  wire  _GEN_8122; // @[Execute.scala 117:10]
  wire  _GEN_8123; // @[Execute.scala 117:10]
  wire  _GEN_8124; // @[Execute.scala 117:10]
  wire  _GEN_8125; // @[Execute.scala 117:10]
  wire  _GEN_8126; // @[Execute.scala 117:10]
  wire  _GEN_8127; // @[Execute.scala 117:10]
  wire  _GEN_8128; // @[Execute.scala 117:10]
  wire  _GEN_8129; // @[Execute.scala 117:10]
  wire  _GEN_8131; // @[Execute.scala 117:10]
  wire  _GEN_8132; // @[Execute.scala 117:10]
  wire  _GEN_8133; // @[Execute.scala 117:10]
  wire  _GEN_8134; // @[Execute.scala 117:10]
  wire  _GEN_8135; // @[Execute.scala 117:10]
  wire  _GEN_8136; // @[Execute.scala 117:10]
  wire  _GEN_8137; // @[Execute.scala 117:10]
  wire  _GEN_8138; // @[Execute.scala 117:10]
  wire  _GEN_8139; // @[Execute.scala 117:10]
  wire  _GEN_8140; // @[Execute.scala 117:10]
  wire  _GEN_8141; // @[Execute.scala 117:10]
  wire  _GEN_8142; // @[Execute.scala 117:10]
  wire  _GEN_8143; // @[Execute.scala 117:10]
  wire  _GEN_8144; // @[Execute.scala 117:10]
  wire  _GEN_8145; // @[Execute.scala 117:10]
  wire  _GEN_8146; // @[Execute.scala 117:10]
  wire  _GEN_8147; // @[Execute.scala 117:10]
  wire  _GEN_8148; // @[Execute.scala 117:10]
  wire  _GEN_8149; // @[Execute.scala 117:10]
  wire  _GEN_8150; // @[Execute.scala 117:10]
  wire  _GEN_8151; // @[Execute.scala 117:10]
  wire  _GEN_8152; // @[Execute.scala 117:10]
  wire  _GEN_8153; // @[Execute.scala 117:10]
  wire  _GEN_8154; // @[Execute.scala 117:10]
  wire  _GEN_8155; // @[Execute.scala 117:10]
  wire  _GEN_8156; // @[Execute.scala 117:10]
  wire  _GEN_8157; // @[Execute.scala 117:10]
  wire  _GEN_8158; // @[Execute.scala 117:10]
  wire  _GEN_8159; // @[Execute.scala 117:10]
  wire  _GEN_8160; // @[Execute.scala 117:10]
  wire  _GEN_8161; // @[Execute.scala 117:10]
  wire  _GEN_8162; // @[Execute.scala 117:10]
  wire  _GEN_8163; // @[Execute.scala 117:10]
  wire  _GEN_8164; // @[Execute.scala 117:10]
  wire  _GEN_8165; // @[Execute.scala 117:10]
  wire  _GEN_8166; // @[Execute.scala 117:10]
  wire  _GEN_8167; // @[Execute.scala 117:10]
  wire  _GEN_8168; // @[Execute.scala 117:10]
  wire  _GEN_8169; // @[Execute.scala 117:10]
  wire  _GEN_8170; // @[Execute.scala 117:10]
  wire  _GEN_8171; // @[Execute.scala 117:10]
  wire  _GEN_8172; // @[Execute.scala 117:10]
  wire  _GEN_8173; // @[Execute.scala 117:10]
  wire  _GEN_8174; // @[Execute.scala 117:10]
  wire  _GEN_8175; // @[Execute.scala 117:10]
  wire  _GEN_8176; // @[Execute.scala 117:10]
  wire  _GEN_8177; // @[Execute.scala 117:10]
  wire  _GEN_8178; // @[Execute.scala 117:10]
  wire  _GEN_8179; // @[Execute.scala 117:10]
  wire  _GEN_8180; // @[Execute.scala 117:10]
  wire  _GEN_8181; // @[Execute.scala 117:10]
  wire  _GEN_8182; // @[Execute.scala 117:10]
  wire  _GEN_8183; // @[Execute.scala 117:10]
  wire  _GEN_8184; // @[Execute.scala 117:10]
  wire  _GEN_8185; // @[Execute.scala 117:10]
  wire  _GEN_8186; // @[Execute.scala 117:10]
  wire  _GEN_8187; // @[Execute.scala 117:10]
  wire  _GEN_8188; // @[Execute.scala 117:10]
  wire  _GEN_8189; // @[Execute.scala 117:10]
  wire  _GEN_8190; // @[Execute.scala 117:10]
  wire  _GEN_8191; // @[Execute.scala 117:10]
  wire  _GEN_8192; // @[Execute.scala 117:10]
  wire  _GEN_8193; // @[Execute.scala 117:10]
  wire  _T_721; // @[Execute.scala 117:10]
  wire  _T_722; // @[Execute.scala 117:15]
  wire [5:0] _T_724; // @[Execute.scala 117:37]
  wire [5:0] _T_728; // @[Execute.scala 117:60]
  wire  _GEN_8195; // @[Execute.scala 117:10]
  wire  _GEN_8196; // @[Execute.scala 117:10]
  wire  _GEN_8197; // @[Execute.scala 117:10]
  wire  _GEN_8198; // @[Execute.scala 117:10]
  wire  _GEN_8199; // @[Execute.scala 117:10]
  wire  _GEN_8200; // @[Execute.scala 117:10]
  wire  _GEN_8201; // @[Execute.scala 117:10]
  wire  _GEN_8202; // @[Execute.scala 117:10]
  wire  _GEN_8203; // @[Execute.scala 117:10]
  wire  _GEN_8204; // @[Execute.scala 117:10]
  wire  _GEN_8205; // @[Execute.scala 117:10]
  wire  _GEN_8206; // @[Execute.scala 117:10]
  wire  _GEN_8207; // @[Execute.scala 117:10]
  wire  _GEN_8208; // @[Execute.scala 117:10]
  wire  _GEN_8209; // @[Execute.scala 117:10]
  wire  _GEN_8210; // @[Execute.scala 117:10]
  wire  _GEN_8211; // @[Execute.scala 117:10]
  wire  _GEN_8212; // @[Execute.scala 117:10]
  wire  _GEN_8213; // @[Execute.scala 117:10]
  wire  _GEN_8214; // @[Execute.scala 117:10]
  wire  _GEN_8215; // @[Execute.scala 117:10]
  wire  _GEN_8216; // @[Execute.scala 117:10]
  wire  _GEN_8217; // @[Execute.scala 117:10]
  wire  _GEN_8218; // @[Execute.scala 117:10]
  wire  _GEN_8219; // @[Execute.scala 117:10]
  wire  _GEN_8220; // @[Execute.scala 117:10]
  wire  _GEN_8221; // @[Execute.scala 117:10]
  wire  _GEN_8222; // @[Execute.scala 117:10]
  wire  _GEN_8223; // @[Execute.scala 117:10]
  wire  _GEN_8224; // @[Execute.scala 117:10]
  wire  _GEN_8225; // @[Execute.scala 117:10]
  wire  _GEN_8226; // @[Execute.scala 117:10]
  wire  _GEN_8227; // @[Execute.scala 117:10]
  wire  _GEN_8228; // @[Execute.scala 117:10]
  wire  _GEN_8229; // @[Execute.scala 117:10]
  wire  _GEN_8230; // @[Execute.scala 117:10]
  wire  _GEN_8231; // @[Execute.scala 117:10]
  wire  _GEN_8232; // @[Execute.scala 117:10]
  wire  _GEN_8233; // @[Execute.scala 117:10]
  wire  _GEN_8234; // @[Execute.scala 117:10]
  wire  _GEN_8235; // @[Execute.scala 117:10]
  wire  _GEN_8236; // @[Execute.scala 117:10]
  wire  _GEN_8237; // @[Execute.scala 117:10]
  wire  _GEN_8238; // @[Execute.scala 117:10]
  wire  _GEN_8239; // @[Execute.scala 117:10]
  wire  _GEN_8240; // @[Execute.scala 117:10]
  wire  _GEN_8241; // @[Execute.scala 117:10]
  wire  _GEN_8242; // @[Execute.scala 117:10]
  wire  _GEN_8243; // @[Execute.scala 117:10]
  wire  _GEN_8244; // @[Execute.scala 117:10]
  wire  _GEN_8245; // @[Execute.scala 117:10]
  wire  _GEN_8246; // @[Execute.scala 117:10]
  wire  _GEN_8247; // @[Execute.scala 117:10]
  wire  _GEN_8248; // @[Execute.scala 117:10]
  wire  _GEN_8249; // @[Execute.scala 117:10]
  wire  _GEN_8250; // @[Execute.scala 117:10]
  wire  _GEN_8251; // @[Execute.scala 117:10]
  wire  _GEN_8252; // @[Execute.scala 117:10]
  wire  _GEN_8253; // @[Execute.scala 117:10]
  wire  _GEN_8254; // @[Execute.scala 117:10]
  wire  _GEN_8255; // @[Execute.scala 117:10]
  wire  _GEN_8256; // @[Execute.scala 117:10]
  wire  _GEN_8257; // @[Execute.scala 117:10]
  wire  _GEN_8259; // @[Execute.scala 117:10]
  wire  _GEN_8260; // @[Execute.scala 117:10]
  wire  _GEN_8261; // @[Execute.scala 117:10]
  wire  _GEN_8262; // @[Execute.scala 117:10]
  wire  _GEN_8263; // @[Execute.scala 117:10]
  wire  _GEN_8264; // @[Execute.scala 117:10]
  wire  _GEN_8265; // @[Execute.scala 117:10]
  wire  _GEN_8266; // @[Execute.scala 117:10]
  wire  _GEN_8267; // @[Execute.scala 117:10]
  wire  _GEN_8268; // @[Execute.scala 117:10]
  wire  _GEN_8269; // @[Execute.scala 117:10]
  wire  _GEN_8270; // @[Execute.scala 117:10]
  wire  _GEN_8271; // @[Execute.scala 117:10]
  wire  _GEN_8272; // @[Execute.scala 117:10]
  wire  _GEN_8273; // @[Execute.scala 117:10]
  wire  _GEN_8274; // @[Execute.scala 117:10]
  wire  _GEN_8275; // @[Execute.scala 117:10]
  wire  _GEN_8276; // @[Execute.scala 117:10]
  wire  _GEN_8277; // @[Execute.scala 117:10]
  wire  _GEN_8278; // @[Execute.scala 117:10]
  wire  _GEN_8279; // @[Execute.scala 117:10]
  wire  _GEN_8280; // @[Execute.scala 117:10]
  wire  _GEN_8281; // @[Execute.scala 117:10]
  wire  _GEN_8282; // @[Execute.scala 117:10]
  wire  _GEN_8283; // @[Execute.scala 117:10]
  wire  _GEN_8284; // @[Execute.scala 117:10]
  wire  _GEN_8285; // @[Execute.scala 117:10]
  wire  _GEN_8286; // @[Execute.scala 117:10]
  wire  _GEN_8287; // @[Execute.scala 117:10]
  wire  _GEN_8288; // @[Execute.scala 117:10]
  wire  _GEN_8289; // @[Execute.scala 117:10]
  wire  _GEN_8290; // @[Execute.scala 117:10]
  wire  _GEN_8291; // @[Execute.scala 117:10]
  wire  _GEN_8292; // @[Execute.scala 117:10]
  wire  _GEN_8293; // @[Execute.scala 117:10]
  wire  _GEN_8294; // @[Execute.scala 117:10]
  wire  _GEN_8295; // @[Execute.scala 117:10]
  wire  _GEN_8296; // @[Execute.scala 117:10]
  wire  _GEN_8297; // @[Execute.scala 117:10]
  wire  _GEN_8298; // @[Execute.scala 117:10]
  wire  _GEN_8299; // @[Execute.scala 117:10]
  wire  _GEN_8300; // @[Execute.scala 117:10]
  wire  _GEN_8301; // @[Execute.scala 117:10]
  wire  _GEN_8302; // @[Execute.scala 117:10]
  wire  _GEN_8303; // @[Execute.scala 117:10]
  wire  _GEN_8304; // @[Execute.scala 117:10]
  wire  _GEN_8305; // @[Execute.scala 117:10]
  wire  _GEN_8306; // @[Execute.scala 117:10]
  wire  _GEN_8307; // @[Execute.scala 117:10]
  wire  _GEN_8308; // @[Execute.scala 117:10]
  wire  _GEN_8309; // @[Execute.scala 117:10]
  wire  _GEN_8310; // @[Execute.scala 117:10]
  wire  _GEN_8311; // @[Execute.scala 117:10]
  wire  _GEN_8312; // @[Execute.scala 117:10]
  wire  _GEN_8313; // @[Execute.scala 117:10]
  wire  _GEN_8314; // @[Execute.scala 117:10]
  wire  _GEN_8315; // @[Execute.scala 117:10]
  wire  _GEN_8316; // @[Execute.scala 117:10]
  wire  _GEN_8317; // @[Execute.scala 117:10]
  wire  _GEN_8318; // @[Execute.scala 117:10]
  wire  _GEN_8319; // @[Execute.scala 117:10]
  wire  _GEN_8320; // @[Execute.scala 117:10]
  wire  _GEN_8321; // @[Execute.scala 117:10]
  wire  _T_731; // @[Execute.scala 117:10]
  wire [7:0] _T_739; // @[Execute.scala 302:55]
  wire [15:0] _T_747; // @[Execute.scala 302:55]
  wire [7:0] _T_754; // @[Execute.scala 302:55]
  wire [31:0] _T_763; // @[Execute.scala 302:55]
  wire [7:0] _T_770; // @[Execute.scala 302:55]
  wire [15:0] _T_778; // @[Execute.scala 302:55]
  wire [7:0] _T_785; // @[Execute.scala 302:55]
  wire [31:0] _T_794; // @[Execute.scala 302:55]
  wire [63:0] _T_795; // @[Execute.scala 302:55]
  wire [63:0] _GEN_8323; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8324; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8325; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8326; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8327; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8328; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8329; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8330; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8331; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8332; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8333; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8334; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8335; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8336; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8337; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8338; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8339; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8340; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8341; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8342; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8343; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8344; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8345; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8346; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8347; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8348; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8349; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8350; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8351; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8352; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8353; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8354; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8355; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8356; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8357; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8358; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8359; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8360; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8361; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8362; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8363; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8364; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8365; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8366; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8367; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8368; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8369; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8370; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8371; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8372; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8373; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8374; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8375; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8376; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8377; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8378; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8379; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8380; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8381; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8382; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8383; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8384; // @[Execute.scala 304:9]
  wire [63:0] _GEN_8385; // @[Execute.scala 304:9]
  wire [5:0] _GEN_10438; // @[Execute.scala 117:37]
  wire [5:0] _T_835; // @[Execute.scala 117:37]
  wire  _GEN_8388; // @[Execute.scala 117:10]
  wire  _GEN_8389; // @[Execute.scala 117:10]
  wire  _GEN_8390; // @[Execute.scala 117:10]
  wire  _GEN_8391; // @[Execute.scala 117:10]
  wire  _GEN_8392; // @[Execute.scala 117:10]
  wire  _GEN_8393; // @[Execute.scala 117:10]
  wire  _GEN_8394; // @[Execute.scala 117:10]
  wire  _GEN_8395; // @[Execute.scala 117:10]
  wire  _GEN_8396; // @[Execute.scala 117:10]
  wire  _GEN_8397; // @[Execute.scala 117:10]
  wire  _GEN_8398; // @[Execute.scala 117:10]
  wire  _GEN_8399; // @[Execute.scala 117:10]
  wire  _GEN_8400; // @[Execute.scala 117:10]
  wire  _GEN_8401; // @[Execute.scala 117:10]
  wire  _GEN_8402; // @[Execute.scala 117:10]
  wire  _GEN_8403; // @[Execute.scala 117:10]
  wire  _GEN_8404; // @[Execute.scala 117:10]
  wire  _GEN_8405; // @[Execute.scala 117:10]
  wire  _GEN_8406; // @[Execute.scala 117:10]
  wire  _GEN_8407; // @[Execute.scala 117:10]
  wire  _GEN_8408; // @[Execute.scala 117:10]
  wire  _GEN_8409; // @[Execute.scala 117:10]
  wire  _GEN_8410; // @[Execute.scala 117:10]
  wire  _GEN_8411; // @[Execute.scala 117:10]
  wire  _GEN_8412; // @[Execute.scala 117:10]
  wire  _GEN_8413; // @[Execute.scala 117:10]
  wire  _GEN_8414; // @[Execute.scala 117:10]
  wire  _GEN_8415; // @[Execute.scala 117:10]
  wire  _GEN_8416; // @[Execute.scala 117:10]
  wire  _GEN_8417; // @[Execute.scala 117:10]
  wire  _GEN_8418; // @[Execute.scala 117:10]
  wire  _T_840; // @[Execute.scala 117:15]
  wire [4:0] _T_842; // @[Execute.scala 117:37]
  wire [4:0] _T_844; // @[Execute.scala 117:60]
  wire  _GEN_8452; // @[Execute.scala 117:10]
  wire  _GEN_8453; // @[Execute.scala 117:10]
  wire  _GEN_8454; // @[Execute.scala 117:10]
  wire  _GEN_8455; // @[Execute.scala 117:10]
  wire  _GEN_8456; // @[Execute.scala 117:10]
  wire  _GEN_8457; // @[Execute.scala 117:10]
  wire  _GEN_8458; // @[Execute.scala 117:10]
  wire  _GEN_8459; // @[Execute.scala 117:10]
  wire  _GEN_8460; // @[Execute.scala 117:10]
  wire  _GEN_8461; // @[Execute.scala 117:10]
  wire  _GEN_8462; // @[Execute.scala 117:10]
  wire  _GEN_8463; // @[Execute.scala 117:10]
  wire  _GEN_8464; // @[Execute.scala 117:10]
  wire  _GEN_8465; // @[Execute.scala 117:10]
  wire  _GEN_8466; // @[Execute.scala 117:10]
  wire  _GEN_8467; // @[Execute.scala 117:10]
  wire  _GEN_8468; // @[Execute.scala 117:10]
  wire  _GEN_8469; // @[Execute.scala 117:10]
  wire  _GEN_8470; // @[Execute.scala 117:10]
  wire  _GEN_8471; // @[Execute.scala 117:10]
  wire  _GEN_8472; // @[Execute.scala 117:10]
  wire  _GEN_8473; // @[Execute.scala 117:10]
  wire  _GEN_8474; // @[Execute.scala 117:10]
  wire  _GEN_8475; // @[Execute.scala 117:10]
  wire  _GEN_8476; // @[Execute.scala 117:10]
  wire  _GEN_8477; // @[Execute.scala 117:10]
  wire  _GEN_8478; // @[Execute.scala 117:10]
  wire  _GEN_8479; // @[Execute.scala 117:10]
  wire  _GEN_8480; // @[Execute.scala 117:10]
  wire  _GEN_8481; // @[Execute.scala 117:10]
  wire  _GEN_8482; // @[Execute.scala 117:10]
  wire  _GEN_8484; // @[Execute.scala 117:10]
  wire  _GEN_8485; // @[Execute.scala 117:10]
  wire  _GEN_8486; // @[Execute.scala 117:10]
  wire  _GEN_8487; // @[Execute.scala 117:10]
  wire  _GEN_8488; // @[Execute.scala 117:10]
  wire  _GEN_8489; // @[Execute.scala 117:10]
  wire  _GEN_8490; // @[Execute.scala 117:10]
  wire  _GEN_8491; // @[Execute.scala 117:10]
  wire  _GEN_8492; // @[Execute.scala 117:10]
  wire  _GEN_8493; // @[Execute.scala 117:10]
  wire  _GEN_8494; // @[Execute.scala 117:10]
  wire  _GEN_8495; // @[Execute.scala 117:10]
  wire  _GEN_8496; // @[Execute.scala 117:10]
  wire  _GEN_8497; // @[Execute.scala 117:10]
  wire  _GEN_8498; // @[Execute.scala 117:10]
  wire  _GEN_8499; // @[Execute.scala 117:10]
  wire  _GEN_8500; // @[Execute.scala 117:10]
  wire  _GEN_8501; // @[Execute.scala 117:10]
  wire  _GEN_8502; // @[Execute.scala 117:10]
  wire  _GEN_8503; // @[Execute.scala 117:10]
  wire  _GEN_8504; // @[Execute.scala 117:10]
  wire  _GEN_8505; // @[Execute.scala 117:10]
  wire  _GEN_8506; // @[Execute.scala 117:10]
  wire  _GEN_8507; // @[Execute.scala 117:10]
  wire  _GEN_8508; // @[Execute.scala 117:10]
  wire  _GEN_8509; // @[Execute.scala 117:10]
  wire  _GEN_8510; // @[Execute.scala 117:10]
  wire  _GEN_8511; // @[Execute.scala 117:10]
  wire  _GEN_8512; // @[Execute.scala 117:10]
  wire  _GEN_8513; // @[Execute.scala 117:10]
  wire  _GEN_8514; // @[Execute.scala 117:10]
  wire  _T_845; // @[Execute.scala 117:10]
  wire  _T_846; // @[Execute.scala 117:15]
  wire [4:0] _T_848; // @[Execute.scala 117:37]
  wire [4:0] _T_850; // @[Execute.scala 117:60]
  wire  _GEN_8516; // @[Execute.scala 117:10]
  wire  _GEN_8517; // @[Execute.scala 117:10]
  wire  _GEN_8518; // @[Execute.scala 117:10]
  wire  _GEN_8519; // @[Execute.scala 117:10]
  wire  _GEN_8520; // @[Execute.scala 117:10]
  wire  _GEN_8521; // @[Execute.scala 117:10]
  wire  _GEN_8522; // @[Execute.scala 117:10]
  wire  _GEN_8523; // @[Execute.scala 117:10]
  wire  _GEN_8524; // @[Execute.scala 117:10]
  wire  _GEN_8525; // @[Execute.scala 117:10]
  wire  _GEN_8526; // @[Execute.scala 117:10]
  wire  _GEN_8527; // @[Execute.scala 117:10]
  wire  _GEN_8528; // @[Execute.scala 117:10]
  wire  _GEN_8529; // @[Execute.scala 117:10]
  wire  _GEN_8530; // @[Execute.scala 117:10]
  wire  _GEN_8531; // @[Execute.scala 117:10]
  wire  _GEN_8532; // @[Execute.scala 117:10]
  wire  _GEN_8533; // @[Execute.scala 117:10]
  wire  _GEN_8534; // @[Execute.scala 117:10]
  wire  _GEN_8535; // @[Execute.scala 117:10]
  wire  _GEN_8536; // @[Execute.scala 117:10]
  wire  _GEN_8537; // @[Execute.scala 117:10]
  wire  _GEN_8538; // @[Execute.scala 117:10]
  wire  _GEN_8539; // @[Execute.scala 117:10]
  wire  _GEN_8540; // @[Execute.scala 117:10]
  wire  _GEN_8541; // @[Execute.scala 117:10]
  wire  _GEN_8542; // @[Execute.scala 117:10]
  wire  _GEN_8543; // @[Execute.scala 117:10]
  wire  _GEN_8544; // @[Execute.scala 117:10]
  wire  _GEN_8545; // @[Execute.scala 117:10]
  wire  _GEN_8546; // @[Execute.scala 117:10]
  wire  _GEN_8548; // @[Execute.scala 117:10]
  wire  _GEN_8549; // @[Execute.scala 117:10]
  wire  _GEN_8550; // @[Execute.scala 117:10]
  wire  _GEN_8551; // @[Execute.scala 117:10]
  wire  _GEN_8552; // @[Execute.scala 117:10]
  wire  _GEN_8553; // @[Execute.scala 117:10]
  wire  _GEN_8554; // @[Execute.scala 117:10]
  wire  _GEN_8555; // @[Execute.scala 117:10]
  wire  _GEN_8556; // @[Execute.scala 117:10]
  wire  _GEN_8557; // @[Execute.scala 117:10]
  wire  _GEN_8558; // @[Execute.scala 117:10]
  wire  _GEN_8559; // @[Execute.scala 117:10]
  wire  _GEN_8560; // @[Execute.scala 117:10]
  wire  _GEN_8561; // @[Execute.scala 117:10]
  wire  _GEN_8562; // @[Execute.scala 117:10]
  wire  _GEN_8563; // @[Execute.scala 117:10]
  wire  _GEN_8564; // @[Execute.scala 117:10]
  wire  _GEN_8565; // @[Execute.scala 117:10]
  wire  _GEN_8566; // @[Execute.scala 117:10]
  wire  _GEN_8567; // @[Execute.scala 117:10]
  wire  _GEN_8568; // @[Execute.scala 117:10]
  wire  _GEN_8569; // @[Execute.scala 117:10]
  wire  _GEN_8570; // @[Execute.scala 117:10]
  wire  _GEN_8571; // @[Execute.scala 117:10]
  wire  _GEN_8572; // @[Execute.scala 117:10]
  wire  _GEN_8573; // @[Execute.scala 117:10]
  wire  _GEN_8574; // @[Execute.scala 117:10]
  wire  _GEN_8575; // @[Execute.scala 117:10]
  wire  _GEN_8576; // @[Execute.scala 117:10]
  wire  _GEN_8577; // @[Execute.scala 117:10]
  wire  _GEN_8578; // @[Execute.scala 117:10]
  wire  _T_851; // @[Execute.scala 117:10]
  wire  _T_852; // @[Execute.scala 117:15]
  wire [4:0] _T_854; // @[Execute.scala 117:37]
  wire [4:0] _T_856; // @[Execute.scala 117:60]
  wire  _GEN_8580; // @[Execute.scala 117:10]
  wire  _GEN_8581; // @[Execute.scala 117:10]
  wire  _GEN_8582; // @[Execute.scala 117:10]
  wire  _GEN_8583; // @[Execute.scala 117:10]
  wire  _GEN_8584; // @[Execute.scala 117:10]
  wire  _GEN_8585; // @[Execute.scala 117:10]
  wire  _GEN_8586; // @[Execute.scala 117:10]
  wire  _GEN_8587; // @[Execute.scala 117:10]
  wire  _GEN_8588; // @[Execute.scala 117:10]
  wire  _GEN_8589; // @[Execute.scala 117:10]
  wire  _GEN_8590; // @[Execute.scala 117:10]
  wire  _GEN_8591; // @[Execute.scala 117:10]
  wire  _GEN_8592; // @[Execute.scala 117:10]
  wire  _GEN_8593; // @[Execute.scala 117:10]
  wire  _GEN_8594; // @[Execute.scala 117:10]
  wire  _GEN_8595; // @[Execute.scala 117:10]
  wire  _GEN_8596; // @[Execute.scala 117:10]
  wire  _GEN_8597; // @[Execute.scala 117:10]
  wire  _GEN_8598; // @[Execute.scala 117:10]
  wire  _GEN_8599; // @[Execute.scala 117:10]
  wire  _GEN_8600; // @[Execute.scala 117:10]
  wire  _GEN_8601; // @[Execute.scala 117:10]
  wire  _GEN_8602; // @[Execute.scala 117:10]
  wire  _GEN_8603; // @[Execute.scala 117:10]
  wire  _GEN_8604; // @[Execute.scala 117:10]
  wire  _GEN_8605; // @[Execute.scala 117:10]
  wire  _GEN_8606; // @[Execute.scala 117:10]
  wire  _GEN_8607; // @[Execute.scala 117:10]
  wire  _GEN_8608; // @[Execute.scala 117:10]
  wire  _GEN_8609; // @[Execute.scala 117:10]
  wire  _GEN_8610; // @[Execute.scala 117:10]
  wire  _GEN_8612; // @[Execute.scala 117:10]
  wire  _GEN_8613; // @[Execute.scala 117:10]
  wire  _GEN_8614; // @[Execute.scala 117:10]
  wire  _GEN_8615; // @[Execute.scala 117:10]
  wire  _GEN_8616; // @[Execute.scala 117:10]
  wire  _GEN_8617; // @[Execute.scala 117:10]
  wire  _GEN_8618; // @[Execute.scala 117:10]
  wire  _GEN_8619; // @[Execute.scala 117:10]
  wire  _GEN_8620; // @[Execute.scala 117:10]
  wire  _GEN_8621; // @[Execute.scala 117:10]
  wire  _GEN_8622; // @[Execute.scala 117:10]
  wire  _GEN_8623; // @[Execute.scala 117:10]
  wire  _GEN_8624; // @[Execute.scala 117:10]
  wire  _GEN_8625; // @[Execute.scala 117:10]
  wire  _GEN_8626; // @[Execute.scala 117:10]
  wire  _GEN_8627; // @[Execute.scala 117:10]
  wire  _GEN_8628; // @[Execute.scala 117:10]
  wire  _GEN_8629; // @[Execute.scala 117:10]
  wire  _GEN_8630; // @[Execute.scala 117:10]
  wire  _GEN_8631; // @[Execute.scala 117:10]
  wire  _GEN_8632; // @[Execute.scala 117:10]
  wire  _GEN_8633; // @[Execute.scala 117:10]
  wire  _GEN_8634; // @[Execute.scala 117:10]
  wire  _GEN_8635; // @[Execute.scala 117:10]
  wire  _GEN_8636; // @[Execute.scala 117:10]
  wire  _GEN_8637; // @[Execute.scala 117:10]
  wire  _GEN_8638; // @[Execute.scala 117:10]
  wire  _GEN_8639; // @[Execute.scala 117:10]
  wire  _GEN_8640; // @[Execute.scala 117:10]
  wire  _GEN_8641; // @[Execute.scala 117:10]
  wire  _GEN_8642; // @[Execute.scala 117:10]
  wire  _T_857; // @[Execute.scala 117:10]
  wire  _T_858; // @[Execute.scala 117:15]
  wire [4:0] _T_860; // @[Execute.scala 117:37]
  wire [4:0] _T_862; // @[Execute.scala 117:60]
  wire  _GEN_8644; // @[Execute.scala 117:10]
  wire  _GEN_8645; // @[Execute.scala 117:10]
  wire  _GEN_8646; // @[Execute.scala 117:10]
  wire  _GEN_8647; // @[Execute.scala 117:10]
  wire  _GEN_8648; // @[Execute.scala 117:10]
  wire  _GEN_8649; // @[Execute.scala 117:10]
  wire  _GEN_8650; // @[Execute.scala 117:10]
  wire  _GEN_8651; // @[Execute.scala 117:10]
  wire  _GEN_8652; // @[Execute.scala 117:10]
  wire  _GEN_8653; // @[Execute.scala 117:10]
  wire  _GEN_8654; // @[Execute.scala 117:10]
  wire  _GEN_8655; // @[Execute.scala 117:10]
  wire  _GEN_8656; // @[Execute.scala 117:10]
  wire  _GEN_8657; // @[Execute.scala 117:10]
  wire  _GEN_8658; // @[Execute.scala 117:10]
  wire  _GEN_8659; // @[Execute.scala 117:10]
  wire  _GEN_8660; // @[Execute.scala 117:10]
  wire  _GEN_8661; // @[Execute.scala 117:10]
  wire  _GEN_8662; // @[Execute.scala 117:10]
  wire  _GEN_8663; // @[Execute.scala 117:10]
  wire  _GEN_8664; // @[Execute.scala 117:10]
  wire  _GEN_8665; // @[Execute.scala 117:10]
  wire  _GEN_8666; // @[Execute.scala 117:10]
  wire  _GEN_8667; // @[Execute.scala 117:10]
  wire  _GEN_8668; // @[Execute.scala 117:10]
  wire  _GEN_8669; // @[Execute.scala 117:10]
  wire  _GEN_8670; // @[Execute.scala 117:10]
  wire  _GEN_8671; // @[Execute.scala 117:10]
  wire  _GEN_8672; // @[Execute.scala 117:10]
  wire  _GEN_8673; // @[Execute.scala 117:10]
  wire  _GEN_8674; // @[Execute.scala 117:10]
  wire  _GEN_8676; // @[Execute.scala 117:10]
  wire  _GEN_8677; // @[Execute.scala 117:10]
  wire  _GEN_8678; // @[Execute.scala 117:10]
  wire  _GEN_8679; // @[Execute.scala 117:10]
  wire  _GEN_8680; // @[Execute.scala 117:10]
  wire  _GEN_8681; // @[Execute.scala 117:10]
  wire  _GEN_8682; // @[Execute.scala 117:10]
  wire  _GEN_8683; // @[Execute.scala 117:10]
  wire  _GEN_8684; // @[Execute.scala 117:10]
  wire  _GEN_8685; // @[Execute.scala 117:10]
  wire  _GEN_8686; // @[Execute.scala 117:10]
  wire  _GEN_8687; // @[Execute.scala 117:10]
  wire  _GEN_8688; // @[Execute.scala 117:10]
  wire  _GEN_8689; // @[Execute.scala 117:10]
  wire  _GEN_8690; // @[Execute.scala 117:10]
  wire  _GEN_8691; // @[Execute.scala 117:10]
  wire  _GEN_8692; // @[Execute.scala 117:10]
  wire  _GEN_8693; // @[Execute.scala 117:10]
  wire  _GEN_8694; // @[Execute.scala 117:10]
  wire  _GEN_8695; // @[Execute.scala 117:10]
  wire  _GEN_8696; // @[Execute.scala 117:10]
  wire  _GEN_8697; // @[Execute.scala 117:10]
  wire  _GEN_8698; // @[Execute.scala 117:10]
  wire  _GEN_8699; // @[Execute.scala 117:10]
  wire  _GEN_8700; // @[Execute.scala 117:10]
  wire  _GEN_8701; // @[Execute.scala 117:10]
  wire  _GEN_8702; // @[Execute.scala 117:10]
  wire  _GEN_8703; // @[Execute.scala 117:10]
  wire  _GEN_8704; // @[Execute.scala 117:10]
  wire  _GEN_8705; // @[Execute.scala 117:10]
  wire  _GEN_8706; // @[Execute.scala 117:10]
  wire  _T_863; // @[Execute.scala 117:10]
  wire  _T_864; // @[Execute.scala 117:15]
  wire [4:0] _T_866; // @[Execute.scala 117:37]
  wire [4:0] _T_868; // @[Execute.scala 117:60]
  wire  _GEN_8708; // @[Execute.scala 117:10]
  wire  _GEN_8709; // @[Execute.scala 117:10]
  wire  _GEN_8710; // @[Execute.scala 117:10]
  wire  _GEN_8711; // @[Execute.scala 117:10]
  wire  _GEN_8712; // @[Execute.scala 117:10]
  wire  _GEN_8713; // @[Execute.scala 117:10]
  wire  _GEN_8714; // @[Execute.scala 117:10]
  wire  _GEN_8715; // @[Execute.scala 117:10]
  wire  _GEN_8716; // @[Execute.scala 117:10]
  wire  _GEN_8717; // @[Execute.scala 117:10]
  wire  _GEN_8718; // @[Execute.scala 117:10]
  wire  _GEN_8719; // @[Execute.scala 117:10]
  wire  _GEN_8720; // @[Execute.scala 117:10]
  wire  _GEN_8721; // @[Execute.scala 117:10]
  wire  _GEN_8722; // @[Execute.scala 117:10]
  wire  _GEN_8723; // @[Execute.scala 117:10]
  wire  _GEN_8724; // @[Execute.scala 117:10]
  wire  _GEN_8725; // @[Execute.scala 117:10]
  wire  _GEN_8726; // @[Execute.scala 117:10]
  wire  _GEN_8727; // @[Execute.scala 117:10]
  wire  _GEN_8728; // @[Execute.scala 117:10]
  wire  _GEN_8729; // @[Execute.scala 117:10]
  wire  _GEN_8730; // @[Execute.scala 117:10]
  wire  _GEN_8731; // @[Execute.scala 117:10]
  wire  _GEN_8732; // @[Execute.scala 117:10]
  wire  _GEN_8733; // @[Execute.scala 117:10]
  wire  _GEN_8734; // @[Execute.scala 117:10]
  wire  _GEN_8735; // @[Execute.scala 117:10]
  wire  _GEN_8736; // @[Execute.scala 117:10]
  wire  _GEN_8737; // @[Execute.scala 117:10]
  wire  _GEN_8738; // @[Execute.scala 117:10]
  wire  _GEN_8740; // @[Execute.scala 117:10]
  wire  _GEN_8741; // @[Execute.scala 117:10]
  wire  _GEN_8742; // @[Execute.scala 117:10]
  wire  _GEN_8743; // @[Execute.scala 117:10]
  wire  _GEN_8744; // @[Execute.scala 117:10]
  wire  _GEN_8745; // @[Execute.scala 117:10]
  wire  _GEN_8746; // @[Execute.scala 117:10]
  wire  _GEN_8747; // @[Execute.scala 117:10]
  wire  _GEN_8748; // @[Execute.scala 117:10]
  wire  _GEN_8749; // @[Execute.scala 117:10]
  wire  _GEN_8750; // @[Execute.scala 117:10]
  wire  _GEN_8751; // @[Execute.scala 117:10]
  wire  _GEN_8752; // @[Execute.scala 117:10]
  wire  _GEN_8753; // @[Execute.scala 117:10]
  wire  _GEN_8754; // @[Execute.scala 117:10]
  wire  _GEN_8755; // @[Execute.scala 117:10]
  wire  _GEN_8756; // @[Execute.scala 117:10]
  wire  _GEN_8757; // @[Execute.scala 117:10]
  wire  _GEN_8758; // @[Execute.scala 117:10]
  wire  _GEN_8759; // @[Execute.scala 117:10]
  wire  _GEN_8760; // @[Execute.scala 117:10]
  wire  _GEN_8761; // @[Execute.scala 117:10]
  wire  _GEN_8762; // @[Execute.scala 117:10]
  wire  _GEN_8763; // @[Execute.scala 117:10]
  wire  _GEN_8764; // @[Execute.scala 117:10]
  wire  _GEN_8765; // @[Execute.scala 117:10]
  wire  _GEN_8766; // @[Execute.scala 117:10]
  wire  _GEN_8767; // @[Execute.scala 117:10]
  wire  _GEN_8768; // @[Execute.scala 117:10]
  wire  _GEN_8769; // @[Execute.scala 117:10]
  wire  _GEN_8770; // @[Execute.scala 117:10]
  wire  _T_869; // @[Execute.scala 117:10]
  wire  _T_870; // @[Execute.scala 117:15]
  wire [4:0] _T_872; // @[Execute.scala 117:37]
  wire [4:0] _T_874; // @[Execute.scala 117:60]
  wire  _GEN_8772; // @[Execute.scala 117:10]
  wire  _GEN_8773; // @[Execute.scala 117:10]
  wire  _GEN_8774; // @[Execute.scala 117:10]
  wire  _GEN_8775; // @[Execute.scala 117:10]
  wire  _GEN_8776; // @[Execute.scala 117:10]
  wire  _GEN_8777; // @[Execute.scala 117:10]
  wire  _GEN_8778; // @[Execute.scala 117:10]
  wire  _GEN_8779; // @[Execute.scala 117:10]
  wire  _GEN_8780; // @[Execute.scala 117:10]
  wire  _GEN_8781; // @[Execute.scala 117:10]
  wire  _GEN_8782; // @[Execute.scala 117:10]
  wire  _GEN_8783; // @[Execute.scala 117:10]
  wire  _GEN_8784; // @[Execute.scala 117:10]
  wire  _GEN_8785; // @[Execute.scala 117:10]
  wire  _GEN_8786; // @[Execute.scala 117:10]
  wire  _GEN_8787; // @[Execute.scala 117:10]
  wire  _GEN_8788; // @[Execute.scala 117:10]
  wire  _GEN_8789; // @[Execute.scala 117:10]
  wire  _GEN_8790; // @[Execute.scala 117:10]
  wire  _GEN_8791; // @[Execute.scala 117:10]
  wire  _GEN_8792; // @[Execute.scala 117:10]
  wire  _GEN_8793; // @[Execute.scala 117:10]
  wire  _GEN_8794; // @[Execute.scala 117:10]
  wire  _GEN_8795; // @[Execute.scala 117:10]
  wire  _GEN_8796; // @[Execute.scala 117:10]
  wire  _GEN_8797; // @[Execute.scala 117:10]
  wire  _GEN_8798; // @[Execute.scala 117:10]
  wire  _GEN_8799; // @[Execute.scala 117:10]
  wire  _GEN_8800; // @[Execute.scala 117:10]
  wire  _GEN_8801; // @[Execute.scala 117:10]
  wire  _GEN_8802; // @[Execute.scala 117:10]
  wire  _GEN_8804; // @[Execute.scala 117:10]
  wire  _GEN_8805; // @[Execute.scala 117:10]
  wire  _GEN_8806; // @[Execute.scala 117:10]
  wire  _GEN_8807; // @[Execute.scala 117:10]
  wire  _GEN_8808; // @[Execute.scala 117:10]
  wire  _GEN_8809; // @[Execute.scala 117:10]
  wire  _GEN_8810; // @[Execute.scala 117:10]
  wire  _GEN_8811; // @[Execute.scala 117:10]
  wire  _GEN_8812; // @[Execute.scala 117:10]
  wire  _GEN_8813; // @[Execute.scala 117:10]
  wire  _GEN_8814; // @[Execute.scala 117:10]
  wire  _GEN_8815; // @[Execute.scala 117:10]
  wire  _GEN_8816; // @[Execute.scala 117:10]
  wire  _GEN_8817; // @[Execute.scala 117:10]
  wire  _GEN_8818; // @[Execute.scala 117:10]
  wire  _GEN_8819; // @[Execute.scala 117:10]
  wire  _GEN_8820; // @[Execute.scala 117:10]
  wire  _GEN_8821; // @[Execute.scala 117:10]
  wire  _GEN_8822; // @[Execute.scala 117:10]
  wire  _GEN_8823; // @[Execute.scala 117:10]
  wire  _GEN_8824; // @[Execute.scala 117:10]
  wire  _GEN_8825; // @[Execute.scala 117:10]
  wire  _GEN_8826; // @[Execute.scala 117:10]
  wire  _GEN_8827; // @[Execute.scala 117:10]
  wire  _GEN_8828; // @[Execute.scala 117:10]
  wire  _GEN_8829; // @[Execute.scala 117:10]
  wire  _GEN_8830; // @[Execute.scala 117:10]
  wire  _GEN_8831; // @[Execute.scala 117:10]
  wire  _GEN_8832; // @[Execute.scala 117:10]
  wire  _GEN_8833; // @[Execute.scala 117:10]
  wire  _GEN_8834; // @[Execute.scala 117:10]
  wire  _T_875; // @[Execute.scala 117:10]
  wire  _T_876; // @[Execute.scala 117:15]
  wire [4:0] _T_878; // @[Execute.scala 117:37]
  wire [4:0] _T_880; // @[Execute.scala 117:60]
  wire  _GEN_8836; // @[Execute.scala 117:10]
  wire  _GEN_8837; // @[Execute.scala 117:10]
  wire  _GEN_8838; // @[Execute.scala 117:10]
  wire  _GEN_8839; // @[Execute.scala 117:10]
  wire  _GEN_8840; // @[Execute.scala 117:10]
  wire  _GEN_8841; // @[Execute.scala 117:10]
  wire  _GEN_8842; // @[Execute.scala 117:10]
  wire  _GEN_8843; // @[Execute.scala 117:10]
  wire  _GEN_8844; // @[Execute.scala 117:10]
  wire  _GEN_8845; // @[Execute.scala 117:10]
  wire  _GEN_8846; // @[Execute.scala 117:10]
  wire  _GEN_8847; // @[Execute.scala 117:10]
  wire  _GEN_8848; // @[Execute.scala 117:10]
  wire  _GEN_8849; // @[Execute.scala 117:10]
  wire  _GEN_8850; // @[Execute.scala 117:10]
  wire  _GEN_8851; // @[Execute.scala 117:10]
  wire  _GEN_8852; // @[Execute.scala 117:10]
  wire  _GEN_8853; // @[Execute.scala 117:10]
  wire  _GEN_8854; // @[Execute.scala 117:10]
  wire  _GEN_8855; // @[Execute.scala 117:10]
  wire  _GEN_8856; // @[Execute.scala 117:10]
  wire  _GEN_8857; // @[Execute.scala 117:10]
  wire  _GEN_8858; // @[Execute.scala 117:10]
  wire  _GEN_8859; // @[Execute.scala 117:10]
  wire  _GEN_8860; // @[Execute.scala 117:10]
  wire  _GEN_8861; // @[Execute.scala 117:10]
  wire  _GEN_8862; // @[Execute.scala 117:10]
  wire  _GEN_8863; // @[Execute.scala 117:10]
  wire  _GEN_8864; // @[Execute.scala 117:10]
  wire  _GEN_8865; // @[Execute.scala 117:10]
  wire  _GEN_8866; // @[Execute.scala 117:10]
  wire  _GEN_8868; // @[Execute.scala 117:10]
  wire  _GEN_8869; // @[Execute.scala 117:10]
  wire  _GEN_8870; // @[Execute.scala 117:10]
  wire  _GEN_8871; // @[Execute.scala 117:10]
  wire  _GEN_8872; // @[Execute.scala 117:10]
  wire  _GEN_8873; // @[Execute.scala 117:10]
  wire  _GEN_8874; // @[Execute.scala 117:10]
  wire  _GEN_8875; // @[Execute.scala 117:10]
  wire  _GEN_8876; // @[Execute.scala 117:10]
  wire  _GEN_8877; // @[Execute.scala 117:10]
  wire  _GEN_8878; // @[Execute.scala 117:10]
  wire  _GEN_8879; // @[Execute.scala 117:10]
  wire  _GEN_8880; // @[Execute.scala 117:10]
  wire  _GEN_8881; // @[Execute.scala 117:10]
  wire  _GEN_8882; // @[Execute.scala 117:10]
  wire  _GEN_8883; // @[Execute.scala 117:10]
  wire  _GEN_8884; // @[Execute.scala 117:10]
  wire  _GEN_8885; // @[Execute.scala 117:10]
  wire  _GEN_8886; // @[Execute.scala 117:10]
  wire  _GEN_8887; // @[Execute.scala 117:10]
  wire  _GEN_8888; // @[Execute.scala 117:10]
  wire  _GEN_8889; // @[Execute.scala 117:10]
  wire  _GEN_8890; // @[Execute.scala 117:10]
  wire  _GEN_8891; // @[Execute.scala 117:10]
  wire  _GEN_8892; // @[Execute.scala 117:10]
  wire  _GEN_8893; // @[Execute.scala 117:10]
  wire  _GEN_8894; // @[Execute.scala 117:10]
  wire  _GEN_8895; // @[Execute.scala 117:10]
  wire  _GEN_8896; // @[Execute.scala 117:10]
  wire  _GEN_8897; // @[Execute.scala 117:10]
  wire  _GEN_8898; // @[Execute.scala 117:10]
  wire  _T_881; // @[Execute.scala 117:10]
  wire  _T_882; // @[Execute.scala 117:15]
  wire [4:0] _T_884; // @[Execute.scala 117:37]
  wire [4:0] _T_886; // @[Execute.scala 117:60]
  wire  _GEN_8900; // @[Execute.scala 117:10]
  wire  _GEN_8901; // @[Execute.scala 117:10]
  wire  _GEN_8902; // @[Execute.scala 117:10]
  wire  _GEN_8903; // @[Execute.scala 117:10]
  wire  _GEN_8904; // @[Execute.scala 117:10]
  wire  _GEN_8905; // @[Execute.scala 117:10]
  wire  _GEN_8906; // @[Execute.scala 117:10]
  wire  _GEN_8907; // @[Execute.scala 117:10]
  wire  _GEN_8908; // @[Execute.scala 117:10]
  wire  _GEN_8909; // @[Execute.scala 117:10]
  wire  _GEN_8910; // @[Execute.scala 117:10]
  wire  _GEN_8911; // @[Execute.scala 117:10]
  wire  _GEN_8912; // @[Execute.scala 117:10]
  wire  _GEN_8913; // @[Execute.scala 117:10]
  wire  _GEN_8914; // @[Execute.scala 117:10]
  wire  _GEN_8915; // @[Execute.scala 117:10]
  wire  _GEN_8916; // @[Execute.scala 117:10]
  wire  _GEN_8917; // @[Execute.scala 117:10]
  wire  _GEN_8918; // @[Execute.scala 117:10]
  wire  _GEN_8919; // @[Execute.scala 117:10]
  wire  _GEN_8920; // @[Execute.scala 117:10]
  wire  _GEN_8921; // @[Execute.scala 117:10]
  wire  _GEN_8922; // @[Execute.scala 117:10]
  wire  _GEN_8923; // @[Execute.scala 117:10]
  wire  _GEN_8924; // @[Execute.scala 117:10]
  wire  _GEN_8925; // @[Execute.scala 117:10]
  wire  _GEN_8926; // @[Execute.scala 117:10]
  wire  _GEN_8927; // @[Execute.scala 117:10]
  wire  _GEN_8928; // @[Execute.scala 117:10]
  wire  _GEN_8929; // @[Execute.scala 117:10]
  wire  _GEN_8930; // @[Execute.scala 117:10]
  wire  _GEN_8932; // @[Execute.scala 117:10]
  wire  _GEN_8933; // @[Execute.scala 117:10]
  wire  _GEN_8934; // @[Execute.scala 117:10]
  wire  _GEN_8935; // @[Execute.scala 117:10]
  wire  _GEN_8936; // @[Execute.scala 117:10]
  wire  _GEN_8937; // @[Execute.scala 117:10]
  wire  _GEN_8938; // @[Execute.scala 117:10]
  wire  _GEN_8939; // @[Execute.scala 117:10]
  wire  _GEN_8940; // @[Execute.scala 117:10]
  wire  _GEN_8941; // @[Execute.scala 117:10]
  wire  _GEN_8942; // @[Execute.scala 117:10]
  wire  _GEN_8943; // @[Execute.scala 117:10]
  wire  _GEN_8944; // @[Execute.scala 117:10]
  wire  _GEN_8945; // @[Execute.scala 117:10]
  wire  _GEN_8946; // @[Execute.scala 117:10]
  wire  _GEN_8947; // @[Execute.scala 117:10]
  wire  _GEN_8948; // @[Execute.scala 117:10]
  wire  _GEN_8949; // @[Execute.scala 117:10]
  wire  _GEN_8950; // @[Execute.scala 117:10]
  wire  _GEN_8951; // @[Execute.scala 117:10]
  wire  _GEN_8952; // @[Execute.scala 117:10]
  wire  _GEN_8953; // @[Execute.scala 117:10]
  wire  _GEN_8954; // @[Execute.scala 117:10]
  wire  _GEN_8955; // @[Execute.scala 117:10]
  wire  _GEN_8956; // @[Execute.scala 117:10]
  wire  _GEN_8957; // @[Execute.scala 117:10]
  wire  _GEN_8958; // @[Execute.scala 117:10]
  wire  _GEN_8959; // @[Execute.scala 117:10]
  wire  _GEN_8960; // @[Execute.scala 117:10]
  wire  _GEN_8961; // @[Execute.scala 117:10]
  wire  _GEN_8962; // @[Execute.scala 117:10]
  wire  _T_887; // @[Execute.scala 117:10]
  wire  _T_888; // @[Execute.scala 117:15]
  wire [4:0] _T_890; // @[Execute.scala 117:37]
  wire [4:0] _T_892; // @[Execute.scala 117:60]
  wire  _GEN_8964; // @[Execute.scala 117:10]
  wire  _GEN_8965; // @[Execute.scala 117:10]
  wire  _GEN_8966; // @[Execute.scala 117:10]
  wire  _GEN_8967; // @[Execute.scala 117:10]
  wire  _GEN_8968; // @[Execute.scala 117:10]
  wire  _GEN_8969; // @[Execute.scala 117:10]
  wire  _GEN_8970; // @[Execute.scala 117:10]
  wire  _GEN_8971; // @[Execute.scala 117:10]
  wire  _GEN_8972; // @[Execute.scala 117:10]
  wire  _GEN_8973; // @[Execute.scala 117:10]
  wire  _GEN_8974; // @[Execute.scala 117:10]
  wire  _GEN_8975; // @[Execute.scala 117:10]
  wire  _GEN_8976; // @[Execute.scala 117:10]
  wire  _GEN_8977; // @[Execute.scala 117:10]
  wire  _GEN_8978; // @[Execute.scala 117:10]
  wire  _GEN_8979; // @[Execute.scala 117:10]
  wire  _GEN_8980; // @[Execute.scala 117:10]
  wire  _GEN_8981; // @[Execute.scala 117:10]
  wire  _GEN_8982; // @[Execute.scala 117:10]
  wire  _GEN_8983; // @[Execute.scala 117:10]
  wire  _GEN_8984; // @[Execute.scala 117:10]
  wire  _GEN_8985; // @[Execute.scala 117:10]
  wire  _GEN_8986; // @[Execute.scala 117:10]
  wire  _GEN_8987; // @[Execute.scala 117:10]
  wire  _GEN_8988; // @[Execute.scala 117:10]
  wire  _GEN_8989; // @[Execute.scala 117:10]
  wire  _GEN_8990; // @[Execute.scala 117:10]
  wire  _GEN_8991; // @[Execute.scala 117:10]
  wire  _GEN_8992; // @[Execute.scala 117:10]
  wire  _GEN_8993; // @[Execute.scala 117:10]
  wire  _GEN_8994; // @[Execute.scala 117:10]
  wire  _GEN_8996; // @[Execute.scala 117:10]
  wire  _GEN_8997; // @[Execute.scala 117:10]
  wire  _GEN_8998; // @[Execute.scala 117:10]
  wire  _GEN_8999; // @[Execute.scala 117:10]
  wire  _GEN_9000; // @[Execute.scala 117:10]
  wire  _GEN_9001; // @[Execute.scala 117:10]
  wire  _GEN_9002; // @[Execute.scala 117:10]
  wire  _GEN_9003; // @[Execute.scala 117:10]
  wire  _GEN_9004; // @[Execute.scala 117:10]
  wire  _GEN_9005; // @[Execute.scala 117:10]
  wire  _GEN_9006; // @[Execute.scala 117:10]
  wire  _GEN_9007; // @[Execute.scala 117:10]
  wire  _GEN_9008; // @[Execute.scala 117:10]
  wire  _GEN_9009; // @[Execute.scala 117:10]
  wire  _GEN_9010; // @[Execute.scala 117:10]
  wire  _GEN_9011; // @[Execute.scala 117:10]
  wire  _GEN_9012; // @[Execute.scala 117:10]
  wire  _GEN_9013; // @[Execute.scala 117:10]
  wire  _GEN_9014; // @[Execute.scala 117:10]
  wire  _GEN_9015; // @[Execute.scala 117:10]
  wire  _GEN_9016; // @[Execute.scala 117:10]
  wire  _GEN_9017; // @[Execute.scala 117:10]
  wire  _GEN_9018; // @[Execute.scala 117:10]
  wire  _GEN_9019; // @[Execute.scala 117:10]
  wire  _GEN_9020; // @[Execute.scala 117:10]
  wire  _GEN_9021; // @[Execute.scala 117:10]
  wire  _GEN_9022; // @[Execute.scala 117:10]
  wire  _GEN_9023; // @[Execute.scala 117:10]
  wire  _GEN_9024; // @[Execute.scala 117:10]
  wire  _GEN_9025; // @[Execute.scala 117:10]
  wire  _GEN_9026; // @[Execute.scala 117:10]
  wire  _T_893; // @[Execute.scala 117:10]
  wire  _T_894; // @[Execute.scala 117:15]
  wire [4:0] _T_896; // @[Execute.scala 117:37]
  wire [4:0] _T_898; // @[Execute.scala 117:60]
  wire  _GEN_9028; // @[Execute.scala 117:10]
  wire  _GEN_9029; // @[Execute.scala 117:10]
  wire  _GEN_9030; // @[Execute.scala 117:10]
  wire  _GEN_9031; // @[Execute.scala 117:10]
  wire  _GEN_9032; // @[Execute.scala 117:10]
  wire  _GEN_9033; // @[Execute.scala 117:10]
  wire  _GEN_9034; // @[Execute.scala 117:10]
  wire  _GEN_9035; // @[Execute.scala 117:10]
  wire  _GEN_9036; // @[Execute.scala 117:10]
  wire  _GEN_9037; // @[Execute.scala 117:10]
  wire  _GEN_9038; // @[Execute.scala 117:10]
  wire  _GEN_9039; // @[Execute.scala 117:10]
  wire  _GEN_9040; // @[Execute.scala 117:10]
  wire  _GEN_9041; // @[Execute.scala 117:10]
  wire  _GEN_9042; // @[Execute.scala 117:10]
  wire  _GEN_9043; // @[Execute.scala 117:10]
  wire  _GEN_9044; // @[Execute.scala 117:10]
  wire  _GEN_9045; // @[Execute.scala 117:10]
  wire  _GEN_9046; // @[Execute.scala 117:10]
  wire  _GEN_9047; // @[Execute.scala 117:10]
  wire  _GEN_9048; // @[Execute.scala 117:10]
  wire  _GEN_9049; // @[Execute.scala 117:10]
  wire  _GEN_9050; // @[Execute.scala 117:10]
  wire  _GEN_9051; // @[Execute.scala 117:10]
  wire  _GEN_9052; // @[Execute.scala 117:10]
  wire  _GEN_9053; // @[Execute.scala 117:10]
  wire  _GEN_9054; // @[Execute.scala 117:10]
  wire  _GEN_9055; // @[Execute.scala 117:10]
  wire  _GEN_9056; // @[Execute.scala 117:10]
  wire  _GEN_9057; // @[Execute.scala 117:10]
  wire  _GEN_9058; // @[Execute.scala 117:10]
  wire  _GEN_9060; // @[Execute.scala 117:10]
  wire  _GEN_9061; // @[Execute.scala 117:10]
  wire  _GEN_9062; // @[Execute.scala 117:10]
  wire  _GEN_9063; // @[Execute.scala 117:10]
  wire  _GEN_9064; // @[Execute.scala 117:10]
  wire  _GEN_9065; // @[Execute.scala 117:10]
  wire  _GEN_9066; // @[Execute.scala 117:10]
  wire  _GEN_9067; // @[Execute.scala 117:10]
  wire  _GEN_9068; // @[Execute.scala 117:10]
  wire  _GEN_9069; // @[Execute.scala 117:10]
  wire  _GEN_9070; // @[Execute.scala 117:10]
  wire  _GEN_9071; // @[Execute.scala 117:10]
  wire  _GEN_9072; // @[Execute.scala 117:10]
  wire  _GEN_9073; // @[Execute.scala 117:10]
  wire  _GEN_9074; // @[Execute.scala 117:10]
  wire  _GEN_9075; // @[Execute.scala 117:10]
  wire  _GEN_9076; // @[Execute.scala 117:10]
  wire  _GEN_9077; // @[Execute.scala 117:10]
  wire  _GEN_9078; // @[Execute.scala 117:10]
  wire  _GEN_9079; // @[Execute.scala 117:10]
  wire  _GEN_9080; // @[Execute.scala 117:10]
  wire  _GEN_9081; // @[Execute.scala 117:10]
  wire  _GEN_9082; // @[Execute.scala 117:10]
  wire  _GEN_9083; // @[Execute.scala 117:10]
  wire  _GEN_9084; // @[Execute.scala 117:10]
  wire  _GEN_9085; // @[Execute.scala 117:10]
  wire  _GEN_9086; // @[Execute.scala 117:10]
  wire  _GEN_9087; // @[Execute.scala 117:10]
  wire  _GEN_9088; // @[Execute.scala 117:10]
  wire  _GEN_9089; // @[Execute.scala 117:10]
  wire  _GEN_9090; // @[Execute.scala 117:10]
  wire  _T_899; // @[Execute.scala 117:10]
  wire  _T_900; // @[Execute.scala 117:15]
  wire [4:0] _T_902; // @[Execute.scala 117:37]
  wire [4:0] _T_904; // @[Execute.scala 117:60]
  wire  _GEN_9092; // @[Execute.scala 117:10]
  wire  _GEN_9093; // @[Execute.scala 117:10]
  wire  _GEN_9094; // @[Execute.scala 117:10]
  wire  _GEN_9095; // @[Execute.scala 117:10]
  wire  _GEN_9096; // @[Execute.scala 117:10]
  wire  _GEN_9097; // @[Execute.scala 117:10]
  wire  _GEN_9098; // @[Execute.scala 117:10]
  wire  _GEN_9099; // @[Execute.scala 117:10]
  wire  _GEN_9100; // @[Execute.scala 117:10]
  wire  _GEN_9101; // @[Execute.scala 117:10]
  wire  _GEN_9102; // @[Execute.scala 117:10]
  wire  _GEN_9103; // @[Execute.scala 117:10]
  wire  _GEN_9104; // @[Execute.scala 117:10]
  wire  _GEN_9105; // @[Execute.scala 117:10]
  wire  _GEN_9106; // @[Execute.scala 117:10]
  wire  _GEN_9107; // @[Execute.scala 117:10]
  wire  _GEN_9108; // @[Execute.scala 117:10]
  wire  _GEN_9109; // @[Execute.scala 117:10]
  wire  _GEN_9110; // @[Execute.scala 117:10]
  wire  _GEN_9111; // @[Execute.scala 117:10]
  wire  _GEN_9112; // @[Execute.scala 117:10]
  wire  _GEN_9113; // @[Execute.scala 117:10]
  wire  _GEN_9114; // @[Execute.scala 117:10]
  wire  _GEN_9115; // @[Execute.scala 117:10]
  wire  _GEN_9116; // @[Execute.scala 117:10]
  wire  _GEN_9117; // @[Execute.scala 117:10]
  wire  _GEN_9118; // @[Execute.scala 117:10]
  wire  _GEN_9119; // @[Execute.scala 117:10]
  wire  _GEN_9120; // @[Execute.scala 117:10]
  wire  _GEN_9121; // @[Execute.scala 117:10]
  wire  _GEN_9122; // @[Execute.scala 117:10]
  wire  _GEN_9124; // @[Execute.scala 117:10]
  wire  _GEN_9125; // @[Execute.scala 117:10]
  wire  _GEN_9126; // @[Execute.scala 117:10]
  wire  _GEN_9127; // @[Execute.scala 117:10]
  wire  _GEN_9128; // @[Execute.scala 117:10]
  wire  _GEN_9129; // @[Execute.scala 117:10]
  wire  _GEN_9130; // @[Execute.scala 117:10]
  wire  _GEN_9131; // @[Execute.scala 117:10]
  wire  _GEN_9132; // @[Execute.scala 117:10]
  wire  _GEN_9133; // @[Execute.scala 117:10]
  wire  _GEN_9134; // @[Execute.scala 117:10]
  wire  _GEN_9135; // @[Execute.scala 117:10]
  wire  _GEN_9136; // @[Execute.scala 117:10]
  wire  _GEN_9137; // @[Execute.scala 117:10]
  wire  _GEN_9138; // @[Execute.scala 117:10]
  wire  _GEN_9139; // @[Execute.scala 117:10]
  wire  _GEN_9140; // @[Execute.scala 117:10]
  wire  _GEN_9141; // @[Execute.scala 117:10]
  wire  _GEN_9142; // @[Execute.scala 117:10]
  wire  _GEN_9143; // @[Execute.scala 117:10]
  wire  _GEN_9144; // @[Execute.scala 117:10]
  wire  _GEN_9145; // @[Execute.scala 117:10]
  wire  _GEN_9146; // @[Execute.scala 117:10]
  wire  _GEN_9147; // @[Execute.scala 117:10]
  wire  _GEN_9148; // @[Execute.scala 117:10]
  wire  _GEN_9149; // @[Execute.scala 117:10]
  wire  _GEN_9150; // @[Execute.scala 117:10]
  wire  _GEN_9151; // @[Execute.scala 117:10]
  wire  _GEN_9152; // @[Execute.scala 117:10]
  wire  _GEN_9153; // @[Execute.scala 117:10]
  wire  _GEN_9154; // @[Execute.scala 117:10]
  wire  _T_905; // @[Execute.scala 117:10]
  wire  _T_906; // @[Execute.scala 117:15]
  wire [4:0] _T_908; // @[Execute.scala 117:37]
  wire [4:0] _T_910; // @[Execute.scala 117:60]
  wire  _GEN_9156; // @[Execute.scala 117:10]
  wire  _GEN_9157; // @[Execute.scala 117:10]
  wire  _GEN_9158; // @[Execute.scala 117:10]
  wire  _GEN_9159; // @[Execute.scala 117:10]
  wire  _GEN_9160; // @[Execute.scala 117:10]
  wire  _GEN_9161; // @[Execute.scala 117:10]
  wire  _GEN_9162; // @[Execute.scala 117:10]
  wire  _GEN_9163; // @[Execute.scala 117:10]
  wire  _GEN_9164; // @[Execute.scala 117:10]
  wire  _GEN_9165; // @[Execute.scala 117:10]
  wire  _GEN_9166; // @[Execute.scala 117:10]
  wire  _GEN_9167; // @[Execute.scala 117:10]
  wire  _GEN_9168; // @[Execute.scala 117:10]
  wire  _GEN_9169; // @[Execute.scala 117:10]
  wire  _GEN_9170; // @[Execute.scala 117:10]
  wire  _GEN_9171; // @[Execute.scala 117:10]
  wire  _GEN_9172; // @[Execute.scala 117:10]
  wire  _GEN_9173; // @[Execute.scala 117:10]
  wire  _GEN_9174; // @[Execute.scala 117:10]
  wire  _GEN_9175; // @[Execute.scala 117:10]
  wire  _GEN_9176; // @[Execute.scala 117:10]
  wire  _GEN_9177; // @[Execute.scala 117:10]
  wire  _GEN_9178; // @[Execute.scala 117:10]
  wire  _GEN_9179; // @[Execute.scala 117:10]
  wire  _GEN_9180; // @[Execute.scala 117:10]
  wire  _GEN_9181; // @[Execute.scala 117:10]
  wire  _GEN_9182; // @[Execute.scala 117:10]
  wire  _GEN_9183; // @[Execute.scala 117:10]
  wire  _GEN_9184; // @[Execute.scala 117:10]
  wire  _GEN_9185; // @[Execute.scala 117:10]
  wire  _GEN_9186; // @[Execute.scala 117:10]
  wire  _GEN_9188; // @[Execute.scala 117:10]
  wire  _GEN_9189; // @[Execute.scala 117:10]
  wire  _GEN_9190; // @[Execute.scala 117:10]
  wire  _GEN_9191; // @[Execute.scala 117:10]
  wire  _GEN_9192; // @[Execute.scala 117:10]
  wire  _GEN_9193; // @[Execute.scala 117:10]
  wire  _GEN_9194; // @[Execute.scala 117:10]
  wire  _GEN_9195; // @[Execute.scala 117:10]
  wire  _GEN_9196; // @[Execute.scala 117:10]
  wire  _GEN_9197; // @[Execute.scala 117:10]
  wire  _GEN_9198; // @[Execute.scala 117:10]
  wire  _GEN_9199; // @[Execute.scala 117:10]
  wire  _GEN_9200; // @[Execute.scala 117:10]
  wire  _GEN_9201; // @[Execute.scala 117:10]
  wire  _GEN_9202; // @[Execute.scala 117:10]
  wire  _GEN_9203; // @[Execute.scala 117:10]
  wire  _GEN_9204; // @[Execute.scala 117:10]
  wire  _GEN_9205; // @[Execute.scala 117:10]
  wire  _GEN_9206; // @[Execute.scala 117:10]
  wire  _GEN_9207; // @[Execute.scala 117:10]
  wire  _GEN_9208; // @[Execute.scala 117:10]
  wire  _GEN_9209; // @[Execute.scala 117:10]
  wire  _GEN_9210; // @[Execute.scala 117:10]
  wire  _GEN_9211; // @[Execute.scala 117:10]
  wire  _GEN_9212; // @[Execute.scala 117:10]
  wire  _GEN_9213; // @[Execute.scala 117:10]
  wire  _GEN_9214; // @[Execute.scala 117:10]
  wire  _GEN_9215; // @[Execute.scala 117:10]
  wire  _GEN_9216; // @[Execute.scala 117:10]
  wire  _GEN_9217; // @[Execute.scala 117:10]
  wire  _GEN_9218; // @[Execute.scala 117:10]
  wire  _T_911; // @[Execute.scala 117:10]
  wire  _T_912; // @[Execute.scala 117:15]
  wire [4:0] _T_914; // @[Execute.scala 117:37]
  wire [4:0] _T_916; // @[Execute.scala 117:60]
  wire  _GEN_9220; // @[Execute.scala 117:10]
  wire  _GEN_9221; // @[Execute.scala 117:10]
  wire  _GEN_9222; // @[Execute.scala 117:10]
  wire  _GEN_9223; // @[Execute.scala 117:10]
  wire  _GEN_9224; // @[Execute.scala 117:10]
  wire  _GEN_9225; // @[Execute.scala 117:10]
  wire  _GEN_9226; // @[Execute.scala 117:10]
  wire  _GEN_9227; // @[Execute.scala 117:10]
  wire  _GEN_9228; // @[Execute.scala 117:10]
  wire  _GEN_9229; // @[Execute.scala 117:10]
  wire  _GEN_9230; // @[Execute.scala 117:10]
  wire  _GEN_9231; // @[Execute.scala 117:10]
  wire  _GEN_9232; // @[Execute.scala 117:10]
  wire  _GEN_9233; // @[Execute.scala 117:10]
  wire  _GEN_9234; // @[Execute.scala 117:10]
  wire  _GEN_9235; // @[Execute.scala 117:10]
  wire  _GEN_9236; // @[Execute.scala 117:10]
  wire  _GEN_9237; // @[Execute.scala 117:10]
  wire  _GEN_9238; // @[Execute.scala 117:10]
  wire  _GEN_9239; // @[Execute.scala 117:10]
  wire  _GEN_9240; // @[Execute.scala 117:10]
  wire  _GEN_9241; // @[Execute.scala 117:10]
  wire  _GEN_9242; // @[Execute.scala 117:10]
  wire  _GEN_9243; // @[Execute.scala 117:10]
  wire  _GEN_9244; // @[Execute.scala 117:10]
  wire  _GEN_9245; // @[Execute.scala 117:10]
  wire  _GEN_9246; // @[Execute.scala 117:10]
  wire  _GEN_9247; // @[Execute.scala 117:10]
  wire  _GEN_9248; // @[Execute.scala 117:10]
  wire  _GEN_9249; // @[Execute.scala 117:10]
  wire  _GEN_9250; // @[Execute.scala 117:10]
  wire  _GEN_9252; // @[Execute.scala 117:10]
  wire  _GEN_9253; // @[Execute.scala 117:10]
  wire  _GEN_9254; // @[Execute.scala 117:10]
  wire  _GEN_9255; // @[Execute.scala 117:10]
  wire  _GEN_9256; // @[Execute.scala 117:10]
  wire  _GEN_9257; // @[Execute.scala 117:10]
  wire  _GEN_9258; // @[Execute.scala 117:10]
  wire  _GEN_9259; // @[Execute.scala 117:10]
  wire  _GEN_9260; // @[Execute.scala 117:10]
  wire  _GEN_9261; // @[Execute.scala 117:10]
  wire  _GEN_9262; // @[Execute.scala 117:10]
  wire  _GEN_9263; // @[Execute.scala 117:10]
  wire  _GEN_9264; // @[Execute.scala 117:10]
  wire  _GEN_9265; // @[Execute.scala 117:10]
  wire  _GEN_9266; // @[Execute.scala 117:10]
  wire  _GEN_9267; // @[Execute.scala 117:10]
  wire  _GEN_9268; // @[Execute.scala 117:10]
  wire  _GEN_9269; // @[Execute.scala 117:10]
  wire  _GEN_9270; // @[Execute.scala 117:10]
  wire  _GEN_9271; // @[Execute.scala 117:10]
  wire  _GEN_9272; // @[Execute.scala 117:10]
  wire  _GEN_9273; // @[Execute.scala 117:10]
  wire  _GEN_9274; // @[Execute.scala 117:10]
  wire  _GEN_9275; // @[Execute.scala 117:10]
  wire  _GEN_9276; // @[Execute.scala 117:10]
  wire  _GEN_9277; // @[Execute.scala 117:10]
  wire  _GEN_9278; // @[Execute.scala 117:10]
  wire  _GEN_9279; // @[Execute.scala 117:10]
  wire  _GEN_9280; // @[Execute.scala 117:10]
  wire  _GEN_9281; // @[Execute.scala 117:10]
  wire  _GEN_9282; // @[Execute.scala 117:10]
  wire  _T_917; // @[Execute.scala 117:10]
  wire  _T_918; // @[Execute.scala 117:15]
  wire [4:0] _T_920; // @[Execute.scala 117:37]
  wire [4:0] _T_922; // @[Execute.scala 117:60]
  wire  _GEN_9284; // @[Execute.scala 117:10]
  wire  _GEN_9285; // @[Execute.scala 117:10]
  wire  _GEN_9286; // @[Execute.scala 117:10]
  wire  _GEN_9287; // @[Execute.scala 117:10]
  wire  _GEN_9288; // @[Execute.scala 117:10]
  wire  _GEN_9289; // @[Execute.scala 117:10]
  wire  _GEN_9290; // @[Execute.scala 117:10]
  wire  _GEN_9291; // @[Execute.scala 117:10]
  wire  _GEN_9292; // @[Execute.scala 117:10]
  wire  _GEN_9293; // @[Execute.scala 117:10]
  wire  _GEN_9294; // @[Execute.scala 117:10]
  wire  _GEN_9295; // @[Execute.scala 117:10]
  wire  _GEN_9296; // @[Execute.scala 117:10]
  wire  _GEN_9297; // @[Execute.scala 117:10]
  wire  _GEN_9298; // @[Execute.scala 117:10]
  wire  _GEN_9299; // @[Execute.scala 117:10]
  wire  _GEN_9300; // @[Execute.scala 117:10]
  wire  _GEN_9301; // @[Execute.scala 117:10]
  wire  _GEN_9302; // @[Execute.scala 117:10]
  wire  _GEN_9303; // @[Execute.scala 117:10]
  wire  _GEN_9304; // @[Execute.scala 117:10]
  wire  _GEN_9305; // @[Execute.scala 117:10]
  wire  _GEN_9306; // @[Execute.scala 117:10]
  wire  _GEN_9307; // @[Execute.scala 117:10]
  wire  _GEN_9308; // @[Execute.scala 117:10]
  wire  _GEN_9309; // @[Execute.scala 117:10]
  wire  _GEN_9310; // @[Execute.scala 117:10]
  wire  _GEN_9311; // @[Execute.scala 117:10]
  wire  _GEN_9312; // @[Execute.scala 117:10]
  wire  _GEN_9313; // @[Execute.scala 117:10]
  wire  _GEN_9314; // @[Execute.scala 117:10]
  wire  _GEN_9316; // @[Execute.scala 117:10]
  wire  _GEN_9317; // @[Execute.scala 117:10]
  wire  _GEN_9318; // @[Execute.scala 117:10]
  wire  _GEN_9319; // @[Execute.scala 117:10]
  wire  _GEN_9320; // @[Execute.scala 117:10]
  wire  _GEN_9321; // @[Execute.scala 117:10]
  wire  _GEN_9322; // @[Execute.scala 117:10]
  wire  _GEN_9323; // @[Execute.scala 117:10]
  wire  _GEN_9324; // @[Execute.scala 117:10]
  wire  _GEN_9325; // @[Execute.scala 117:10]
  wire  _GEN_9326; // @[Execute.scala 117:10]
  wire  _GEN_9327; // @[Execute.scala 117:10]
  wire  _GEN_9328; // @[Execute.scala 117:10]
  wire  _GEN_9329; // @[Execute.scala 117:10]
  wire  _GEN_9330; // @[Execute.scala 117:10]
  wire  _GEN_9331; // @[Execute.scala 117:10]
  wire  _GEN_9332; // @[Execute.scala 117:10]
  wire  _GEN_9333; // @[Execute.scala 117:10]
  wire  _GEN_9334; // @[Execute.scala 117:10]
  wire  _GEN_9335; // @[Execute.scala 117:10]
  wire  _GEN_9336; // @[Execute.scala 117:10]
  wire  _GEN_9337; // @[Execute.scala 117:10]
  wire  _GEN_9338; // @[Execute.scala 117:10]
  wire  _GEN_9339; // @[Execute.scala 117:10]
  wire  _GEN_9340; // @[Execute.scala 117:10]
  wire  _GEN_9341; // @[Execute.scala 117:10]
  wire  _GEN_9342; // @[Execute.scala 117:10]
  wire  _GEN_9343; // @[Execute.scala 117:10]
  wire  _GEN_9344; // @[Execute.scala 117:10]
  wire  _GEN_9345; // @[Execute.scala 117:10]
  wire  _GEN_9346; // @[Execute.scala 117:10]
  wire  _T_923; // @[Execute.scala 117:10]
  wire  _T_924; // @[Execute.scala 117:15]
  wire [4:0] _T_926; // @[Execute.scala 117:37]
  wire [4:0] _T_928; // @[Execute.scala 117:60]
  wire  _GEN_9348; // @[Execute.scala 117:10]
  wire  _GEN_9349; // @[Execute.scala 117:10]
  wire  _GEN_9350; // @[Execute.scala 117:10]
  wire  _GEN_9351; // @[Execute.scala 117:10]
  wire  _GEN_9352; // @[Execute.scala 117:10]
  wire  _GEN_9353; // @[Execute.scala 117:10]
  wire  _GEN_9354; // @[Execute.scala 117:10]
  wire  _GEN_9355; // @[Execute.scala 117:10]
  wire  _GEN_9356; // @[Execute.scala 117:10]
  wire  _GEN_9357; // @[Execute.scala 117:10]
  wire  _GEN_9358; // @[Execute.scala 117:10]
  wire  _GEN_9359; // @[Execute.scala 117:10]
  wire  _GEN_9360; // @[Execute.scala 117:10]
  wire  _GEN_9361; // @[Execute.scala 117:10]
  wire  _GEN_9362; // @[Execute.scala 117:10]
  wire  _GEN_9363; // @[Execute.scala 117:10]
  wire  _GEN_9364; // @[Execute.scala 117:10]
  wire  _GEN_9365; // @[Execute.scala 117:10]
  wire  _GEN_9366; // @[Execute.scala 117:10]
  wire  _GEN_9367; // @[Execute.scala 117:10]
  wire  _GEN_9368; // @[Execute.scala 117:10]
  wire  _GEN_9369; // @[Execute.scala 117:10]
  wire  _GEN_9370; // @[Execute.scala 117:10]
  wire  _GEN_9371; // @[Execute.scala 117:10]
  wire  _GEN_9372; // @[Execute.scala 117:10]
  wire  _GEN_9373; // @[Execute.scala 117:10]
  wire  _GEN_9374; // @[Execute.scala 117:10]
  wire  _GEN_9375; // @[Execute.scala 117:10]
  wire  _GEN_9376; // @[Execute.scala 117:10]
  wire  _GEN_9377; // @[Execute.scala 117:10]
  wire  _GEN_9378; // @[Execute.scala 117:10]
  wire  _GEN_9380; // @[Execute.scala 117:10]
  wire  _GEN_9381; // @[Execute.scala 117:10]
  wire  _GEN_9382; // @[Execute.scala 117:10]
  wire  _GEN_9383; // @[Execute.scala 117:10]
  wire  _GEN_9384; // @[Execute.scala 117:10]
  wire  _GEN_9385; // @[Execute.scala 117:10]
  wire  _GEN_9386; // @[Execute.scala 117:10]
  wire  _GEN_9387; // @[Execute.scala 117:10]
  wire  _GEN_9388; // @[Execute.scala 117:10]
  wire  _GEN_9389; // @[Execute.scala 117:10]
  wire  _GEN_9390; // @[Execute.scala 117:10]
  wire  _GEN_9391; // @[Execute.scala 117:10]
  wire  _GEN_9392; // @[Execute.scala 117:10]
  wire  _GEN_9393; // @[Execute.scala 117:10]
  wire  _GEN_9394; // @[Execute.scala 117:10]
  wire  _GEN_9395; // @[Execute.scala 117:10]
  wire  _GEN_9396; // @[Execute.scala 117:10]
  wire  _GEN_9397; // @[Execute.scala 117:10]
  wire  _GEN_9398; // @[Execute.scala 117:10]
  wire  _GEN_9399; // @[Execute.scala 117:10]
  wire  _GEN_9400; // @[Execute.scala 117:10]
  wire  _GEN_9401; // @[Execute.scala 117:10]
  wire  _GEN_9402; // @[Execute.scala 117:10]
  wire  _GEN_9403; // @[Execute.scala 117:10]
  wire  _GEN_9404; // @[Execute.scala 117:10]
  wire  _GEN_9405; // @[Execute.scala 117:10]
  wire  _GEN_9406; // @[Execute.scala 117:10]
  wire  _GEN_9407; // @[Execute.scala 117:10]
  wire  _GEN_9408; // @[Execute.scala 117:10]
  wire  _GEN_9409; // @[Execute.scala 117:10]
  wire  _GEN_9410; // @[Execute.scala 117:10]
  wire  _T_929; // @[Execute.scala 117:10]
  wire  _T_930; // @[Execute.scala 117:15]
  wire [4:0] _T_932; // @[Execute.scala 117:37]
  wire [4:0] _T_934; // @[Execute.scala 117:60]
  wire  _GEN_9412; // @[Execute.scala 117:10]
  wire  _GEN_9413; // @[Execute.scala 117:10]
  wire  _GEN_9414; // @[Execute.scala 117:10]
  wire  _GEN_9415; // @[Execute.scala 117:10]
  wire  _GEN_9416; // @[Execute.scala 117:10]
  wire  _GEN_9417; // @[Execute.scala 117:10]
  wire  _GEN_9418; // @[Execute.scala 117:10]
  wire  _GEN_9419; // @[Execute.scala 117:10]
  wire  _GEN_9420; // @[Execute.scala 117:10]
  wire  _GEN_9421; // @[Execute.scala 117:10]
  wire  _GEN_9422; // @[Execute.scala 117:10]
  wire  _GEN_9423; // @[Execute.scala 117:10]
  wire  _GEN_9424; // @[Execute.scala 117:10]
  wire  _GEN_9425; // @[Execute.scala 117:10]
  wire  _GEN_9426; // @[Execute.scala 117:10]
  wire  _GEN_9427; // @[Execute.scala 117:10]
  wire  _GEN_9428; // @[Execute.scala 117:10]
  wire  _GEN_9429; // @[Execute.scala 117:10]
  wire  _GEN_9430; // @[Execute.scala 117:10]
  wire  _GEN_9431; // @[Execute.scala 117:10]
  wire  _GEN_9432; // @[Execute.scala 117:10]
  wire  _GEN_9433; // @[Execute.scala 117:10]
  wire  _GEN_9434; // @[Execute.scala 117:10]
  wire  _GEN_9435; // @[Execute.scala 117:10]
  wire  _GEN_9436; // @[Execute.scala 117:10]
  wire  _GEN_9437; // @[Execute.scala 117:10]
  wire  _GEN_9438; // @[Execute.scala 117:10]
  wire  _GEN_9439; // @[Execute.scala 117:10]
  wire  _GEN_9440; // @[Execute.scala 117:10]
  wire  _GEN_9441; // @[Execute.scala 117:10]
  wire  _GEN_9442; // @[Execute.scala 117:10]
  wire  _GEN_9444; // @[Execute.scala 117:10]
  wire  _GEN_9445; // @[Execute.scala 117:10]
  wire  _GEN_9446; // @[Execute.scala 117:10]
  wire  _GEN_9447; // @[Execute.scala 117:10]
  wire  _GEN_9448; // @[Execute.scala 117:10]
  wire  _GEN_9449; // @[Execute.scala 117:10]
  wire  _GEN_9450; // @[Execute.scala 117:10]
  wire  _GEN_9451; // @[Execute.scala 117:10]
  wire  _GEN_9452; // @[Execute.scala 117:10]
  wire  _GEN_9453; // @[Execute.scala 117:10]
  wire  _GEN_9454; // @[Execute.scala 117:10]
  wire  _GEN_9455; // @[Execute.scala 117:10]
  wire  _GEN_9456; // @[Execute.scala 117:10]
  wire  _GEN_9457; // @[Execute.scala 117:10]
  wire  _GEN_9458; // @[Execute.scala 117:10]
  wire  _GEN_9459; // @[Execute.scala 117:10]
  wire  _GEN_9460; // @[Execute.scala 117:10]
  wire  _GEN_9461; // @[Execute.scala 117:10]
  wire  _GEN_9462; // @[Execute.scala 117:10]
  wire  _GEN_9463; // @[Execute.scala 117:10]
  wire  _GEN_9464; // @[Execute.scala 117:10]
  wire  _GEN_9465; // @[Execute.scala 117:10]
  wire  _GEN_9466; // @[Execute.scala 117:10]
  wire  _GEN_9467; // @[Execute.scala 117:10]
  wire  _GEN_9468; // @[Execute.scala 117:10]
  wire  _GEN_9469; // @[Execute.scala 117:10]
  wire  _GEN_9470; // @[Execute.scala 117:10]
  wire  _GEN_9471; // @[Execute.scala 117:10]
  wire  _GEN_9472; // @[Execute.scala 117:10]
  wire  _GEN_9473; // @[Execute.scala 117:10]
  wire  _GEN_9474; // @[Execute.scala 117:10]
  wire  _T_935; // @[Execute.scala 117:10]
  wire  _T_936; // @[Execute.scala 117:15]
  wire [4:0] _T_938; // @[Execute.scala 117:37]
  wire [4:0] _T_940; // @[Execute.scala 117:60]
  wire  _GEN_9476; // @[Execute.scala 117:10]
  wire  _GEN_9477; // @[Execute.scala 117:10]
  wire  _GEN_9478; // @[Execute.scala 117:10]
  wire  _GEN_9479; // @[Execute.scala 117:10]
  wire  _GEN_9480; // @[Execute.scala 117:10]
  wire  _GEN_9481; // @[Execute.scala 117:10]
  wire  _GEN_9482; // @[Execute.scala 117:10]
  wire  _GEN_9483; // @[Execute.scala 117:10]
  wire  _GEN_9484; // @[Execute.scala 117:10]
  wire  _GEN_9485; // @[Execute.scala 117:10]
  wire  _GEN_9486; // @[Execute.scala 117:10]
  wire  _GEN_9487; // @[Execute.scala 117:10]
  wire  _GEN_9488; // @[Execute.scala 117:10]
  wire  _GEN_9489; // @[Execute.scala 117:10]
  wire  _GEN_9490; // @[Execute.scala 117:10]
  wire  _GEN_9491; // @[Execute.scala 117:10]
  wire  _GEN_9492; // @[Execute.scala 117:10]
  wire  _GEN_9493; // @[Execute.scala 117:10]
  wire  _GEN_9494; // @[Execute.scala 117:10]
  wire  _GEN_9495; // @[Execute.scala 117:10]
  wire  _GEN_9496; // @[Execute.scala 117:10]
  wire  _GEN_9497; // @[Execute.scala 117:10]
  wire  _GEN_9498; // @[Execute.scala 117:10]
  wire  _GEN_9499; // @[Execute.scala 117:10]
  wire  _GEN_9500; // @[Execute.scala 117:10]
  wire  _GEN_9501; // @[Execute.scala 117:10]
  wire  _GEN_9502; // @[Execute.scala 117:10]
  wire  _GEN_9503; // @[Execute.scala 117:10]
  wire  _GEN_9504; // @[Execute.scala 117:10]
  wire  _GEN_9505; // @[Execute.scala 117:10]
  wire  _GEN_9506; // @[Execute.scala 117:10]
  wire  _GEN_9508; // @[Execute.scala 117:10]
  wire  _GEN_9509; // @[Execute.scala 117:10]
  wire  _GEN_9510; // @[Execute.scala 117:10]
  wire  _GEN_9511; // @[Execute.scala 117:10]
  wire  _GEN_9512; // @[Execute.scala 117:10]
  wire  _GEN_9513; // @[Execute.scala 117:10]
  wire  _GEN_9514; // @[Execute.scala 117:10]
  wire  _GEN_9515; // @[Execute.scala 117:10]
  wire  _GEN_9516; // @[Execute.scala 117:10]
  wire  _GEN_9517; // @[Execute.scala 117:10]
  wire  _GEN_9518; // @[Execute.scala 117:10]
  wire  _GEN_9519; // @[Execute.scala 117:10]
  wire  _GEN_9520; // @[Execute.scala 117:10]
  wire  _GEN_9521; // @[Execute.scala 117:10]
  wire  _GEN_9522; // @[Execute.scala 117:10]
  wire  _GEN_9523; // @[Execute.scala 117:10]
  wire  _GEN_9524; // @[Execute.scala 117:10]
  wire  _GEN_9525; // @[Execute.scala 117:10]
  wire  _GEN_9526; // @[Execute.scala 117:10]
  wire  _GEN_9527; // @[Execute.scala 117:10]
  wire  _GEN_9528; // @[Execute.scala 117:10]
  wire  _GEN_9529; // @[Execute.scala 117:10]
  wire  _GEN_9530; // @[Execute.scala 117:10]
  wire  _GEN_9531; // @[Execute.scala 117:10]
  wire  _GEN_9532; // @[Execute.scala 117:10]
  wire  _GEN_9533; // @[Execute.scala 117:10]
  wire  _GEN_9534; // @[Execute.scala 117:10]
  wire  _GEN_9535; // @[Execute.scala 117:10]
  wire  _GEN_9536; // @[Execute.scala 117:10]
  wire  _GEN_9537; // @[Execute.scala 117:10]
  wire  _GEN_9538; // @[Execute.scala 117:10]
  wire  _T_941; // @[Execute.scala 117:10]
  wire  _T_942; // @[Execute.scala 117:15]
  wire [4:0] _T_944; // @[Execute.scala 117:37]
  wire [4:0] _T_946; // @[Execute.scala 117:60]
  wire  _GEN_9540; // @[Execute.scala 117:10]
  wire  _GEN_9541; // @[Execute.scala 117:10]
  wire  _GEN_9542; // @[Execute.scala 117:10]
  wire  _GEN_9543; // @[Execute.scala 117:10]
  wire  _GEN_9544; // @[Execute.scala 117:10]
  wire  _GEN_9545; // @[Execute.scala 117:10]
  wire  _GEN_9546; // @[Execute.scala 117:10]
  wire  _GEN_9547; // @[Execute.scala 117:10]
  wire  _GEN_9548; // @[Execute.scala 117:10]
  wire  _GEN_9549; // @[Execute.scala 117:10]
  wire  _GEN_9550; // @[Execute.scala 117:10]
  wire  _GEN_9551; // @[Execute.scala 117:10]
  wire  _GEN_9552; // @[Execute.scala 117:10]
  wire  _GEN_9553; // @[Execute.scala 117:10]
  wire  _GEN_9554; // @[Execute.scala 117:10]
  wire  _GEN_9555; // @[Execute.scala 117:10]
  wire  _GEN_9556; // @[Execute.scala 117:10]
  wire  _GEN_9557; // @[Execute.scala 117:10]
  wire  _GEN_9558; // @[Execute.scala 117:10]
  wire  _GEN_9559; // @[Execute.scala 117:10]
  wire  _GEN_9560; // @[Execute.scala 117:10]
  wire  _GEN_9561; // @[Execute.scala 117:10]
  wire  _GEN_9562; // @[Execute.scala 117:10]
  wire  _GEN_9563; // @[Execute.scala 117:10]
  wire  _GEN_9564; // @[Execute.scala 117:10]
  wire  _GEN_9565; // @[Execute.scala 117:10]
  wire  _GEN_9566; // @[Execute.scala 117:10]
  wire  _GEN_9567; // @[Execute.scala 117:10]
  wire  _GEN_9568; // @[Execute.scala 117:10]
  wire  _GEN_9569; // @[Execute.scala 117:10]
  wire  _GEN_9570; // @[Execute.scala 117:10]
  wire  _GEN_9572; // @[Execute.scala 117:10]
  wire  _GEN_9573; // @[Execute.scala 117:10]
  wire  _GEN_9574; // @[Execute.scala 117:10]
  wire  _GEN_9575; // @[Execute.scala 117:10]
  wire  _GEN_9576; // @[Execute.scala 117:10]
  wire  _GEN_9577; // @[Execute.scala 117:10]
  wire  _GEN_9578; // @[Execute.scala 117:10]
  wire  _GEN_9579; // @[Execute.scala 117:10]
  wire  _GEN_9580; // @[Execute.scala 117:10]
  wire  _GEN_9581; // @[Execute.scala 117:10]
  wire  _GEN_9582; // @[Execute.scala 117:10]
  wire  _GEN_9583; // @[Execute.scala 117:10]
  wire  _GEN_9584; // @[Execute.scala 117:10]
  wire  _GEN_9585; // @[Execute.scala 117:10]
  wire  _GEN_9586; // @[Execute.scala 117:10]
  wire  _GEN_9587; // @[Execute.scala 117:10]
  wire  _GEN_9588; // @[Execute.scala 117:10]
  wire  _GEN_9589; // @[Execute.scala 117:10]
  wire  _GEN_9590; // @[Execute.scala 117:10]
  wire  _GEN_9591; // @[Execute.scala 117:10]
  wire  _GEN_9592; // @[Execute.scala 117:10]
  wire  _GEN_9593; // @[Execute.scala 117:10]
  wire  _GEN_9594; // @[Execute.scala 117:10]
  wire  _GEN_9595; // @[Execute.scala 117:10]
  wire  _GEN_9596; // @[Execute.scala 117:10]
  wire  _GEN_9597; // @[Execute.scala 117:10]
  wire  _GEN_9598; // @[Execute.scala 117:10]
  wire  _GEN_9599; // @[Execute.scala 117:10]
  wire  _GEN_9600; // @[Execute.scala 117:10]
  wire  _GEN_9601; // @[Execute.scala 117:10]
  wire  _GEN_9602; // @[Execute.scala 117:10]
  wire  _T_947; // @[Execute.scala 117:10]
  wire  _T_948; // @[Execute.scala 117:15]
  wire [4:0] _T_950; // @[Execute.scala 117:37]
  wire [4:0] _T_952; // @[Execute.scala 117:60]
  wire  _GEN_9604; // @[Execute.scala 117:10]
  wire  _GEN_9605; // @[Execute.scala 117:10]
  wire  _GEN_9606; // @[Execute.scala 117:10]
  wire  _GEN_9607; // @[Execute.scala 117:10]
  wire  _GEN_9608; // @[Execute.scala 117:10]
  wire  _GEN_9609; // @[Execute.scala 117:10]
  wire  _GEN_9610; // @[Execute.scala 117:10]
  wire  _GEN_9611; // @[Execute.scala 117:10]
  wire  _GEN_9612; // @[Execute.scala 117:10]
  wire  _GEN_9613; // @[Execute.scala 117:10]
  wire  _GEN_9614; // @[Execute.scala 117:10]
  wire  _GEN_9615; // @[Execute.scala 117:10]
  wire  _GEN_9616; // @[Execute.scala 117:10]
  wire  _GEN_9617; // @[Execute.scala 117:10]
  wire  _GEN_9618; // @[Execute.scala 117:10]
  wire  _GEN_9619; // @[Execute.scala 117:10]
  wire  _GEN_9620; // @[Execute.scala 117:10]
  wire  _GEN_9621; // @[Execute.scala 117:10]
  wire  _GEN_9622; // @[Execute.scala 117:10]
  wire  _GEN_9623; // @[Execute.scala 117:10]
  wire  _GEN_9624; // @[Execute.scala 117:10]
  wire  _GEN_9625; // @[Execute.scala 117:10]
  wire  _GEN_9626; // @[Execute.scala 117:10]
  wire  _GEN_9627; // @[Execute.scala 117:10]
  wire  _GEN_9628; // @[Execute.scala 117:10]
  wire  _GEN_9629; // @[Execute.scala 117:10]
  wire  _GEN_9630; // @[Execute.scala 117:10]
  wire  _GEN_9631; // @[Execute.scala 117:10]
  wire  _GEN_9632; // @[Execute.scala 117:10]
  wire  _GEN_9633; // @[Execute.scala 117:10]
  wire  _GEN_9634; // @[Execute.scala 117:10]
  wire  _GEN_9636; // @[Execute.scala 117:10]
  wire  _GEN_9637; // @[Execute.scala 117:10]
  wire  _GEN_9638; // @[Execute.scala 117:10]
  wire  _GEN_9639; // @[Execute.scala 117:10]
  wire  _GEN_9640; // @[Execute.scala 117:10]
  wire  _GEN_9641; // @[Execute.scala 117:10]
  wire  _GEN_9642; // @[Execute.scala 117:10]
  wire  _GEN_9643; // @[Execute.scala 117:10]
  wire  _GEN_9644; // @[Execute.scala 117:10]
  wire  _GEN_9645; // @[Execute.scala 117:10]
  wire  _GEN_9646; // @[Execute.scala 117:10]
  wire  _GEN_9647; // @[Execute.scala 117:10]
  wire  _GEN_9648; // @[Execute.scala 117:10]
  wire  _GEN_9649; // @[Execute.scala 117:10]
  wire  _GEN_9650; // @[Execute.scala 117:10]
  wire  _GEN_9651; // @[Execute.scala 117:10]
  wire  _GEN_9652; // @[Execute.scala 117:10]
  wire  _GEN_9653; // @[Execute.scala 117:10]
  wire  _GEN_9654; // @[Execute.scala 117:10]
  wire  _GEN_9655; // @[Execute.scala 117:10]
  wire  _GEN_9656; // @[Execute.scala 117:10]
  wire  _GEN_9657; // @[Execute.scala 117:10]
  wire  _GEN_9658; // @[Execute.scala 117:10]
  wire  _GEN_9659; // @[Execute.scala 117:10]
  wire  _GEN_9660; // @[Execute.scala 117:10]
  wire  _GEN_9661; // @[Execute.scala 117:10]
  wire  _GEN_9662; // @[Execute.scala 117:10]
  wire  _GEN_9663; // @[Execute.scala 117:10]
  wire  _GEN_9664; // @[Execute.scala 117:10]
  wire  _GEN_9665; // @[Execute.scala 117:10]
  wire  _GEN_9666; // @[Execute.scala 117:10]
  wire  _T_953; // @[Execute.scala 117:10]
  wire  _T_954; // @[Execute.scala 117:15]
  wire [4:0] _T_956; // @[Execute.scala 117:37]
  wire [4:0] _T_958; // @[Execute.scala 117:60]
  wire  _GEN_9668; // @[Execute.scala 117:10]
  wire  _GEN_9669; // @[Execute.scala 117:10]
  wire  _GEN_9670; // @[Execute.scala 117:10]
  wire  _GEN_9671; // @[Execute.scala 117:10]
  wire  _GEN_9672; // @[Execute.scala 117:10]
  wire  _GEN_9673; // @[Execute.scala 117:10]
  wire  _GEN_9674; // @[Execute.scala 117:10]
  wire  _GEN_9675; // @[Execute.scala 117:10]
  wire  _GEN_9676; // @[Execute.scala 117:10]
  wire  _GEN_9677; // @[Execute.scala 117:10]
  wire  _GEN_9678; // @[Execute.scala 117:10]
  wire  _GEN_9679; // @[Execute.scala 117:10]
  wire  _GEN_9680; // @[Execute.scala 117:10]
  wire  _GEN_9681; // @[Execute.scala 117:10]
  wire  _GEN_9682; // @[Execute.scala 117:10]
  wire  _GEN_9683; // @[Execute.scala 117:10]
  wire  _GEN_9684; // @[Execute.scala 117:10]
  wire  _GEN_9685; // @[Execute.scala 117:10]
  wire  _GEN_9686; // @[Execute.scala 117:10]
  wire  _GEN_9687; // @[Execute.scala 117:10]
  wire  _GEN_9688; // @[Execute.scala 117:10]
  wire  _GEN_9689; // @[Execute.scala 117:10]
  wire  _GEN_9690; // @[Execute.scala 117:10]
  wire  _GEN_9691; // @[Execute.scala 117:10]
  wire  _GEN_9692; // @[Execute.scala 117:10]
  wire  _GEN_9693; // @[Execute.scala 117:10]
  wire  _GEN_9694; // @[Execute.scala 117:10]
  wire  _GEN_9695; // @[Execute.scala 117:10]
  wire  _GEN_9696; // @[Execute.scala 117:10]
  wire  _GEN_9697; // @[Execute.scala 117:10]
  wire  _GEN_9698; // @[Execute.scala 117:10]
  wire  _GEN_9700; // @[Execute.scala 117:10]
  wire  _GEN_9701; // @[Execute.scala 117:10]
  wire  _GEN_9702; // @[Execute.scala 117:10]
  wire  _GEN_9703; // @[Execute.scala 117:10]
  wire  _GEN_9704; // @[Execute.scala 117:10]
  wire  _GEN_9705; // @[Execute.scala 117:10]
  wire  _GEN_9706; // @[Execute.scala 117:10]
  wire  _GEN_9707; // @[Execute.scala 117:10]
  wire  _GEN_9708; // @[Execute.scala 117:10]
  wire  _GEN_9709; // @[Execute.scala 117:10]
  wire  _GEN_9710; // @[Execute.scala 117:10]
  wire  _GEN_9711; // @[Execute.scala 117:10]
  wire  _GEN_9712; // @[Execute.scala 117:10]
  wire  _GEN_9713; // @[Execute.scala 117:10]
  wire  _GEN_9714; // @[Execute.scala 117:10]
  wire  _GEN_9715; // @[Execute.scala 117:10]
  wire  _GEN_9716; // @[Execute.scala 117:10]
  wire  _GEN_9717; // @[Execute.scala 117:10]
  wire  _GEN_9718; // @[Execute.scala 117:10]
  wire  _GEN_9719; // @[Execute.scala 117:10]
  wire  _GEN_9720; // @[Execute.scala 117:10]
  wire  _GEN_9721; // @[Execute.scala 117:10]
  wire  _GEN_9722; // @[Execute.scala 117:10]
  wire  _GEN_9723; // @[Execute.scala 117:10]
  wire  _GEN_9724; // @[Execute.scala 117:10]
  wire  _GEN_9725; // @[Execute.scala 117:10]
  wire  _GEN_9726; // @[Execute.scala 117:10]
  wire  _GEN_9727; // @[Execute.scala 117:10]
  wire  _GEN_9728; // @[Execute.scala 117:10]
  wire  _GEN_9729; // @[Execute.scala 117:10]
  wire  _GEN_9730; // @[Execute.scala 117:10]
  wire  _T_959; // @[Execute.scala 117:10]
  wire  _T_960; // @[Execute.scala 117:15]
  wire [4:0] _T_962; // @[Execute.scala 117:37]
  wire [4:0] _T_964; // @[Execute.scala 117:60]
  wire  _GEN_9732; // @[Execute.scala 117:10]
  wire  _GEN_9733; // @[Execute.scala 117:10]
  wire  _GEN_9734; // @[Execute.scala 117:10]
  wire  _GEN_9735; // @[Execute.scala 117:10]
  wire  _GEN_9736; // @[Execute.scala 117:10]
  wire  _GEN_9737; // @[Execute.scala 117:10]
  wire  _GEN_9738; // @[Execute.scala 117:10]
  wire  _GEN_9739; // @[Execute.scala 117:10]
  wire  _GEN_9740; // @[Execute.scala 117:10]
  wire  _GEN_9741; // @[Execute.scala 117:10]
  wire  _GEN_9742; // @[Execute.scala 117:10]
  wire  _GEN_9743; // @[Execute.scala 117:10]
  wire  _GEN_9744; // @[Execute.scala 117:10]
  wire  _GEN_9745; // @[Execute.scala 117:10]
  wire  _GEN_9746; // @[Execute.scala 117:10]
  wire  _GEN_9747; // @[Execute.scala 117:10]
  wire  _GEN_9748; // @[Execute.scala 117:10]
  wire  _GEN_9749; // @[Execute.scala 117:10]
  wire  _GEN_9750; // @[Execute.scala 117:10]
  wire  _GEN_9751; // @[Execute.scala 117:10]
  wire  _GEN_9752; // @[Execute.scala 117:10]
  wire  _GEN_9753; // @[Execute.scala 117:10]
  wire  _GEN_9754; // @[Execute.scala 117:10]
  wire  _GEN_9755; // @[Execute.scala 117:10]
  wire  _GEN_9756; // @[Execute.scala 117:10]
  wire  _GEN_9757; // @[Execute.scala 117:10]
  wire  _GEN_9758; // @[Execute.scala 117:10]
  wire  _GEN_9759; // @[Execute.scala 117:10]
  wire  _GEN_9760; // @[Execute.scala 117:10]
  wire  _GEN_9761; // @[Execute.scala 117:10]
  wire  _GEN_9762; // @[Execute.scala 117:10]
  wire  _GEN_9764; // @[Execute.scala 117:10]
  wire  _GEN_9765; // @[Execute.scala 117:10]
  wire  _GEN_9766; // @[Execute.scala 117:10]
  wire  _GEN_9767; // @[Execute.scala 117:10]
  wire  _GEN_9768; // @[Execute.scala 117:10]
  wire  _GEN_9769; // @[Execute.scala 117:10]
  wire  _GEN_9770; // @[Execute.scala 117:10]
  wire  _GEN_9771; // @[Execute.scala 117:10]
  wire  _GEN_9772; // @[Execute.scala 117:10]
  wire  _GEN_9773; // @[Execute.scala 117:10]
  wire  _GEN_9774; // @[Execute.scala 117:10]
  wire  _GEN_9775; // @[Execute.scala 117:10]
  wire  _GEN_9776; // @[Execute.scala 117:10]
  wire  _GEN_9777; // @[Execute.scala 117:10]
  wire  _GEN_9778; // @[Execute.scala 117:10]
  wire  _GEN_9779; // @[Execute.scala 117:10]
  wire  _GEN_9780; // @[Execute.scala 117:10]
  wire  _GEN_9781; // @[Execute.scala 117:10]
  wire  _GEN_9782; // @[Execute.scala 117:10]
  wire  _GEN_9783; // @[Execute.scala 117:10]
  wire  _GEN_9784; // @[Execute.scala 117:10]
  wire  _GEN_9785; // @[Execute.scala 117:10]
  wire  _GEN_9786; // @[Execute.scala 117:10]
  wire  _GEN_9787; // @[Execute.scala 117:10]
  wire  _GEN_9788; // @[Execute.scala 117:10]
  wire  _GEN_9789; // @[Execute.scala 117:10]
  wire  _GEN_9790; // @[Execute.scala 117:10]
  wire  _GEN_9791; // @[Execute.scala 117:10]
  wire  _GEN_9792; // @[Execute.scala 117:10]
  wire  _GEN_9793; // @[Execute.scala 117:10]
  wire  _GEN_9794; // @[Execute.scala 117:10]
  wire  _T_965; // @[Execute.scala 117:10]
  wire  _T_966; // @[Execute.scala 117:15]
  wire [4:0] _T_968; // @[Execute.scala 117:37]
  wire [4:0] _T_970; // @[Execute.scala 117:60]
  wire  _GEN_9796; // @[Execute.scala 117:10]
  wire  _GEN_9797; // @[Execute.scala 117:10]
  wire  _GEN_9798; // @[Execute.scala 117:10]
  wire  _GEN_9799; // @[Execute.scala 117:10]
  wire  _GEN_9800; // @[Execute.scala 117:10]
  wire  _GEN_9801; // @[Execute.scala 117:10]
  wire  _GEN_9802; // @[Execute.scala 117:10]
  wire  _GEN_9803; // @[Execute.scala 117:10]
  wire  _GEN_9804; // @[Execute.scala 117:10]
  wire  _GEN_9805; // @[Execute.scala 117:10]
  wire  _GEN_9806; // @[Execute.scala 117:10]
  wire  _GEN_9807; // @[Execute.scala 117:10]
  wire  _GEN_9808; // @[Execute.scala 117:10]
  wire  _GEN_9809; // @[Execute.scala 117:10]
  wire  _GEN_9810; // @[Execute.scala 117:10]
  wire  _GEN_9811; // @[Execute.scala 117:10]
  wire  _GEN_9812; // @[Execute.scala 117:10]
  wire  _GEN_9813; // @[Execute.scala 117:10]
  wire  _GEN_9814; // @[Execute.scala 117:10]
  wire  _GEN_9815; // @[Execute.scala 117:10]
  wire  _GEN_9816; // @[Execute.scala 117:10]
  wire  _GEN_9817; // @[Execute.scala 117:10]
  wire  _GEN_9818; // @[Execute.scala 117:10]
  wire  _GEN_9819; // @[Execute.scala 117:10]
  wire  _GEN_9820; // @[Execute.scala 117:10]
  wire  _GEN_9821; // @[Execute.scala 117:10]
  wire  _GEN_9822; // @[Execute.scala 117:10]
  wire  _GEN_9823; // @[Execute.scala 117:10]
  wire  _GEN_9824; // @[Execute.scala 117:10]
  wire  _GEN_9825; // @[Execute.scala 117:10]
  wire  _GEN_9826; // @[Execute.scala 117:10]
  wire  _GEN_9828; // @[Execute.scala 117:10]
  wire  _GEN_9829; // @[Execute.scala 117:10]
  wire  _GEN_9830; // @[Execute.scala 117:10]
  wire  _GEN_9831; // @[Execute.scala 117:10]
  wire  _GEN_9832; // @[Execute.scala 117:10]
  wire  _GEN_9833; // @[Execute.scala 117:10]
  wire  _GEN_9834; // @[Execute.scala 117:10]
  wire  _GEN_9835; // @[Execute.scala 117:10]
  wire  _GEN_9836; // @[Execute.scala 117:10]
  wire  _GEN_9837; // @[Execute.scala 117:10]
  wire  _GEN_9838; // @[Execute.scala 117:10]
  wire  _GEN_9839; // @[Execute.scala 117:10]
  wire  _GEN_9840; // @[Execute.scala 117:10]
  wire  _GEN_9841; // @[Execute.scala 117:10]
  wire  _GEN_9842; // @[Execute.scala 117:10]
  wire  _GEN_9843; // @[Execute.scala 117:10]
  wire  _GEN_9844; // @[Execute.scala 117:10]
  wire  _GEN_9845; // @[Execute.scala 117:10]
  wire  _GEN_9846; // @[Execute.scala 117:10]
  wire  _GEN_9847; // @[Execute.scala 117:10]
  wire  _GEN_9848; // @[Execute.scala 117:10]
  wire  _GEN_9849; // @[Execute.scala 117:10]
  wire  _GEN_9850; // @[Execute.scala 117:10]
  wire  _GEN_9851; // @[Execute.scala 117:10]
  wire  _GEN_9852; // @[Execute.scala 117:10]
  wire  _GEN_9853; // @[Execute.scala 117:10]
  wire  _GEN_9854; // @[Execute.scala 117:10]
  wire  _GEN_9855; // @[Execute.scala 117:10]
  wire  _GEN_9856; // @[Execute.scala 117:10]
  wire  _GEN_9857; // @[Execute.scala 117:10]
  wire  _GEN_9858; // @[Execute.scala 117:10]
  wire  _T_971; // @[Execute.scala 117:10]
  wire  _T_972; // @[Execute.scala 117:15]
  wire [4:0] _T_974; // @[Execute.scala 117:37]
  wire [4:0] _T_976; // @[Execute.scala 117:60]
  wire  _GEN_9860; // @[Execute.scala 117:10]
  wire  _GEN_9861; // @[Execute.scala 117:10]
  wire  _GEN_9862; // @[Execute.scala 117:10]
  wire  _GEN_9863; // @[Execute.scala 117:10]
  wire  _GEN_9864; // @[Execute.scala 117:10]
  wire  _GEN_9865; // @[Execute.scala 117:10]
  wire  _GEN_9866; // @[Execute.scala 117:10]
  wire  _GEN_9867; // @[Execute.scala 117:10]
  wire  _GEN_9868; // @[Execute.scala 117:10]
  wire  _GEN_9869; // @[Execute.scala 117:10]
  wire  _GEN_9870; // @[Execute.scala 117:10]
  wire  _GEN_9871; // @[Execute.scala 117:10]
  wire  _GEN_9872; // @[Execute.scala 117:10]
  wire  _GEN_9873; // @[Execute.scala 117:10]
  wire  _GEN_9874; // @[Execute.scala 117:10]
  wire  _GEN_9875; // @[Execute.scala 117:10]
  wire  _GEN_9876; // @[Execute.scala 117:10]
  wire  _GEN_9877; // @[Execute.scala 117:10]
  wire  _GEN_9878; // @[Execute.scala 117:10]
  wire  _GEN_9879; // @[Execute.scala 117:10]
  wire  _GEN_9880; // @[Execute.scala 117:10]
  wire  _GEN_9881; // @[Execute.scala 117:10]
  wire  _GEN_9882; // @[Execute.scala 117:10]
  wire  _GEN_9883; // @[Execute.scala 117:10]
  wire  _GEN_9884; // @[Execute.scala 117:10]
  wire  _GEN_9885; // @[Execute.scala 117:10]
  wire  _GEN_9886; // @[Execute.scala 117:10]
  wire  _GEN_9887; // @[Execute.scala 117:10]
  wire  _GEN_9888; // @[Execute.scala 117:10]
  wire  _GEN_9889; // @[Execute.scala 117:10]
  wire  _GEN_9890; // @[Execute.scala 117:10]
  wire  _GEN_9892; // @[Execute.scala 117:10]
  wire  _GEN_9893; // @[Execute.scala 117:10]
  wire  _GEN_9894; // @[Execute.scala 117:10]
  wire  _GEN_9895; // @[Execute.scala 117:10]
  wire  _GEN_9896; // @[Execute.scala 117:10]
  wire  _GEN_9897; // @[Execute.scala 117:10]
  wire  _GEN_9898; // @[Execute.scala 117:10]
  wire  _GEN_9899; // @[Execute.scala 117:10]
  wire  _GEN_9900; // @[Execute.scala 117:10]
  wire  _GEN_9901; // @[Execute.scala 117:10]
  wire  _GEN_9902; // @[Execute.scala 117:10]
  wire  _GEN_9903; // @[Execute.scala 117:10]
  wire  _GEN_9904; // @[Execute.scala 117:10]
  wire  _GEN_9905; // @[Execute.scala 117:10]
  wire  _GEN_9906; // @[Execute.scala 117:10]
  wire  _GEN_9907; // @[Execute.scala 117:10]
  wire  _GEN_9908; // @[Execute.scala 117:10]
  wire  _GEN_9909; // @[Execute.scala 117:10]
  wire  _GEN_9910; // @[Execute.scala 117:10]
  wire  _GEN_9911; // @[Execute.scala 117:10]
  wire  _GEN_9912; // @[Execute.scala 117:10]
  wire  _GEN_9913; // @[Execute.scala 117:10]
  wire  _GEN_9914; // @[Execute.scala 117:10]
  wire  _GEN_9915; // @[Execute.scala 117:10]
  wire  _GEN_9916; // @[Execute.scala 117:10]
  wire  _GEN_9917; // @[Execute.scala 117:10]
  wire  _GEN_9918; // @[Execute.scala 117:10]
  wire  _GEN_9919; // @[Execute.scala 117:10]
  wire  _GEN_9920; // @[Execute.scala 117:10]
  wire  _GEN_9921; // @[Execute.scala 117:10]
  wire  _GEN_9922; // @[Execute.scala 117:10]
  wire  _T_977; // @[Execute.scala 117:10]
  wire  _T_978; // @[Execute.scala 117:15]
  wire [4:0] _T_980; // @[Execute.scala 117:37]
  wire [4:0] _T_982; // @[Execute.scala 117:60]
  wire  _GEN_9924; // @[Execute.scala 117:10]
  wire  _GEN_9925; // @[Execute.scala 117:10]
  wire  _GEN_9926; // @[Execute.scala 117:10]
  wire  _GEN_9927; // @[Execute.scala 117:10]
  wire  _GEN_9928; // @[Execute.scala 117:10]
  wire  _GEN_9929; // @[Execute.scala 117:10]
  wire  _GEN_9930; // @[Execute.scala 117:10]
  wire  _GEN_9931; // @[Execute.scala 117:10]
  wire  _GEN_9932; // @[Execute.scala 117:10]
  wire  _GEN_9933; // @[Execute.scala 117:10]
  wire  _GEN_9934; // @[Execute.scala 117:10]
  wire  _GEN_9935; // @[Execute.scala 117:10]
  wire  _GEN_9936; // @[Execute.scala 117:10]
  wire  _GEN_9937; // @[Execute.scala 117:10]
  wire  _GEN_9938; // @[Execute.scala 117:10]
  wire  _GEN_9939; // @[Execute.scala 117:10]
  wire  _GEN_9940; // @[Execute.scala 117:10]
  wire  _GEN_9941; // @[Execute.scala 117:10]
  wire  _GEN_9942; // @[Execute.scala 117:10]
  wire  _GEN_9943; // @[Execute.scala 117:10]
  wire  _GEN_9944; // @[Execute.scala 117:10]
  wire  _GEN_9945; // @[Execute.scala 117:10]
  wire  _GEN_9946; // @[Execute.scala 117:10]
  wire  _GEN_9947; // @[Execute.scala 117:10]
  wire  _GEN_9948; // @[Execute.scala 117:10]
  wire  _GEN_9949; // @[Execute.scala 117:10]
  wire  _GEN_9950; // @[Execute.scala 117:10]
  wire  _GEN_9951; // @[Execute.scala 117:10]
  wire  _GEN_9952; // @[Execute.scala 117:10]
  wire  _GEN_9953; // @[Execute.scala 117:10]
  wire  _GEN_9954; // @[Execute.scala 117:10]
  wire  _GEN_9956; // @[Execute.scala 117:10]
  wire  _GEN_9957; // @[Execute.scala 117:10]
  wire  _GEN_9958; // @[Execute.scala 117:10]
  wire  _GEN_9959; // @[Execute.scala 117:10]
  wire  _GEN_9960; // @[Execute.scala 117:10]
  wire  _GEN_9961; // @[Execute.scala 117:10]
  wire  _GEN_9962; // @[Execute.scala 117:10]
  wire  _GEN_9963; // @[Execute.scala 117:10]
  wire  _GEN_9964; // @[Execute.scala 117:10]
  wire  _GEN_9965; // @[Execute.scala 117:10]
  wire  _GEN_9966; // @[Execute.scala 117:10]
  wire  _GEN_9967; // @[Execute.scala 117:10]
  wire  _GEN_9968; // @[Execute.scala 117:10]
  wire  _GEN_9969; // @[Execute.scala 117:10]
  wire  _GEN_9970; // @[Execute.scala 117:10]
  wire  _GEN_9971; // @[Execute.scala 117:10]
  wire  _GEN_9972; // @[Execute.scala 117:10]
  wire  _GEN_9973; // @[Execute.scala 117:10]
  wire  _GEN_9974; // @[Execute.scala 117:10]
  wire  _GEN_9975; // @[Execute.scala 117:10]
  wire  _GEN_9976; // @[Execute.scala 117:10]
  wire  _GEN_9977; // @[Execute.scala 117:10]
  wire  _GEN_9978; // @[Execute.scala 117:10]
  wire  _GEN_9979; // @[Execute.scala 117:10]
  wire  _GEN_9980; // @[Execute.scala 117:10]
  wire  _GEN_9981; // @[Execute.scala 117:10]
  wire  _GEN_9982; // @[Execute.scala 117:10]
  wire  _GEN_9983; // @[Execute.scala 117:10]
  wire  _GEN_9984; // @[Execute.scala 117:10]
  wire  _GEN_9985; // @[Execute.scala 117:10]
  wire  _GEN_9986; // @[Execute.scala 117:10]
  wire  _T_983; // @[Execute.scala 117:10]
  wire  _T_984; // @[Execute.scala 117:15]
  wire [4:0] _T_986; // @[Execute.scala 117:37]
  wire [4:0] _T_988; // @[Execute.scala 117:60]
  wire  _GEN_9988; // @[Execute.scala 117:10]
  wire  _GEN_9989; // @[Execute.scala 117:10]
  wire  _GEN_9990; // @[Execute.scala 117:10]
  wire  _GEN_9991; // @[Execute.scala 117:10]
  wire  _GEN_9992; // @[Execute.scala 117:10]
  wire  _GEN_9993; // @[Execute.scala 117:10]
  wire  _GEN_9994; // @[Execute.scala 117:10]
  wire  _GEN_9995; // @[Execute.scala 117:10]
  wire  _GEN_9996; // @[Execute.scala 117:10]
  wire  _GEN_9997; // @[Execute.scala 117:10]
  wire  _GEN_9998; // @[Execute.scala 117:10]
  wire  _GEN_9999; // @[Execute.scala 117:10]
  wire  _GEN_10000; // @[Execute.scala 117:10]
  wire  _GEN_10001; // @[Execute.scala 117:10]
  wire  _GEN_10002; // @[Execute.scala 117:10]
  wire  _GEN_10003; // @[Execute.scala 117:10]
  wire  _GEN_10004; // @[Execute.scala 117:10]
  wire  _GEN_10005; // @[Execute.scala 117:10]
  wire  _GEN_10006; // @[Execute.scala 117:10]
  wire  _GEN_10007; // @[Execute.scala 117:10]
  wire  _GEN_10008; // @[Execute.scala 117:10]
  wire  _GEN_10009; // @[Execute.scala 117:10]
  wire  _GEN_10010; // @[Execute.scala 117:10]
  wire  _GEN_10011; // @[Execute.scala 117:10]
  wire  _GEN_10012; // @[Execute.scala 117:10]
  wire  _GEN_10013; // @[Execute.scala 117:10]
  wire  _GEN_10014; // @[Execute.scala 117:10]
  wire  _GEN_10015; // @[Execute.scala 117:10]
  wire  _GEN_10016; // @[Execute.scala 117:10]
  wire  _GEN_10017; // @[Execute.scala 117:10]
  wire  _GEN_10018; // @[Execute.scala 117:10]
  wire  _GEN_10020; // @[Execute.scala 117:10]
  wire  _GEN_10021; // @[Execute.scala 117:10]
  wire  _GEN_10022; // @[Execute.scala 117:10]
  wire  _GEN_10023; // @[Execute.scala 117:10]
  wire  _GEN_10024; // @[Execute.scala 117:10]
  wire  _GEN_10025; // @[Execute.scala 117:10]
  wire  _GEN_10026; // @[Execute.scala 117:10]
  wire  _GEN_10027; // @[Execute.scala 117:10]
  wire  _GEN_10028; // @[Execute.scala 117:10]
  wire  _GEN_10029; // @[Execute.scala 117:10]
  wire  _GEN_10030; // @[Execute.scala 117:10]
  wire  _GEN_10031; // @[Execute.scala 117:10]
  wire  _GEN_10032; // @[Execute.scala 117:10]
  wire  _GEN_10033; // @[Execute.scala 117:10]
  wire  _GEN_10034; // @[Execute.scala 117:10]
  wire  _GEN_10035; // @[Execute.scala 117:10]
  wire  _GEN_10036; // @[Execute.scala 117:10]
  wire  _GEN_10037; // @[Execute.scala 117:10]
  wire  _GEN_10038; // @[Execute.scala 117:10]
  wire  _GEN_10039; // @[Execute.scala 117:10]
  wire  _GEN_10040; // @[Execute.scala 117:10]
  wire  _GEN_10041; // @[Execute.scala 117:10]
  wire  _GEN_10042; // @[Execute.scala 117:10]
  wire  _GEN_10043; // @[Execute.scala 117:10]
  wire  _GEN_10044; // @[Execute.scala 117:10]
  wire  _GEN_10045; // @[Execute.scala 117:10]
  wire  _GEN_10046; // @[Execute.scala 117:10]
  wire  _GEN_10047; // @[Execute.scala 117:10]
  wire  _GEN_10048; // @[Execute.scala 117:10]
  wire  _GEN_10049; // @[Execute.scala 117:10]
  wire  _GEN_10050; // @[Execute.scala 117:10]
  wire  _T_989; // @[Execute.scala 117:10]
  wire  _T_990; // @[Execute.scala 117:15]
  wire [4:0] _T_992; // @[Execute.scala 117:37]
  wire [4:0] _T_994; // @[Execute.scala 117:60]
  wire  _GEN_10052; // @[Execute.scala 117:10]
  wire  _GEN_10053; // @[Execute.scala 117:10]
  wire  _GEN_10054; // @[Execute.scala 117:10]
  wire  _GEN_10055; // @[Execute.scala 117:10]
  wire  _GEN_10056; // @[Execute.scala 117:10]
  wire  _GEN_10057; // @[Execute.scala 117:10]
  wire  _GEN_10058; // @[Execute.scala 117:10]
  wire  _GEN_10059; // @[Execute.scala 117:10]
  wire  _GEN_10060; // @[Execute.scala 117:10]
  wire  _GEN_10061; // @[Execute.scala 117:10]
  wire  _GEN_10062; // @[Execute.scala 117:10]
  wire  _GEN_10063; // @[Execute.scala 117:10]
  wire  _GEN_10064; // @[Execute.scala 117:10]
  wire  _GEN_10065; // @[Execute.scala 117:10]
  wire  _GEN_10066; // @[Execute.scala 117:10]
  wire  _GEN_10067; // @[Execute.scala 117:10]
  wire  _GEN_10068; // @[Execute.scala 117:10]
  wire  _GEN_10069; // @[Execute.scala 117:10]
  wire  _GEN_10070; // @[Execute.scala 117:10]
  wire  _GEN_10071; // @[Execute.scala 117:10]
  wire  _GEN_10072; // @[Execute.scala 117:10]
  wire  _GEN_10073; // @[Execute.scala 117:10]
  wire  _GEN_10074; // @[Execute.scala 117:10]
  wire  _GEN_10075; // @[Execute.scala 117:10]
  wire  _GEN_10076; // @[Execute.scala 117:10]
  wire  _GEN_10077; // @[Execute.scala 117:10]
  wire  _GEN_10078; // @[Execute.scala 117:10]
  wire  _GEN_10079; // @[Execute.scala 117:10]
  wire  _GEN_10080; // @[Execute.scala 117:10]
  wire  _GEN_10081; // @[Execute.scala 117:10]
  wire  _GEN_10082; // @[Execute.scala 117:10]
  wire  _GEN_10084; // @[Execute.scala 117:10]
  wire  _GEN_10085; // @[Execute.scala 117:10]
  wire  _GEN_10086; // @[Execute.scala 117:10]
  wire  _GEN_10087; // @[Execute.scala 117:10]
  wire  _GEN_10088; // @[Execute.scala 117:10]
  wire  _GEN_10089; // @[Execute.scala 117:10]
  wire  _GEN_10090; // @[Execute.scala 117:10]
  wire  _GEN_10091; // @[Execute.scala 117:10]
  wire  _GEN_10092; // @[Execute.scala 117:10]
  wire  _GEN_10093; // @[Execute.scala 117:10]
  wire  _GEN_10094; // @[Execute.scala 117:10]
  wire  _GEN_10095; // @[Execute.scala 117:10]
  wire  _GEN_10096; // @[Execute.scala 117:10]
  wire  _GEN_10097; // @[Execute.scala 117:10]
  wire  _GEN_10098; // @[Execute.scala 117:10]
  wire  _GEN_10099; // @[Execute.scala 117:10]
  wire  _GEN_10100; // @[Execute.scala 117:10]
  wire  _GEN_10101; // @[Execute.scala 117:10]
  wire  _GEN_10102; // @[Execute.scala 117:10]
  wire  _GEN_10103; // @[Execute.scala 117:10]
  wire  _GEN_10104; // @[Execute.scala 117:10]
  wire  _GEN_10105; // @[Execute.scala 117:10]
  wire  _GEN_10106; // @[Execute.scala 117:10]
  wire  _GEN_10107; // @[Execute.scala 117:10]
  wire  _GEN_10108; // @[Execute.scala 117:10]
  wire  _GEN_10109; // @[Execute.scala 117:10]
  wire  _GEN_10110; // @[Execute.scala 117:10]
  wire  _GEN_10111; // @[Execute.scala 117:10]
  wire  _GEN_10112; // @[Execute.scala 117:10]
  wire  _GEN_10113; // @[Execute.scala 117:10]
  wire  _GEN_10114; // @[Execute.scala 117:10]
  wire  _T_995; // @[Execute.scala 117:10]
  wire  _T_996; // @[Execute.scala 117:15]
  wire [4:0] _T_998; // @[Execute.scala 117:37]
  wire [4:0] _T_1000; // @[Execute.scala 117:60]
  wire  _GEN_10116; // @[Execute.scala 117:10]
  wire  _GEN_10117; // @[Execute.scala 117:10]
  wire  _GEN_10118; // @[Execute.scala 117:10]
  wire  _GEN_10119; // @[Execute.scala 117:10]
  wire  _GEN_10120; // @[Execute.scala 117:10]
  wire  _GEN_10121; // @[Execute.scala 117:10]
  wire  _GEN_10122; // @[Execute.scala 117:10]
  wire  _GEN_10123; // @[Execute.scala 117:10]
  wire  _GEN_10124; // @[Execute.scala 117:10]
  wire  _GEN_10125; // @[Execute.scala 117:10]
  wire  _GEN_10126; // @[Execute.scala 117:10]
  wire  _GEN_10127; // @[Execute.scala 117:10]
  wire  _GEN_10128; // @[Execute.scala 117:10]
  wire  _GEN_10129; // @[Execute.scala 117:10]
  wire  _GEN_10130; // @[Execute.scala 117:10]
  wire  _GEN_10131; // @[Execute.scala 117:10]
  wire  _GEN_10132; // @[Execute.scala 117:10]
  wire  _GEN_10133; // @[Execute.scala 117:10]
  wire  _GEN_10134; // @[Execute.scala 117:10]
  wire  _GEN_10135; // @[Execute.scala 117:10]
  wire  _GEN_10136; // @[Execute.scala 117:10]
  wire  _GEN_10137; // @[Execute.scala 117:10]
  wire  _GEN_10138; // @[Execute.scala 117:10]
  wire  _GEN_10139; // @[Execute.scala 117:10]
  wire  _GEN_10140; // @[Execute.scala 117:10]
  wire  _GEN_10141; // @[Execute.scala 117:10]
  wire  _GEN_10142; // @[Execute.scala 117:10]
  wire  _GEN_10143; // @[Execute.scala 117:10]
  wire  _GEN_10144; // @[Execute.scala 117:10]
  wire  _GEN_10145; // @[Execute.scala 117:10]
  wire  _GEN_10146; // @[Execute.scala 117:10]
  wire  _GEN_10148; // @[Execute.scala 117:10]
  wire  _GEN_10149; // @[Execute.scala 117:10]
  wire  _GEN_10150; // @[Execute.scala 117:10]
  wire  _GEN_10151; // @[Execute.scala 117:10]
  wire  _GEN_10152; // @[Execute.scala 117:10]
  wire  _GEN_10153; // @[Execute.scala 117:10]
  wire  _GEN_10154; // @[Execute.scala 117:10]
  wire  _GEN_10155; // @[Execute.scala 117:10]
  wire  _GEN_10156; // @[Execute.scala 117:10]
  wire  _GEN_10157; // @[Execute.scala 117:10]
  wire  _GEN_10158; // @[Execute.scala 117:10]
  wire  _GEN_10159; // @[Execute.scala 117:10]
  wire  _GEN_10160; // @[Execute.scala 117:10]
  wire  _GEN_10161; // @[Execute.scala 117:10]
  wire  _GEN_10162; // @[Execute.scala 117:10]
  wire  _GEN_10163; // @[Execute.scala 117:10]
  wire  _GEN_10164; // @[Execute.scala 117:10]
  wire  _GEN_10165; // @[Execute.scala 117:10]
  wire  _GEN_10166; // @[Execute.scala 117:10]
  wire  _GEN_10167; // @[Execute.scala 117:10]
  wire  _GEN_10168; // @[Execute.scala 117:10]
  wire  _GEN_10169; // @[Execute.scala 117:10]
  wire  _GEN_10170; // @[Execute.scala 117:10]
  wire  _GEN_10171; // @[Execute.scala 117:10]
  wire  _GEN_10172; // @[Execute.scala 117:10]
  wire  _GEN_10173; // @[Execute.scala 117:10]
  wire  _GEN_10174; // @[Execute.scala 117:10]
  wire  _GEN_10175; // @[Execute.scala 117:10]
  wire  _GEN_10176; // @[Execute.scala 117:10]
  wire  _GEN_10177; // @[Execute.scala 117:10]
  wire  _GEN_10178; // @[Execute.scala 117:10]
  wire  _T_1001; // @[Execute.scala 117:10]
  wire  _T_1002; // @[Execute.scala 117:15]
  wire [4:0] _T_1004; // @[Execute.scala 117:37]
  wire [4:0] _T_1006; // @[Execute.scala 117:60]
  wire  _GEN_10180; // @[Execute.scala 117:10]
  wire  _GEN_10181; // @[Execute.scala 117:10]
  wire  _GEN_10182; // @[Execute.scala 117:10]
  wire  _GEN_10183; // @[Execute.scala 117:10]
  wire  _GEN_10184; // @[Execute.scala 117:10]
  wire  _GEN_10185; // @[Execute.scala 117:10]
  wire  _GEN_10186; // @[Execute.scala 117:10]
  wire  _GEN_10187; // @[Execute.scala 117:10]
  wire  _GEN_10188; // @[Execute.scala 117:10]
  wire  _GEN_10189; // @[Execute.scala 117:10]
  wire  _GEN_10190; // @[Execute.scala 117:10]
  wire  _GEN_10191; // @[Execute.scala 117:10]
  wire  _GEN_10192; // @[Execute.scala 117:10]
  wire  _GEN_10193; // @[Execute.scala 117:10]
  wire  _GEN_10194; // @[Execute.scala 117:10]
  wire  _GEN_10195; // @[Execute.scala 117:10]
  wire  _GEN_10196; // @[Execute.scala 117:10]
  wire  _GEN_10197; // @[Execute.scala 117:10]
  wire  _GEN_10198; // @[Execute.scala 117:10]
  wire  _GEN_10199; // @[Execute.scala 117:10]
  wire  _GEN_10200; // @[Execute.scala 117:10]
  wire  _GEN_10201; // @[Execute.scala 117:10]
  wire  _GEN_10202; // @[Execute.scala 117:10]
  wire  _GEN_10203; // @[Execute.scala 117:10]
  wire  _GEN_10204; // @[Execute.scala 117:10]
  wire  _GEN_10205; // @[Execute.scala 117:10]
  wire  _GEN_10206; // @[Execute.scala 117:10]
  wire  _GEN_10207; // @[Execute.scala 117:10]
  wire  _GEN_10208; // @[Execute.scala 117:10]
  wire  _GEN_10209; // @[Execute.scala 117:10]
  wire  _GEN_10210; // @[Execute.scala 117:10]
  wire  _GEN_10212; // @[Execute.scala 117:10]
  wire  _GEN_10213; // @[Execute.scala 117:10]
  wire  _GEN_10214; // @[Execute.scala 117:10]
  wire  _GEN_10215; // @[Execute.scala 117:10]
  wire  _GEN_10216; // @[Execute.scala 117:10]
  wire  _GEN_10217; // @[Execute.scala 117:10]
  wire  _GEN_10218; // @[Execute.scala 117:10]
  wire  _GEN_10219; // @[Execute.scala 117:10]
  wire  _GEN_10220; // @[Execute.scala 117:10]
  wire  _GEN_10221; // @[Execute.scala 117:10]
  wire  _GEN_10222; // @[Execute.scala 117:10]
  wire  _GEN_10223; // @[Execute.scala 117:10]
  wire  _GEN_10224; // @[Execute.scala 117:10]
  wire  _GEN_10225; // @[Execute.scala 117:10]
  wire  _GEN_10226; // @[Execute.scala 117:10]
  wire  _GEN_10227; // @[Execute.scala 117:10]
  wire  _GEN_10228; // @[Execute.scala 117:10]
  wire  _GEN_10229; // @[Execute.scala 117:10]
  wire  _GEN_10230; // @[Execute.scala 117:10]
  wire  _GEN_10231; // @[Execute.scala 117:10]
  wire  _GEN_10232; // @[Execute.scala 117:10]
  wire  _GEN_10233; // @[Execute.scala 117:10]
  wire  _GEN_10234; // @[Execute.scala 117:10]
  wire  _GEN_10235; // @[Execute.scala 117:10]
  wire  _GEN_10236; // @[Execute.scala 117:10]
  wire  _GEN_10237; // @[Execute.scala 117:10]
  wire  _GEN_10238; // @[Execute.scala 117:10]
  wire  _GEN_10239; // @[Execute.scala 117:10]
  wire  _GEN_10240; // @[Execute.scala 117:10]
  wire  _GEN_10241; // @[Execute.scala 117:10]
  wire  _GEN_10242; // @[Execute.scala 117:10]
  wire  _T_1007; // @[Execute.scala 117:10]
  wire  _T_1008; // @[Execute.scala 117:15]
  wire [4:0] _T_1010; // @[Execute.scala 117:37]
  wire [4:0] _T_1012; // @[Execute.scala 117:60]
  wire  _GEN_10244; // @[Execute.scala 117:10]
  wire  _GEN_10245; // @[Execute.scala 117:10]
  wire  _GEN_10246; // @[Execute.scala 117:10]
  wire  _GEN_10247; // @[Execute.scala 117:10]
  wire  _GEN_10248; // @[Execute.scala 117:10]
  wire  _GEN_10249; // @[Execute.scala 117:10]
  wire  _GEN_10250; // @[Execute.scala 117:10]
  wire  _GEN_10251; // @[Execute.scala 117:10]
  wire  _GEN_10252; // @[Execute.scala 117:10]
  wire  _GEN_10253; // @[Execute.scala 117:10]
  wire  _GEN_10254; // @[Execute.scala 117:10]
  wire  _GEN_10255; // @[Execute.scala 117:10]
  wire  _GEN_10256; // @[Execute.scala 117:10]
  wire  _GEN_10257; // @[Execute.scala 117:10]
  wire  _GEN_10258; // @[Execute.scala 117:10]
  wire  _GEN_10259; // @[Execute.scala 117:10]
  wire  _GEN_10260; // @[Execute.scala 117:10]
  wire  _GEN_10261; // @[Execute.scala 117:10]
  wire  _GEN_10262; // @[Execute.scala 117:10]
  wire  _GEN_10263; // @[Execute.scala 117:10]
  wire  _GEN_10264; // @[Execute.scala 117:10]
  wire  _GEN_10265; // @[Execute.scala 117:10]
  wire  _GEN_10266; // @[Execute.scala 117:10]
  wire  _GEN_10267; // @[Execute.scala 117:10]
  wire  _GEN_10268; // @[Execute.scala 117:10]
  wire  _GEN_10269; // @[Execute.scala 117:10]
  wire  _GEN_10270; // @[Execute.scala 117:10]
  wire  _GEN_10271; // @[Execute.scala 117:10]
  wire  _GEN_10272; // @[Execute.scala 117:10]
  wire  _GEN_10273; // @[Execute.scala 117:10]
  wire  _GEN_10274; // @[Execute.scala 117:10]
  wire  _GEN_10276; // @[Execute.scala 117:10]
  wire  _GEN_10277; // @[Execute.scala 117:10]
  wire  _GEN_10278; // @[Execute.scala 117:10]
  wire  _GEN_10279; // @[Execute.scala 117:10]
  wire  _GEN_10280; // @[Execute.scala 117:10]
  wire  _GEN_10281; // @[Execute.scala 117:10]
  wire  _GEN_10282; // @[Execute.scala 117:10]
  wire  _GEN_10283; // @[Execute.scala 117:10]
  wire  _GEN_10284; // @[Execute.scala 117:10]
  wire  _GEN_10285; // @[Execute.scala 117:10]
  wire  _GEN_10286; // @[Execute.scala 117:10]
  wire  _GEN_10287; // @[Execute.scala 117:10]
  wire  _GEN_10288; // @[Execute.scala 117:10]
  wire  _GEN_10289; // @[Execute.scala 117:10]
  wire  _GEN_10290; // @[Execute.scala 117:10]
  wire  _GEN_10291; // @[Execute.scala 117:10]
  wire  _GEN_10292; // @[Execute.scala 117:10]
  wire  _GEN_10293; // @[Execute.scala 117:10]
  wire  _GEN_10294; // @[Execute.scala 117:10]
  wire  _GEN_10295; // @[Execute.scala 117:10]
  wire  _GEN_10296; // @[Execute.scala 117:10]
  wire  _GEN_10297; // @[Execute.scala 117:10]
  wire  _GEN_10298; // @[Execute.scala 117:10]
  wire  _GEN_10299; // @[Execute.scala 117:10]
  wire  _GEN_10300; // @[Execute.scala 117:10]
  wire  _GEN_10301; // @[Execute.scala 117:10]
  wire  _GEN_10302; // @[Execute.scala 117:10]
  wire  _GEN_10303; // @[Execute.scala 117:10]
  wire  _GEN_10304; // @[Execute.scala 117:10]
  wire  _GEN_10305; // @[Execute.scala 117:10]
  wire  _GEN_10306; // @[Execute.scala 117:10]
  wire  _T_1013; // @[Execute.scala 117:10]
  wire  _T_1014; // @[Execute.scala 117:15]
  wire [4:0] _T_1016; // @[Execute.scala 117:37]
  wire [4:0] _T_1018; // @[Execute.scala 117:60]
  wire  _GEN_10308; // @[Execute.scala 117:10]
  wire  _GEN_10309; // @[Execute.scala 117:10]
  wire  _GEN_10310; // @[Execute.scala 117:10]
  wire  _GEN_10311; // @[Execute.scala 117:10]
  wire  _GEN_10312; // @[Execute.scala 117:10]
  wire  _GEN_10313; // @[Execute.scala 117:10]
  wire  _GEN_10314; // @[Execute.scala 117:10]
  wire  _GEN_10315; // @[Execute.scala 117:10]
  wire  _GEN_10316; // @[Execute.scala 117:10]
  wire  _GEN_10317; // @[Execute.scala 117:10]
  wire  _GEN_10318; // @[Execute.scala 117:10]
  wire  _GEN_10319; // @[Execute.scala 117:10]
  wire  _GEN_10320; // @[Execute.scala 117:10]
  wire  _GEN_10321; // @[Execute.scala 117:10]
  wire  _GEN_10322; // @[Execute.scala 117:10]
  wire  _GEN_10323; // @[Execute.scala 117:10]
  wire  _GEN_10324; // @[Execute.scala 117:10]
  wire  _GEN_10325; // @[Execute.scala 117:10]
  wire  _GEN_10326; // @[Execute.scala 117:10]
  wire  _GEN_10327; // @[Execute.scala 117:10]
  wire  _GEN_10328; // @[Execute.scala 117:10]
  wire  _GEN_10329; // @[Execute.scala 117:10]
  wire  _GEN_10330; // @[Execute.scala 117:10]
  wire  _GEN_10331; // @[Execute.scala 117:10]
  wire  _GEN_10332; // @[Execute.scala 117:10]
  wire  _GEN_10333; // @[Execute.scala 117:10]
  wire  _GEN_10334; // @[Execute.scala 117:10]
  wire  _GEN_10335; // @[Execute.scala 117:10]
  wire  _GEN_10336; // @[Execute.scala 117:10]
  wire  _GEN_10337; // @[Execute.scala 117:10]
  wire  _GEN_10338; // @[Execute.scala 117:10]
  wire  _GEN_10340; // @[Execute.scala 117:10]
  wire  _GEN_10341; // @[Execute.scala 117:10]
  wire  _GEN_10342; // @[Execute.scala 117:10]
  wire  _GEN_10343; // @[Execute.scala 117:10]
  wire  _GEN_10344; // @[Execute.scala 117:10]
  wire  _GEN_10345; // @[Execute.scala 117:10]
  wire  _GEN_10346; // @[Execute.scala 117:10]
  wire  _GEN_10347; // @[Execute.scala 117:10]
  wire  _GEN_10348; // @[Execute.scala 117:10]
  wire  _GEN_10349; // @[Execute.scala 117:10]
  wire  _GEN_10350; // @[Execute.scala 117:10]
  wire  _GEN_10351; // @[Execute.scala 117:10]
  wire  _GEN_10352; // @[Execute.scala 117:10]
  wire  _GEN_10353; // @[Execute.scala 117:10]
  wire  _GEN_10354; // @[Execute.scala 117:10]
  wire  _GEN_10355; // @[Execute.scala 117:10]
  wire  _GEN_10356; // @[Execute.scala 117:10]
  wire  _GEN_10357; // @[Execute.scala 117:10]
  wire  _GEN_10358; // @[Execute.scala 117:10]
  wire  _GEN_10359; // @[Execute.scala 117:10]
  wire  _GEN_10360; // @[Execute.scala 117:10]
  wire  _GEN_10361; // @[Execute.scala 117:10]
  wire  _GEN_10362; // @[Execute.scala 117:10]
  wire  _GEN_10363; // @[Execute.scala 117:10]
  wire  _GEN_10364; // @[Execute.scala 117:10]
  wire  _GEN_10365; // @[Execute.scala 117:10]
  wire  _GEN_10366; // @[Execute.scala 117:10]
  wire  _GEN_10367; // @[Execute.scala 117:10]
  wire  _GEN_10368; // @[Execute.scala 117:10]
  wire  _GEN_10369; // @[Execute.scala 117:10]
  wire  _GEN_10370; // @[Execute.scala 117:10]
  wire  _T_1019; // @[Execute.scala 117:10]
  wire  _T_1020; // @[Execute.scala 117:15]
  wire [4:0] _T_1022; // @[Execute.scala 117:37]
  wire [4:0] _T_1024; // @[Execute.scala 117:60]
  wire  _GEN_10372; // @[Execute.scala 117:10]
  wire  _GEN_10373; // @[Execute.scala 117:10]
  wire  _GEN_10374; // @[Execute.scala 117:10]
  wire  _GEN_10375; // @[Execute.scala 117:10]
  wire  _GEN_10376; // @[Execute.scala 117:10]
  wire  _GEN_10377; // @[Execute.scala 117:10]
  wire  _GEN_10378; // @[Execute.scala 117:10]
  wire  _GEN_10379; // @[Execute.scala 117:10]
  wire  _GEN_10380; // @[Execute.scala 117:10]
  wire  _GEN_10381; // @[Execute.scala 117:10]
  wire  _GEN_10382; // @[Execute.scala 117:10]
  wire  _GEN_10383; // @[Execute.scala 117:10]
  wire  _GEN_10384; // @[Execute.scala 117:10]
  wire  _GEN_10385; // @[Execute.scala 117:10]
  wire  _GEN_10386; // @[Execute.scala 117:10]
  wire  _GEN_10387; // @[Execute.scala 117:10]
  wire  _GEN_10388; // @[Execute.scala 117:10]
  wire  _GEN_10389; // @[Execute.scala 117:10]
  wire  _GEN_10390; // @[Execute.scala 117:10]
  wire  _GEN_10391; // @[Execute.scala 117:10]
  wire  _GEN_10392; // @[Execute.scala 117:10]
  wire  _GEN_10393; // @[Execute.scala 117:10]
  wire  _GEN_10394; // @[Execute.scala 117:10]
  wire  _GEN_10395; // @[Execute.scala 117:10]
  wire  _GEN_10396; // @[Execute.scala 117:10]
  wire  _GEN_10397; // @[Execute.scala 117:10]
  wire  _GEN_10398; // @[Execute.scala 117:10]
  wire  _GEN_10399; // @[Execute.scala 117:10]
  wire  _GEN_10400; // @[Execute.scala 117:10]
  wire  _GEN_10401; // @[Execute.scala 117:10]
  wire  _GEN_10402; // @[Execute.scala 117:10]
  wire  _GEN_10404; // @[Execute.scala 117:10]
  wire  _GEN_10405; // @[Execute.scala 117:10]
  wire  _GEN_10406; // @[Execute.scala 117:10]
  wire  _GEN_10407; // @[Execute.scala 117:10]
  wire  _GEN_10408; // @[Execute.scala 117:10]
  wire  _GEN_10409; // @[Execute.scala 117:10]
  wire  _GEN_10410; // @[Execute.scala 117:10]
  wire  _GEN_10411; // @[Execute.scala 117:10]
  wire  _GEN_10412; // @[Execute.scala 117:10]
  wire  _GEN_10413; // @[Execute.scala 117:10]
  wire  _GEN_10414; // @[Execute.scala 117:10]
  wire  _GEN_10415; // @[Execute.scala 117:10]
  wire  _GEN_10416; // @[Execute.scala 117:10]
  wire  _GEN_10417; // @[Execute.scala 117:10]
  wire  _GEN_10418; // @[Execute.scala 117:10]
  wire  _GEN_10419; // @[Execute.scala 117:10]
  wire  _GEN_10420; // @[Execute.scala 117:10]
  wire  _GEN_10421; // @[Execute.scala 117:10]
  wire  _GEN_10422; // @[Execute.scala 117:10]
  wire  _GEN_10423; // @[Execute.scala 117:10]
  wire  _GEN_10424; // @[Execute.scala 117:10]
  wire  _GEN_10425; // @[Execute.scala 117:10]
  wire  _GEN_10426; // @[Execute.scala 117:10]
  wire  _GEN_10427; // @[Execute.scala 117:10]
  wire  _GEN_10428; // @[Execute.scala 117:10]
  wire  _GEN_10429; // @[Execute.scala 117:10]
  wire  _GEN_10430; // @[Execute.scala 117:10]
  wire  _GEN_10431; // @[Execute.scala 117:10]
  wire  _GEN_10432; // @[Execute.scala 117:10]
  wire  _GEN_10433; // @[Execute.scala 117:10]
  wire  _GEN_10434; // @[Execute.scala 117:10]
  wire  _T_1025; // @[Execute.scala 117:10]
  wire [7:0] _T_1033; // @[Execute.scala 311:68]
  wire [15:0] _T_1041; // @[Execute.scala 311:68]
  wire [7:0] _T_1048; // @[Execute.scala 311:68]
  wire [31:0] _T_1057; // @[Execute.scala 311:68]
  wire [63:0] _T_1058; // @[Execute.scala 311:78]
  assign _T = ~io_imms; // @[Execute.scala 289:54]
  assign toBeEncoded = {io_immn,_T}; // @[Cat.scala 29:58]
  assign _T_10 = toBeEncoded[2] ? 2'h2 : {{1'd0}, toBeEncoded[1]}; // @[Mux.scala 47:69]
  assign _T_11 = toBeEncoded[3] ? 2'h3 : _T_10; // @[Mux.scala 47:69]
  assign _T_12 = toBeEncoded[4] ? 3'h4 : {{1'd0}, _T_11}; // @[Mux.scala 47:69]
  assign _T_13 = toBeEncoded[5] ? 3'h5 : _T_12; // @[Mux.scala 47:69]
  assign len = toBeEncoded[6] ? 3'h6 : _T_13; // @[Mux.scala 47:69]
  assign _T_15 = {{4'd0}, len};
  assign _GEN_1 = 7'h1 == _T_15 ? 64'h1 : 64'h0; // @[Execute.scala 291:39]
  assign _GEN_2 = 7'h2 == _T_15 ? 64'h3 : _GEN_1; // @[Execute.scala 291:39]
  assign _GEN_3 = 7'h3 == _T_15 ? 64'h7 : _GEN_2; // @[Execute.scala 291:39]
  assign _GEN_4 = 7'h4 == _T_15 ? 64'hf : _GEN_3; // @[Execute.scala 291:39]
  assign _GEN_5 = 7'h5 == _T_15 ? 64'h1f : _GEN_4; // @[Execute.scala 291:39]
  assign _GEN_6 = 7'h6 == _T_15 ? 64'h3f : _GEN_5; // @[Execute.scala 291:39]
  assign _GEN_7 = 7'h7 == _T_15 ? 64'h7f : _GEN_6; // @[Execute.scala 291:39]
  assign _GEN_8 = 7'h8 == _T_15 ? 64'hff : _GEN_7; // @[Execute.scala 291:39]
  assign _GEN_9 = 7'h9 == _T_15 ? 64'h1ff : _GEN_8; // @[Execute.scala 291:39]
  assign _GEN_10 = 7'ha == _T_15 ? 64'h3ff : _GEN_9; // @[Execute.scala 291:39]
  assign _GEN_11 = 7'hb == _T_15 ? 64'h7ff : _GEN_10; // @[Execute.scala 291:39]
  assign _GEN_12 = 7'hc == _T_15 ? 64'hfff : _GEN_11; // @[Execute.scala 291:39]
  assign _GEN_13 = 7'hd == _T_15 ? 64'h1fff : _GEN_12; // @[Execute.scala 291:39]
  assign _GEN_14 = 7'he == _T_15 ? 64'h3fff : _GEN_13; // @[Execute.scala 291:39]
  assign _GEN_15 = 7'hf == _T_15 ? 64'h7fff : _GEN_14; // @[Execute.scala 291:39]
  assign _GEN_16 = 7'h10 == _T_15 ? 64'hffff : _GEN_15; // @[Execute.scala 291:39]
  assign _GEN_17 = 7'h11 == _T_15 ? 64'h1ffff : _GEN_16; // @[Execute.scala 291:39]
  assign _GEN_18 = 7'h12 == _T_15 ? 64'h3ffff : _GEN_17; // @[Execute.scala 291:39]
  assign _GEN_19 = 7'h13 == _T_15 ? 64'h7ffff : _GEN_18; // @[Execute.scala 291:39]
  assign _GEN_20 = 7'h14 == _T_15 ? 64'hfffff : _GEN_19; // @[Execute.scala 291:39]
  assign _GEN_21 = 7'h15 == _T_15 ? 64'h1fffff : _GEN_20; // @[Execute.scala 291:39]
  assign _GEN_22 = 7'h16 == _T_15 ? 64'h3fffff : _GEN_21; // @[Execute.scala 291:39]
  assign _GEN_23 = 7'h17 == _T_15 ? 64'h7fffff : _GEN_22; // @[Execute.scala 291:39]
  assign _GEN_24 = 7'h18 == _T_15 ? 64'hffffff : _GEN_23; // @[Execute.scala 291:39]
  assign _GEN_25 = 7'h19 == _T_15 ? 64'h1ffffff : _GEN_24; // @[Execute.scala 291:39]
  assign _GEN_26 = 7'h1a == _T_15 ? 64'h3ffffff : _GEN_25; // @[Execute.scala 291:39]
  assign _GEN_27 = 7'h1b == _T_15 ? 64'h7ffffff : _GEN_26; // @[Execute.scala 291:39]
  assign _GEN_28 = 7'h1c == _T_15 ? 64'hfffffff : _GEN_27; // @[Execute.scala 291:39]
  assign _GEN_29 = 7'h1d == _T_15 ? 64'h1fffffff : _GEN_28; // @[Execute.scala 291:39]
  assign _GEN_30 = 7'h1e == _T_15 ? 64'h3fffffff : _GEN_29; // @[Execute.scala 291:39]
  assign _GEN_31 = 7'h1f == _T_15 ? 64'h7fffffff : _GEN_30; // @[Execute.scala 291:39]
  assign _GEN_32 = 7'h20 == _T_15 ? 64'hffffffff : _GEN_31; // @[Execute.scala 291:39]
  assign _GEN_33 = 7'h21 == _T_15 ? 64'h1ffffffff : _GEN_32; // @[Execute.scala 291:39]
  assign _GEN_34 = 7'h22 == _T_15 ? 64'h3ffffffff : _GEN_33; // @[Execute.scala 291:39]
  assign _GEN_35 = 7'h23 == _T_15 ? 64'h7ffffffff : _GEN_34; // @[Execute.scala 291:39]
  assign _GEN_36 = 7'h24 == _T_15 ? 64'hfffffffff : _GEN_35; // @[Execute.scala 291:39]
  assign _GEN_37 = 7'h25 == _T_15 ? 64'h1fffffffff : _GEN_36; // @[Execute.scala 291:39]
  assign _GEN_38 = 7'h26 == _T_15 ? 64'h3fffffffff : _GEN_37; // @[Execute.scala 291:39]
  assign _GEN_39 = 7'h27 == _T_15 ? 64'h7fffffffff : _GEN_38; // @[Execute.scala 291:39]
  assign _GEN_40 = 7'h28 == _T_15 ? 64'hffffffffff : _GEN_39; // @[Execute.scala 291:39]
  assign _GEN_41 = 7'h29 == _T_15 ? 64'h1ffffffffff : _GEN_40; // @[Execute.scala 291:39]
  assign _GEN_42 = 7'h2a == _T_15 ? 64'h3ffffffffff : _GEN_41; // @[Execute.scala 291:39]
  assign _GEN_43 = 7'h2b == _T_15 ? 64'h7ffffffffff : _GEN_42; // @[Execute.scala 291:39]
  assign _GEN_44 = 7'h2c == _T_15 ? 64'hfffffffffff : _GEN_43; // @[Execute.scala 291:39]
  assign _GEN_45 = 7'h2d == _T_15 ? 64'h1fffffffffff : _GEN_44; // @[Execute.scala 291:39]
  assign _GEN_46 = 7'h2e == _T_15 ? 64'h3fffffffffff : _GEN_45; // @[Execute.scala 291:39]
  assign _GEN_47 = 7'h2f == _T_15 ? 64'h7fffffffffff : _GEN_46; // @[Execute.scala 291:39]
  assign _GEN_48 = 7'h30 == _T_15 ? 64'hffffffffffff : _GEN_47; // @[Execute.scala 291:39]
  assign _GEN_49 = 7'h31 == _T_15 ? 64'h1ffffffffffff : _GEN_48; // @[Execute.scala 291:39]
  assign _GEN_50 = 7'h32 == _T_15 ? 64'h3ffffffffffff : _GEN_49; // @[Execute.scala 291:39]
  assign _GEN_51 = 7'h33 == _T_15 ? 64'h7ffffffffffff : _GEN_50; // @[Execute.scala 291:39]
  assign _GEN_52 = 7'h34 == _T_15 ? 64'hfffffffffffff : _GEN_51; // @[Execute.scala 291:39]
  assign _GEN_53 = 7'h35 == _T_15 ? 64'h1fffffffffffff : _GEN_52; // @[Execute.scala 291:39]
  assign _GEN_54 = 7'h36 == _T_15 ? 64'h3fffffffffffff : _GEN_53; // @[Execute.scala 291:39]
  assign _GEN_55 = 7'h37 == _T_15 ? 64'h7fffffffffffff : _GEN_54; // @[Execute.scala 291:39]
  assign _GEN_56 = 7'h38 == _T_15 ? 64'hffffffffffffff : _GEN_55; // @[Execute.scala 291:39]
  assign _GEN_57 = 7'h39 == _T_15 ? 64'h1ffffffffffffff : _GEN_56; // @[Execute.scala 291:39]
  assign _GEN_58 = 7'h3a == _T_15 ? 64'h3ffffffffffffff : _GEN_57; // @[Execute.scala 291:39]
  assign _GEN_59 = 7'h3b == _T_15 ? 64'h7ffffffffffffff : _GEN_58; // @[Execute.scala 291:39]
  assign _GEN_60 = 7'h3c == _T_15 ? 64'hfffffffffffffff : _GEN_59; // @[Execute.scala 291:39]
  assign _GEN_61 = 7'h3d == _T_15 ? 64'h1fffffffffffffff : _GEN_60; // @[Execute.scala 291:39]
  assign _GEN_62 = 7'h3e == _T_15 ? 64'h3fffffffffffffff : _GEN_61; // @[Execute.scala 291:39]
  assign _GEN_63 = 7'h3f == _T_15 ? 64'h7fffffffffffffff : _GEN_62; // @[Execute.scala 291:39]
  assign _GEN_64 = 7'h40 == _T_15 ? 64'hffffffffffffffff : _GEN_63; // @[Execute.scala 291:39]
  assign levels = _GEN_64[5:0]; // @[Execute.scala 291:39]
  assign s = io_imms & levels; // @[Execute.scala 293:28]
  assign r = io_immr & levels; // @[Execute.scala 294:28]
  assign diff = s - r; // @[Execute.scala 295:25]
  assign _GEN_10436 = {{1'd0}, levels}; // @[Execute.scala 297:25]
  assign d = diff & _GEN_10436; // @[Execute.scala 297:25]
  assign onesS = s + 6'h1; // @[Execute.scala 298:26]
  assign onesD = d + 7'h1; // @[Execute.scala 299:26]
  assign _GEN_66 = 7'h1 == onesS ? 64'h1 : 64'h0; // @[Execute.scala 301:9]
  assign _GEN_67 = 7'h2 == onesS ? 64'h3 : _GEN_66; // @[Execute.scala 301:9]
  assign _GEN_68 = 7'h3 == onesS ? 64'h7 : _GEN_67; // @[Execute.scala 301:9]
  assign _GEN_69 = 7'h4 == onesS ? 64'hf : _GEN_68; // @[Execute.scala 301:9]
  assign _GEN_70 = 7'h5 == onesS ? 64'h1f : _GEN_69; // @[Execute.scala 301:9]
  assign _GEN_71 = 7'h6 == onesS ? 64'h3f : _GEN_70; // @[Execute.scala 301:9]
  assign _GEN_72 = 7'h7 == onesS ? 64'h7f : _GEN_71; // @[Execute.scala 301:9]
  assign _GEN_73 = 7'h8 == onesS ? 64'hff : _GEN_72; // @[Execute.scala 301:9]
  assign _GEN_74 = 7'h9 == onesS ? 64'h1ff : _GEN_73; // @[Execute.scala 301:9]
  assign _GEN_75 = 7'ha == onesS ? 64'h3ff : _GEN_74; // @[Execute.scala 301:9]
  assign _GEN_76 = 7'hb == onesS ? 64'h7ff : _GEN_75; // @[Execute.scala 301:9]
  assign _GEN_77 = 7'hc == onesS ? 64'hfff : _GEN_76; // @[Execute.scala 301:9]
  assign _GEN_78 = 7'hd == onesS ? 64'h1fff : _GEN_77; // @[Execute.scala 301:9]
  assign _GEN_79 = 7'he == onesS ? 64'h3fff : _GEN_78; // @[Execute.scala 301:9]
  assign _GEN_80 = 7'hf == onesS ? 64'h7fff : _GEN_79; // @[Execute.scala 301:9]
  assign _GEN_81 = 7'h10 == onesS ? 64'hffff : _GEN_80; // @[Execute.scala 301:9]
  assign _GEN_82 = 7'h11 == onesS ? 64'h1ffff : _GEN_81; // @[Execute.scala 301:9]
  assign _GEN_83 = 7'h12 == onesS ? 64'h3ffff : _GEN_82; // @[Execute.scala 301:9]
  assign _GEN_84 = 7'h13 == onesS ? 64'h7ffff : _GEN_83; // @[Execute.scala 301:9]
  assign _GEN_85 = 7'h14 == onesS ? 64'hfffff : _GEN_84; // @[Execute.scala 301:9]
  assign _GEN_86 = 7'h15 == onesS ? 64'h1fffff : _GEN_85; // @[Execute.scala 301:9]
  assign _GEN_87 = 7'h16 == onesS ? 64'h3fffff : _GEN_86; // @[Execute.scala 301:9]
  assign _GEN_88 = 7'h17 == onesS ? 64'h7fffff : _GEN_87; // @[Execute.scala 301:9]
  assign _GEN_89 = 7'h18 == onesS ? 64'hffffff : _GEN_88; // @[Execute.scala 301:9]
  assign _GEN_90 = 7'h19 == onesS ? 64'h1ffffff : _GEN_89; // @[Execute.scala 301:9]
  assign _GEN_91 = 7'h1a == onesS ? 64'h3ffffff : _GEN_90; // @[Execute.scala 301:9]
  assign _GEN_92 = 7'h1b == onesS ? 64'h7ffffff : _GEN_91; // @[Execute.scala 301:9]
  assign _GEN_93 = 7'h1c == onesS ? 64'hfffffff : _GEN_92; // @[Execute.scala 301:9]
  assign _GEN_94 = 7'h1d == onesS ? 64'h1fffffff : _GEN_93; // @[Execute.scala 301:9]
  assign _GEN_95 = 7'h1e == onesS ? 64'h3fffffff : _GEN_94; // @[Execute.scala 301:9]
  assign _GEN_96 = 7'h1f == onesS ? 64'h7fffffff : _GEN_95; // @[Execute.scala 301:9]
  assign _GEN_97 = 7'h20 == onesS ? 64'hffffffff : _GEN_96; // @[Execute.scala 301:9]
  assign _GEN_98 = 7'h21 == onesS ? 64'h1ffffffff : _GEN_97; // @[Execute.scala 301:9]
  assign _GEN_99 = 7'h22 == onesS ? 64'h3ffffffff : _GEN_98; // @[Execute.scala 301:9]
  assign _GEN_100 = 7'h23 == onesS ? 64'h7ffffffff : _GEN_99; // @[Execute.scala 301:9]
  assign _GEN_101 = 7'h24 == onesS ? 64'hfffffffff : _GEN_100; // @[Execute.scala 301:9]
  assign _GEN_102 = 7'h25 == onesS ? 64'h1fffffffff : _GEN_101; // @[Execute.scala 301:9]
  assign _GEN_103 = 7'h26 == onesS ? 64'h3fffffffff : _GEN_102; // @[Execute.scala 301:9]
  assign _GEN_104 = 7'h27 == onesS ? 64'h7fffffffff : _GEN_103; // @[Execute.scala 301:9]
  assign _GEN_105 = 7'h28 == onesS ? 64'hffffffffff : _GEN_104; // @[Execute.scala 301:9]
  assign _GEN_106 = 7'h29 == onesS ? 64'h1ffffffffff : _GEN_105; // @[Execute.scala 301:9]
  assign _GEN_107 = 7'h2a == onesS ? 64'h3ffffffffff : _GEN_106; // @[Execute.scala 301:9]
  assign _GEN_108 = 7'h2b == onesS ? 64'h7ffffffffff : _GEN_107; // @[Execute.scala 301:9]
  assign _GEN_109 = 7'h2c == onesS ? 64'hfffffffffff : _GEN_108; // @[Execute.scala 301:9]
  assign _GEN_110 = 7'h2d == onesS ? 64'h1fffffffffff : _GEN_109; // @[Execute.scala 301:9]
  assign _GEN_111 = 7'h2e == onesS ? 64'h3fffffffffff : _GEN_110; // @[Execute.scala 301:9]
  assign _GEN_112 = 7'h2f == onesS ? 64'h7fffffffffff : _GEN_111; // @[Execute.scala 301:9]
  assign _GEN_113 = 7'h30 == onesS ? 64'hffffffffffff : _GEN_112; // @[Execute.scala 301:9]
  assign _GEN_114 = 7'h31 == onesS ? 64'h1ffffffffffff : _GEN_113; // @[Execute.scala 301:9]
  assign _GEN_115 = 7'h32 == onesS ? 64'h3ffffffffffff : _GEN_114; // @[Execute.scala 301:9]
  assign _GEN_116 = 7'h33 == onesS ? 64'h7ffffffffffff : _GEN_115; // @[Execute.scala 301:9]
  assign _GEN_117 = 7'h34 == onesS ? 64'hfffffffffffff : _GEN_116; // @[Execute.scala 301:9]
  assign _GEN_118 = 7'h35 == onesS ? 64'h1fffffffffffff : _GEN_117; // @[Execute.scala 301:9]
  assign _GEN_119 = 7'h36 == onesS ? 64'h3fffffffffffff : _GEN_118; // @[Execute.scala 301:9]
  assign _GEN_120 = 7'h37 == onesS ? 64'h7fffffffffffff : _GEN_119; // @[Execute.scala 301:9]
  assign _GEN_121 = 7'h38 == onesS ? 64'hffffffffffffff : _GEN_120; // @[Execute.scala 301:9]
  assign _GEN_122 = 7'h39 == onesS ? 64'h1ffffffffffffff : _GEN_121; // @[Execute.scala 301:9]
  assign _GEN_123 = 7'h3a == onesS ? 64'h3ffffffffffffff : _GEN_122; // @[Execute.scala 301:9]
  assign _GEN_124 = 7'h3b == onesS ? 64'h7ffffffffffffff : _GEN_123; // @[Execute.scala 301:9]
  assign _GEN_125 = 7'h3c == onesS ? 64'hfffffffffffffff : _GEN_124; // @[Execute.scala 301:9]
  assign _GEN_126 = 7'h3d == onesS ? 64'h1fffffffffffffff : _GEN_125; // @[Execute.scala 301:9]
  assign _GEN_127 = 7'h3e == onesS ? 64'h3fffffffffffffff : _GEN_126; // @[Execute.scala 301:9]
  assign _GEN_128 = 7'h3f == onesS ? 64'h7fffffffffffffff : _GEN_127; // @[Execute.scala 301:9]
  assign welem = 7'h40 == onesS ? 64'hffffffffffffffff : _GEN_128; // @[Execute.scala 301:9]
  assign _GEN_10437 = {{1'd0}, r}; // @[Execute.scala 117:37]
  assign _T_94 = _GEN_10437 - 7'h40; // @[Execute.scala 117:37]
  assign _GEN_131 = 6'h1 == _T_94[5:0] ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_132 = 6'h2 == _T_94[5:0] ? welem[2] : _GEN_131; // @[Execute.scala 117:10]
  assign _GEN_133 = 6'h3 == _T_94[5:0] ? welem[3] : _GEN_132; // @[Execute.scala 117:10]
  assign _GEN_134 = 6'h4 == _T_94[5:0] ? welem[4] : _GEN_133; // @[Execute.scala 117:10]
  assign _GEN_135 = 6'h5 == _T_94[5:0] ? welem[5] : _GEN_134; // @[Execute.scala 117:10]
  assign _GEN_136 = 6'h6 == _T_94[5:0] ? welem[6] : _GEN_135; // @[Execute.scala 117:10]
  assign _GEN_137 = 6'h7 == _T_94[5:0] ? welem[7] : _GEN_136; // @[Execute.scala 117:10]
  assign _GEN_138 = 6'h8 == _T_94[5:0] ? welem[8] : _GEN_137; // @[Execute.scala 117:10]
  assign _GEN_139 = 6'h9 == _T_94[5:0] ? welem[9] : _GEN_138; // @[Execute.scala 117:10]
  assign _GEN_140 = 6'ha == _T_94[5:0] ? welem[10] : _GEN_139; // @[Execute.scala 117:10]
  assign _GEN_141 = 6'hb == _T_94[5:0] ? welem[11] : _GEN_140; // @[Execute.scala 117:10]
  assign _GEN_142 = 6'hc == _T_94[5:0] ? welem[12] : _GEN_141; // @[Execute.scala 117:10]
  assign _GEN_143 = 6'hd == _T_94[5:0] ? welem[13] : _GEN_142; // @[Execute.scala 117:10]
  assign _GEN_144 = 6'he == _T_94[5:0] ? welem[14] : _GEN_143; // @[Execute.scala 117:10]
  assign _GEN_145 = 6'hf == _T_94[5:0] ? welem[15] : _GEN_144; // @[Execute.scala 117:10]
  assign _GEN_146 = 6'h10 == _T_94[5:0] ? welem[16] : _GEN_145; // @[Execute.scala 117:10]
  assign _GEN_147 = 6'h11 == _T_94[5:0] ? welem[17] : _GEN_146; // @[Execute.scala 117:10]
  assign _GEN_148 = 6'h12 == _T_94[5:0] ? welem[18] : _GEN_147; // @[Execute.scala 117:10]
  assign _GEN_149 = 6'h13 == _T_94[5:0] ? welem[19] : _GEN_148; // @[Execute.scala 117:10]
  assign _GEN_150 = 6'h14 == _T_94[5:0] ? welem[20] : _GEN_149; // @[Execute.scala 117:10]
  assign _GEN_151 = 6'h15 == _T_94[5:0] ? welem[21] : _GEN_150; // @[Execute.scala 117:10]
  assign _GEN_152 = 6'h16 == _T_94[5:0] ? welem[22] : _GEN_151; // @[Execute.scala 117:10]
  assign _GEN_153 = 6'h17 == _T_94[5:0] ? welem[23] : _GEN_152; // @[Execute.scala 117:10]
  assign _GEN_154 = 6'h18 == _T_94[5:0] ? welem[24] : _GEN_153; // @[Execute.scala 117:10]
  assign _GEN_155 = 6'h19 == _T_94[5:0] ? welem[25] : _GEN_154; // @[Execute.scala 117:10]
  assign _GEN_156 = 6'h1a == _T_94[5:0] ? welem[26] : _GEN_155; // @[Execute.scala 117:10]
  assign _GEN_157 = 6'h1b == _T_94[5:0] ? welem[27] : _GEN_156; // @[Execute.scala 117:10]
  assign _GEN_158 = 6'h1c == _T_94[5:0] ? welem[28] : _GEN_157; // @[Execute.scala 117:10]
  assign _GEN_159 = 6'h1d == _T_94[5:0] ? welem[29] : _GEN_158; // @[Execute.scala 117:10]
  assign _GEN_160 = 6'h1e == _T_94[5:0] ? welem[30] : _GEN_159; // @[Execute.scala 117:10]
  assign _GEN_161 = 6'h1f == _T_94[5:0] ? welem[31] : _GEN_160; // @[Execute.scala 117:10]
  assign _GEN_162 = 6'h20 == _T_94[5:0] ? welem[32] : _GEN_161; // @[Execute.scala 117:10]
  assign _GEN_163 = 6'h21 == _T_94[5:0] ? welem[33] : _GEN_162; // @[Execute.scala 117:10]
  assign _GEN_164 = 6'h22 == _T_94[5:0] ? welem[34] : _GEN_163; // @[Execute.scala 117:10]
  assign _GEN_165 = 6'h23 == _T_94[5:0] ? welem[35] : _GEN_164; // @[Execute.scala 117:10]
  assign _GEN_166 = 6'h24 == _T_94[5:0] ? welem[36] : _GEN_165; // @[Execute.scala 117:10]
  assign _GEN_167 = 6'h25 == _T_94[5:0] ? welem[37] : _GEN_166; // @[Execute.scala 117:10]
  assign _GEN_168 = 6'h26 == _T_94[5:0] ? welem[38] : _GEN_167; // @[Execute.scala 117:10]
  assign _GEN_169 = 6'h27 == _T_94[5:0] ? welem[39] : _GEN_168; // @[Execute.scala 117:10]
  assign _GEN_170 = 6'h28 == _T_94[5:0] ? welem[40] : _GEN_169; // @[Execute.scala 117:10]
  assign _GEN_171 = 6'h29 == _T_94[5:0] ? welem[41] : _GEN_170; // @[Execute.scala 117:10]
  assign _GEN_172 = 6'h2a == _T_94[5:0] ? welem[42] : _GEN_171; // @[Execute.scala 117:10]
  assign _GEN_173 = 6'h2b == _T_94[5:0] ? welem[43] : _GEN_172; // @[Execute.scala 117:10]
  assign _GEN_174 = 6'h2c == _T_94[5:0] ? welem[44] : _GEN_173; // @[Execute.scala 117:10]
  assign _GEN_175 = 6'h2d == _T_94[5:0] ? welem[45] : _GEN_174; // @[Execute.scala 117:10]
  assign _GEN_176 = 6'h2e == _T_94[5:0] ? welem[46] : _GEN_175; // @[Execute.scala 117:10]
  assign _GEN_177 = 6'h2f == _T_94[5:0] ? welem[47] : _GEN_176; // @[Execute.scala 117:10]
  assign _GEN_178 = 6'h30 == _T_94[5:0] ? welem[48] : _GEN_177; // @[Execute.scala 117:10]
  assign _GEN_179 = 6'h31 == _T_94[5:0] ? welem[49] : _GEN_178; // @[Execute.scala 117:10]
  assign _GEN_180 = 6'h32 == _T_94[5:0] ? welem[50] : _GEN_179; // @[Execute.scala 117:10]
  assign _GEN_181 = 6'h33 == _T_94[5:0] ? welem[51] : _GEN_180; // @[Execute.scala 117:10]
  assign _GEN_182 = 6'h34 == _T_94[5:0] ? welem[52] : _GEN_181; // @[Execute.scala 117:10]
  assign _GEN_183 = 6'h35 == _T_94[5:0] ? welem[53] : _GEN_182; // @[Execute.scala 117:10]
  assign _GEN_184 = 6'h36 == _T_94[5:0] ? welem[54] : _GEN_183; // @[Execute.scala 117:10]
  assign _GEN_185 = 6'h37 == _T_94[5:0] ? welem[55] : _GEN_184; // @[Execute.scala 117:10]
  assign _GEN_186 = 6'h38 == _T_94[5:0] ? welem[56] : _GEN_185; // @[Execute.scala 117:10]
  assign _GEN_187 = 6'h39 == _T_94[5:0] ? welem[57] : _GEN_186; // @[Execute.scala 117:10]
  assign _GEN_188 = 6'h3a == _T_94[5:0] ? welem[58] : _GEN_187; // @[Execute.scala 117:10]
  assign _GEN_189 = 6'h3b == _T_94[5:0] ? welem[59] : _GEN_188; // @[Execute.scala 117:10]
  assign _GEN_190 = 6'h3c == _T_94[5:0] ? welem[60] : _GEN_189; // @[Execute.scala 117:10]
  assign _GEN_191 = 6'h3d == _T_94[5:0] ? welem[61] : _GEN_190; // @[Execute.scala 117:10]
  assign _GEN_192 = 6'h3e == _T_94[5:0] ? welem[62] : _GEN_191; // @[Execute.scala 117:10]
  assign _GEN_193 = 6'h3f == _T_94[5:0] ? welem[63] : _GEN_192; // @[Execute.scala 117:10]
  assign _T_102 = r < 6'h3f; // @[Execute.scala 117:15]
  assign _T_104 = r - 6'h3f; // @[Execute.scala 117:37]
  assign _T_108 = 6'h1 + r; // @[Execute.scala 117:60]
  assign _GEN_259 = 6'h1 == _T_104 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_260 = 6'h2 == _T_104 ? welem[2] : _GEN_259; // @[Execute.scala 117:10]
  assign _GEN_261 = 6'h3 == _T_104 ? welem[3] : _GEN_260; // @[Execute.scala 117:10]
  assign _GEN_262 = 6'h4 == _T_104 ? welem[4] : _GEN_261; // @[Execute.scala 117:10]
  assign _GEN_263 = 6'h5 == _T_104 ? welem[5] : _GEN_262; // @[Execute.scala 117:10]
  assign _GEN_264 = 6'h6 == _T_104 ? welem[6] : _GEN_263; // @[Execute.scala 117:10]
  assign _GEN_265 = 6'h7 == _T_104 ? welem[7] : _GEN_264; // @[Execute.scala 117:10]
  assign _GEN_266 = 6'h8 == _T_104 ? welem[8] : _GEN_265; // @[Execute.scala 117:10]
  assign _GEN_267 = 6'h9 == _T_104 ? welem[9] : _GEN_266; // @[Execute.scala 117:10]
  assign _GEN_268 = 6'ha == _T_104 ? welem[10] : _GEN_267; // @[Execute.scala 117:10]
  assign _GEN_269 = 6'hb == _T_104 ? welem[11] : _GEN_268; // @[Execute.scala 117:10]
  assign _GEN_270 = 6'hc == _T_104 ? welem[12] : _GEN_269; // @[Execute.scala 117:10]
  assign _GEN_271 = 6'hd == _T_104 ? welem[13] : _GEN_270; // @[Execute.scala 117:10]
  assign _GEN_272 = 6'he == _T_104 ? welem[14] : _GEN_271; // @[Execute.scala 117:10]
  assign _GEN_273 = 6'hf == _T_104 ? welem[15] : _GEN_272; // @[Execute.scala 117:10]
  assign _GEN_274 = 6'h10 == _T_104 ? welem[16] : _GEN_273; // @[Execute.scala 117:10]
  assign _GEN_275 = 6'h11 == _T_104 ? welem[17] : _GEN_274; // @[Execute.scala 117:10]
  assign _GEN_276 = 6'h12 == _T_104 ? welem[18] : _GEN_275; // @[Execute.scala 117:10]
  assign _GEN_277 = 6'h13 == _T_104 ? welem[19] : _GEN_276; // @[Execute.scala 117:10]
  assign _GEN_278 = 6'h14 == _T_104 ? welem[20] : _GEN_277; // @[Execute.scala 117:10]
  assign _GEN_279 = 6'h15 == _T_104 ? welem[21] : _GEN_278; // @[Execute.scala 117:10]
  assign _GEN_280 = 6'h16 == _T_104 ? welem[22] : _GEN_279; // @[Execute.scala 117:10]
  assign _GEN_281 = 6'h17 == _T_104 ? welem[23] : _GEN_280; // @[Execute.scala 117:10]
  assign _GEN_282 = 6'h18 == _T_104 ? welem[24] : _GEN_281; // @[Execute.scala 117:10]
  assign _GEN_283 = 6'h19 == _T_104 ? welem[25] : _GEN_282; // @[Execute.scala 117:10]
  assign _GEN_284 = 6'h1a == _T_104 ? welem[26] : _GEN_283; // @[Execute.scala 117:10]
  assign _GEN_285 = 6'h1b == _T_104 ? welem[27] : _GEN_284; // @[Execute.scala 117:10]
  assign _GEN_286 = 6'h1c == _T_104 ? welem[28] : _GEN_285; // @[Execute.scala 117:10]
  assign _GEN_287 = 6'h1d == _T_104 ? welem[29] : _GEN_286; // @[Execute.scala 117:10]
  assign _GEN_288 = 6'h1e == _T_104 ? welem[30] : _GEN_287; // @[Execute.scala 117:10]
  assign _GEN_289 = 6'h1f == _T_104 ? welem[31] : _GEN_288; // @[Execute.scala 117:10]
  assign _GEN_290 = 6'h20 == _T_104 ? welem[32] : _GEN_289; // @[Execute.scala 117:10]
  assign _GEN_291 = 6'h21 == _T_104 ? welem[33] : _GEN_290; // @[Execute.scala 117:10]
  assign _GEN_292 = 6'h22 == _T_104 ? welem[34] : _GEN_291; // @[Execute.scala 117:10]
  assign _GEN_293 = 6'h23 == _T_104 ? welem[35] : _GEN_292; // @[Execute.scala 117:10]
  assign _GEN_294 = 6'h24 == _T_104 ? welem[36] : _GEN_293; // @[Execute.scala 117:10]
  assign _GEN_295 = 6'h25 == _T_104 ? welem[37] : _GEN_294; // @[Execute.scala 117:10]
  assign _GEN_296 = 6'h26 == _T_104 ? welem[38] : _GEN_295; // @[Execute.scala 117:10]
  assign _GEN_297 = 6'h27 == _T_104 ? welem[39] : _GEN_296; // @[Execute.scala 117:10]
  assign _GEN_298 = 6'h28 == _T_104 ? welem[40] : _GEN_297; // @[Execute.scala 117:10]
  assign _GEN_299 = 6'h29 == _T_104 ? welem[41] : _GEN_298; // @[Execute.scala 117:10]
  assign _GEN_300 = 6'h2a == _T_104 ? welem[42] : _GEN_299; // @[Execute.scala 117:10]
  assign _GEN_301 = 6'h2b == _T_104 ? welem[43] : _GEN_300; // @[Execute.scala 117:10]
  assign _GEN_302 = 6'h2c == _T_104 ? welem[44] : _GEN_301; // @[Execute.scala 117:10]
  assign _GEN_303 = 6'h2d == _T_104 ? welem[45] : _GEN_302; // @[Execute.scala 117:10]
  assign _GEN_304 = 6'h2e == _T_104 ? welem[46] : _GEN_303; // @[Execute.scala 117:10]
  assign _GEN_305 = 6'h2f == _T_104 ? welem[47] : _GEN_304; // @[Execute.scala 117:10]
  assign _GEN_306 = 6'h30 == _T_104 ? welem[48] : _GEN_305; // @[Execute.scala 117:10]
  assign _GEN_307 = 6'h31 == _T_104 ? welem[49] : _GEN_306; // @[Execute.scala 117:10]
  assign _GEN_308 = 6'h32 == _T_104 ? welem[50] : _GEN_307; // @[Execute.scala 117:10]
  assign _GEN_309 = 6'h33 == _T_104 ? welem[51] : _GEN_308; // @[Execute.scala 117:10]
  assign _GEN_310 = 6'h34 == _T_104 ? welem[52] : _GEN_309; // @[Execute.scala 117:10]
  assign _GEN_311 = 6'h35 == _T_104 ? welem[53] : _GEN_310; // @[Execute.scala 117:10]
  assign _GEN_312 = 6'h36 == _T_104 ? welem[54] : _GEN_311; // @[Execute.scala 117:10]
  assign _GEN_313 = 6'h37 == _T_104 ? welem[55] : _GEN_312; // @[Execute.scala 117:10]
  assign _GEN_314 = 6'h38 == _T_104 ? welem[56] : _GEN_313; // @[Execute.scala 117:10]
  assign _GEN_315 = 6'h39 == _T_104 ? welem[57] : _GEN_314; // @[Execute.scala 117:10]
  assign _GEN_316 = 6'h3a == _T_104 ? welem[58] : _GEN_315; // @[Execute.scala 117:10]
  assign _GEN_317 = 6'h3b == _T_104 ? welem[59] : _GEN_316; // @[Execute.scala 117:10]
  assign _GEN_318 = 6'h3c == _T_104 ? welem[60] : _GEN_317; // @[Execute.scala 117:10]
  assign _GEN_319 = 6'h3d == _T_104 ? welem[61] : _GEN_318; // @[Execute.scala 117:10]
  assign _GEN_320 = 6'h3e == _T_104 ? welem[62] : _GEN_319; // @[Execute.scala 117:10]
  assign _GEN_321 = 6'h3f == _T_104 ? welem[63] : _GEN_320; // @[Execute.scala 117:10]
  assign _GEN_323 = 6'h1 == _T_108 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_324 = 6'h2 == _T_108 ? welem[2] : _GEN_323; // @[Execute.scala 117:10]
  assign _GEN_325 = 6'h3 == _T_108 ? welem[3] : _GEN_324; // @[Execute.scala 117:10]
  assign _GEN_326 = 6'h4 == _T_108 ? welem[4] : _GEN_325; // @[Execute.scala 117:10]
  assign _GEN_327 = 6'h5 == _T_108 ? welem[5] : _GEN_326; // @[Execute.scala 117:10]
  assign _GEN_328 = 6'h6 == _T_108 ? welem[6] : _GEN_327; // @[Execute.scala 117:10]
  assign _GEN_329 = 6'h7 == _T_108 ? welem[7] : _GEN_328; // @[Execute.scala 117:10]
  assign _GEN_330 = 6'h8 == _T_108 ? welem[8] : _GEN_329; // @[Execute.scala 117:10]
  assign _GEN_331 = 6'h9 == _T_108 ? welem[9] : _GEN_330; // @[Execute.scala 117:10]
  assign _GEN_332 = 6'ha == _T_108 ? welem[10] : _GEN_331; // @[Execute.scala 117:10]
  assign _GEN_333 = 6'hb == _T_108 ? welem[11] : _GEN_332; // @[Execute.scala 117:10]
  assign _GEN_334 = 6'hc == _T_108 ? welem[12] : _GEN_333; // @[Execute.scala 117:10]
  assign _GEN_335 = 6'hd == _T_108 ? welem[13] : _GEN_334; // @[Execute.scala 117:10]
  assign _GEN_336 = 6'he == _T_108 ? welem[14] : _GEN_335; // @[Execute.scala 117:10]
  assign _GEN_337 = 6'hf == _T_108 ? welem[15] : _GEN_336; // @[Execute.scala 117:10]
  assign _GEN_338 = 6'h10 == _T_108 ? welem[16] : _GEN_337; // @[Execute.scala 117:10]
  assign _GEN_339 = 6'h11 == _T_108 ? welem[17] : _GEN_338; // @[Execute.scala 117:10]
  assign _GEN_340 = 6'h12 == _T_108 ? welem[18] : _GEN_339; // @[Execute.scala 117:10]
  assign _GEN_341 = 6'h13 == _T_108 ? welem[19] : _GEN_340; // @[Execute.scala 117:10]
  assign _GEN_342 = 6'h14 == _T_108 ? welem[20] : _GEN_341; // @[Execute.scala 117:10]
  assign _GEN_343 = 6'h15 == _T_108 ? welem[21] : _GEN_342; // @[Execute.scala 117:10]
  assign _GEN_344 = 6'h16 == _T_108 ? welem[22] : _GEN_343; // @[Execute.scala 117:10]
  assign _GEN_345 = 6'h17 == _T_108 ? welem[23] : _GEN_344; // @[Execute.scala 117:10]
  assign _GEN_346 = 6'h18 == _T_108 ? welem[24] : _GEN_345; // @[Execute.scala 117:10]
  assign _GEN_347 = 6'h19 == _T_108 ? welem[25] : _GEN_346; // @[Execute.scala 117:10]
  assign _GEN_348 = 6'h1a == _T_108 ? welem[26] : _GEN_347; // @[Execute.scala 117:10]
  assign _GEN_349 = 6'h1b == _T_108 ? welem[27] : _GEN_348; // @[Execute.scala 117:10]
  assign _GEN_350 = 6'h1c == _T_108 ? welem[28] : _GEN_349; // @[Execute.scala 117:10]
  assign _GEN_351 = 6'h1d == _T_108 ? welem[29] : _GEN_350; // @[Execute.scala 117:10]
  assign _GEN_352 = 6'h1e == _T_108 ? welem[30] : _GEN_351; // @[Execute.scala 117:10]
  assign _GEN_353 = 6'h1f == _T_108 ? welem[31] : _GEN_352; // @[Execute.scala 117:10]
  assign _GEN_354 = 6'h20 == _T_108 ? welem[32] : _GEN_353; // @[Execute.scala 117:10]
  assign _GEN_355 = 6'h21 == _T_108 ? welem[33] : _GEN_354; // @[Execute.scala 117:10]
  assign _GEN_356 = 6'h22 == _T_108 ? welem[34] : _GEN_355; // @[Execute.scala 117:10]
  assign _GEN_357 = 6'h23 == _T_108 ? welem[35] : _GEN_356; // @[Execute.scala 117:10]
  assign _GEN_358 = 6'h24 == _T_108 ? welem[36] : _GEN_357; // @[Execute.scala 117:10]
  assign _GEN_359 = 6'h25 == _T_108 ? welem[37] : _GEN_358; // @[Execute.scala 117:10]
  assign _GEN_360 = 6'h26 == _T_108 ? welem[38] : _GEN_359; // @[Execute.scala 117:10]
  assign _GEN_361 = 6'h27 == _T_108 ? welem[39] : _GEN_360; // @[Execute.scala 117:10]
  assign _GEN_362 = 6'h28 == _T_108 ? welem[40] : _GEN_361; // @[Execute.scala 117:10]
  assign _GEN_363 = 6'h29 == _T_108 ? welem[41] : _GEN_362; // @[Execute.scala 117:10]
  assign _GEN_364 = 6'h2a == _T_108 ? welem[42] : _GEN_363; // @[Execute.scala 117:10]
  assign _GEN_365 = 6'h2b == _T_108 ? welem[43] : _GEN_364; // @[Execute.scala 117:10]
  assign _GEN_366 = 6'h2c == _T_108 ? welem[44] : _GEN_365; // @[Execute.scala 117:10]
  assign _GEN_367 = 6'h2d == _T_108 ? welem[45] : _GEN_366; // @[Execute.scala 117:10]
  assign _GEN_368 = 6'h2e == _T_108 ? welem[46] : _GEN_367; // @[Execute.scala 117:10]
  assign _GEN_369 = 6'h2f == _T_108 ? welem[47] : _GEN_368; // @[Execute.scala 117:10]
  assign _GEN_370 = 6'h30 == _T_108 ? welem[48] : _GEN_369; // @[Execute.scala 117:10]
  assign _GEN_371 = 6'h31 == _T_108 ? welem[49] : _GEN_370; // @[Execute.scala 117:10]
  assign _GEN_372 = 6'h32 == _T_108 ? welem[50] : _GEN_371; // @[Execute.scala 117:10]
  assign _GEN_373 = 6'h33 == _T_108 ? welem[51] : _GEN_372; // @[Execute.scala 117:10]
  assign _GEN_374 = 6'h34 == _T_108 ? welem[52] : _GEN_373; // @[Execute.scala 117:10]
  assign _GEN_375 = 6'h35 == _T_108 ? welem[53] : _GEN_374; // @[Execute.scala 117:10]
  assign _GEN_376 = 6'h36 == _T_108 ? welem[54] : _GEN_375; // @[Execute.scala 117:10]
  assign _GEN_377 = 6'h37 == _T_108 ? welem[55] : _GEN_376; // @[Execute.scala 117:10]
  assign _GEN_378 = 6'h38 == _T_108 ? welem[56] : _GEN_377; // @[Execute.scala 117:10]
  assign _GEN_379 = 6'h39 == _T_108 ? welem[57] : _GEN_378; // @[Execute.scala 117:10]
  assign _GEN_380 = 6'h3a == _T_108 ? welem[58] : _GEN_379; // @[Execute.scala 117:10]
  assign _GEN_381 = 6'h3b == _T_108 ? welem[59] : _GEN_380; // @[Execute.scala 117:10]
  assign _GEN_382 = 6'h3c == _T_108 ? welem[60] : _GEN_381; // @[Execute.scala 117:10]
  assign _GEN_383 = 6'h3d == _T_108 ? welem[61] : _GEN_382; // @[Execute.scala 117:10]
  assign _GEN_384 = 6'h3e == _T_108 ? welem[62] : _GEN_383; // @[Execute.scala 117:10]
  assign _GEN_385 = 6'h3f == _T_108 ? welem[63] : _GEN_384; // @[Execute.scala 117:10]
  assign _T_111 = _T_102 ? _GEN_321 : _GEN_385; // @[Execute.scala 117:10]
  assign _T_112 = r < 6'h3e; // @[Execute.scala 117:15]
  assign _T_114 = r - 6'h3e; // @[Execute.scala 117:37]
  assign _T_118 = 6'h2 + r; // @[Execute.scala 117:60]
  assign _GEN_387 = 6'h1 == _T_114 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_388 = 6'h2 == _T_114 ? welem[2] : _GEN_387; // @[Execute.scala 117:10]
  assign _GEN_389 = 6'h3 == _T_114 ? welem[3] : _GEN_388; // @[Execute.scala 117:10]
  assign _GEN_390 = 6'h4 == _T_114 ? welem[4] : _GEN_389; // @[Execute.scala 117:10]
  assign _GEN_391 = 6'h5 == _T_114 ? welem[5] : _GEN_390; // @[Execute.scala 117:10]
  assign _GEN_392 = 6'h6 == _T_114 ? welem[6] : _GEN_391; // @[Execute.scala 117:10]
  assign _GEN_393 = 6'h7 == _T_114 ? welem[7] : _GEN_392; // @[Execute.scala 117:10]
  assign _GEN_394 = 6'h8 == _T_114 ? welem[8] : _GEN_393; // @[Execute.scala 117:10]
  assign _GEN_395 = 6'h9 == _T_114 ? welem[9] : _GEN_394; // @[Execute.scala 117:10]
  assign _GEN_396 = 6'ha == _T_114 ? welem[10] : _GEN_395; // @[Execute.scala 117:10]
  assign _GEN_397 = 6'hb == _T_114 ? welem[11] : _GEN_396; // @[Execute.scala 117:10]
  assign _GEN_398 = 6'hc == _T_114 ? welem[12] : _GEN_397; // @[Execute.scala 117:10]
  assign _GEN_399 = 6'hd == _T_114 ? welem[13] : _GEN_398; // @[Execute.scala 117:10]
  assign _GEN_400 = 6'he == _T_114 ? welem[14] : _GEN_399; // @[Execute.scala 117:10]
  assign _GEN_401 = 6'hf == _T_114 ? welem[15] : _GEN_400; // @[Execute.scala 117:10]
  assign _GEN_402 = 6'h10 == _T_114 ? welem[16] : _GEN_401; // @[Execute.scala 117:10]
  assign _GEN_403 = 6'h11 == _T_114 ? welem[17] : _GEN_402; // @[Execute.scala 117:10]
  assign _GEN_404 = 6'h12 == _T_114 ? welem[18] : _GEN_403; // @[Execute.scala 117:10]
  assign _GEN_405 = 6'h13 == _T_114 ? welem[19] : _GEN_404; // @[Execute.scala 117:10]
  assign _GEN_406 = 6'h14 == _T_114 ? welem[20] : _GEN_405; // @[Execute.scala 117:10]
  assign _GEN_407 = 6'h15 == _T_114 ? welem[21] : _GEN_406; // @[Execute.scala 117:10]
  assign _GEN_408 = 6'h16 == _T_114 ? welem[22] : _GEN_407; // @[Execute.scala 117:10]
  assign _GEN_409 = 6'h17 == _T_114 ? welem[23] : _GEN_408; // @[Execute.scala 117:10]
  assign _GEN_410 = 6'h18 == _T_114 ? welem[24] : _GEN_409; // @[Execute.scala 117:10]
  assign _GEN_411 = 6'h19 == _T_114 ? welem[25] : _GEN_410; // @[Execute.scala 117:10]
  assign _GEN_412 = 6'h1a == _T_114 ? welem[26] : _GEN_411; // @[Execute.scala 117:10]
  assign _GEN_413 = 6'h1b == _T_114 ? welem[27] : _GEN_412; // @[Execute.scala 117:10]
  assign _GEN_414 = 6'h1c == _T_114 ? welem[28] : _GEN_413; // @[Execute.scala 117:10]
  assign _GEN_415 = 6'h1d == _T_114 ? welem[29] : _GEN_414; // @[Execute.scala 117:10]
  assign _GEN_416 = 6'h1e == _T_114 ? welem[30] : _GEN_415; // @[Execute.scala 117:10]
  assign _GEN_417 = 6'h1f == _T_114 ? welem[31] : _GEN_416; // @[Execute.scala 117:10]
  assign _GEN_418 = 6'h20 == _T_114 ? welem[32] : _GEN_417; // @[Execute.scala 117:10]
  assign _GEN_419 = 6'h21 == _T_114 ? welem[33] : _GEN_418; // @[Execute.scala 117:10]
  assign _GEN_420 = 6'h22 == _T_114 ? welem[34] : _GEN_419; // @[Execute.scala 117:10]
  assign _GEN_421 = 6'h23 == _T_114 ? welem[35] : _GEN_420; // @[Execute.scala 117:10]
  assign _GEN_422 = 6'h24 == _T_114 ? welem[36] : _GEN_421; // @[Execute.scala 117:10]
  assign _GEN_423 = 6'h25 == _T_114 ? welem[37] : _GEN_422; // @[Execute.scala 117:10]
  assign _GEN_424 = 6'h26 == _T_114 ? welem[38] : _GEN_423; // @[Execute.scala 117:10]
  assign _GEN_425 = 6'h27 == _T_114 ? welem[39] : _GEN_424; // @[Execute.scala 117:10]
  assign _GEN_426 = 6'h28 == _T_114 ? welem[40] : _GEN_425; // @[Execute.scala 117:10]
  assign _GEN_427 = 6'h29 == _T_114 ? welem[41] : _GEN_426; // @[Execute.scala 117:10]
  assign _GEN_428 = 6'h2a == _T_114 ? welem[42] : _GEN_427; // @[Execute.scala 117:10]
  assign _GEN_429 = 6'h2b == _T_114 ? welem[43] : _GEN_428; // @[Execute.scala 117:10]
  assign _GEN_430 = 6'h2c == _T_114 ? welem[44] : _GEN_429; // @[Execute.scala 117:10]
  assign _GEN_431 = 6'h2d == _T_114 ? welem[45] : _GEN_430; // @[Execute.scala 117:10]
  assign _GEN_432 = 6'h2e == _T_114 ? welem[46] : _GEN_431; // @[Execute.scala 117:10]
  assign _GEN_433 = 6'h2f == _T_114 ? welem[47] : _GEN_432; // @[Execute.scala 117:10]
  assign _GEN_434 = 6'h30 == _T_114 ? welem[48] : _GEN_433; // @[Execute.scala 117:10]
  assign _GEN_435 = 6'h31 == _T_114 ? welem[49] : _GEN_434; // @[Execute.scala 117:10]
  assign _GEN_436 = 6'h32 == _T_114 ? welem[50] : _GEN_435; // @[Execute.scala 117:10]
  assign _GEN_437 = 6'h33 == _T_114 ? welem[51] : _GEN_436; // @[Execute.scala 117:10]
  assign _GEN_438 = 6'h34 == _T_114 ? welem[52] : _GEN_437; // @[Execute.scala 117:10]
  assign _GEN_439 = 6'h35 == _T_114 ? welem[53] : _GEN_438; // @[Execute.scala 117:10]
  assign _GEN_440 = 6'h36 == _T_114 ? welem[54] : _GEN_439; // @[Execute.scala 117:10]
  assign _GEN_441 = 6'h37 == _T_114 ? welem[55] : _GEN_440; // @[Execute.scala 117:10]
  assign _GEN_442 = 6'h38 == _T_114 ? welem[56] : _GEN_441; // @[Execute.scala 117:10]
  assign _GEN_443 = 6'h39 == _T_114 ? welem[57] : _GEN_442; // @[Execute.scala 117:10]
  assign _GEN_444 = 6'h3a == _T_114 ? welem[58] : _GEN_443; // @[Execute.scala 117:10]
  assign _GEN_445 = 6'h3b == _T_114 ? welem[59] : _GEN_444; // @[Execute.scala 117:10]
  assign _GEN_446 = 6'h3c == _T_114 ? welem[60] : _GEN_445; // @[Execute.scala 117:10]
  assign _GEN_447 = 6'h3d == _T_114 ? welem[61] : _GEN_446; // @[Execute.scala 117:10]
  assign _GEN_448 = 6'h3e == _T_114 ? welem[62] : _GEN_447; // @[Execute.scala 117:10]
  assign _GEN_449 = 6'h3f == _T_114 ? welem[63] : _GEN_448; // @[Execute.scala 117:10]
  assign _GEN_451 = 6'h1 == _T_118 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_452 = 6'h2 == _T_118 ? welem[2] : _GEN_451; // @[Execute.scala 117:10]
  assign _GEN_453 = 6'h3 == _T_118 ? welem[3] : _GEN_452; // @[Execute.scala 117:10]
  assign _GEN_454 = 6'h4 == _T_118 ? welem[4] : _GEN_453; // @[Execute.scala 117:10]
  assign _GEN_455 = 6'h5 == _T_118 ? welem[5] : _GEN_454; // @[Execute.scala 117:10]
  assign _GEN_456 = 6'h6 == _T_118 ? welem[6] : _GEN_455; // @[Execute.scala 117:10]
  assign _GEN_457 = 6'h7 == _T_118 ? welem[7] : _GEN_456; // @[Execute.scala 117:10]
  assign _GEN_458 = 6'h8 == _T_118 ? welem[8] : _GEN_457; // @[Execute.scala 117:10]
  assign _GEN_459 = 6'h9 == _T_118 ? welem[9] : _GEN_458; // @[Execute.scala 117:10]
  assign _GEN_460 = 6'ha == _T_118 ? welem[10] : _GEN_459; // @[Execute.scala 117:10]
  assign _GEN_461 = 6'hb == _T_118 ? welem[11] : _GEN_460; // @[Execute.scala 117:10]
  assign _GEN_462 = 6'hc == _T_118 ? welem[12] : _GEN_461; // @[Execute.scala 117:10]
  assign _GEN_463 = 6'hd == _T_118 ? welem[13] : _GEN_462; // @[Execute.scala 117:10]
  assign _GEN_464 = 6'he == _T_118 ? welem[14] : _GEN_463; // @[Execute.scala 117:10]
  assign _GEN_465 = 6'hf == _T_118 ? welem[15] : _GEN_464; // @[Execute.scala 117:10]
  assign _GEN_466 = 6'h10 == _T_118 ? welem[16] : _GEN_465; // @[Execute.scala 117:10]
  assign _GEN_467 = 6'h11 == _T_118 ? welem[17] : _GEN_466; // @[Execute.scala 117:10]
  assign _GEN_468 = 6'h12 == _T_118 ? welem[18] : _GEN_467; // @[Execute.scala 117:10]
  assign _GEN_469 = 6'h13 == _T_118 ? welem[19] : _GEN_468; // @[Execute.scala 117:10]
  assign _GEN_470 = 6'h14 == _T_118 ? welem[20] : _GEN_469; // @[Execute.scala 117:10]
  assign _GEN_471 = 6'h15 == _T_118 ? welem[21] : _GEN_470; // @[Execute.scala 117:10]
  assign _GEN_472 = 6'h16 == _T_118 ? welem[22] : _GEN_471; // @[Execute.scala 117:10]
  assign _GEN_473 = 6'h17 == _T_118 ? welem[23] : _GEN_472; // @[Execute.scala 117:10]
  assign _GEN_474 = 6'h18 == _T_118 ? welem[24] : _GEN_473; // @[Execute.scala 117:10]
  assign _GEN_475 = 6'h19 == _T_118 ? welem[25] : _GEN_474; // @[Execute.scala 117:10]
  assign _GEN_476 = 6'h1a == _T_118 ? welem[26] : _GEN_475; // @[Execute.scala 117:10]
  assign _GEN_477 = 6'h1b == _T_118 ? welem[27] : _GEN_476; // @[Execute.scala 117:10]
  assign _GEN_478 = 6'h1c == _T_118 ? welem[28] : _GEN_477; // @[Execute.scala 117:10]
  assign _GEN_479 = 6'h1d == _T_118 ? welem[29] : _GEN_478; // @[Execute.scala 117:10]
  assign _GEN_480 = 6'h1e == _T_118 ? welem[30] : _GEN_479; // @[Execute.scala 117:10]
  assign _GEN_481 = 6'h1f == _T_118 ? welem[31] : _GEN_480; // @[Execute.scala 117:10]
  assign _GEN_482 = 6'h20 == _T_118 ? welem[32] : _GEN_481; // @[Execute.scala 117:10]
  assign _GEN_483 = 6'h21 == _T_118 ? welem[33] : _GEN_482; // @[Execute.scala 117:10]
  assign _GEN_484 = 6'h22 == _T_118 ? welem[34] : _GEN_483; // @[Execute.scala 117:10]
  assign _GEN_485 = 6'h23 == _T_118 ? welem[35] : _GEN_484; // @[Execute.scala 117:10]
  assign _GEN_486 = 6'h24 == _T_118 ? welem[36] : _GEN_485; // @[Execute.scala 117:10]
  assign _GEN_487 = 6'h25 == _T_118 ? welem[37] : _GEN_486; // @[Execute.scala 117:10]
  assign _GEN_488 = 6'h26 == _T_118 ? welem[38] : _GEN_487; // @[Execute.scala 117:10]
  assign _GEN_489 = 6'h27 == _T_118 ? welem[39] : _GEN_488; // @[Execute.scala 117:10]
  assign _GEN_490 = 6'h28 == _T_118 ? welem[40] : _GEN_489; // @[Execute.scala 117:10]
  assign _GEN_491 = 6'h29 == _T_118 ? welem[41] : _GEN_490; // @[Execute.scala 117:10]
  assign _GEN_492 = 6'h2a == _T_118 ? welem[42] : _GEN_491; // @[Execute.scala 117:10]
  assign _GEN_493 = 6'h2b == _T_118 ? welem[43] : _GEN_492; // @[Execute.scala 117:10]
  assign _GEN_494 = 6'h2c == _T_118 ? welem[44] : _GEN_493; // @[Execute.scala 117:10]
  assign _GEN_495 = 6'h2d == _T_118 ? welem[45] : _GEN_494; // @[Execute.scala 117:10]
  assign _GEN_496 = 6'h2e == _T_118 ? welem[46] : _GEN_495; // @[Execute.scala 117:10]
  assign _GEN_497 = 6'h2f == _T_118 ? welem[47] : _GEN_496; // @[Execute.scala 117:10]
  assign _GEN_498 = 6'h30 == _T_118 ? welem[48] : _GEN_497; // @[Execute.scala 117:10]
  assign _GEN_499 = 6'h31 == _T_118 ? welem[49] : _GEN_498; // @[Execute.scala 117:10]
  assign _GEN_500 = 6'h32 == _T_118 ? welem[50] : _GEN_499; // @[Execute.scala 117:10]
  assign _GEN_501 = 6'h33 == _T_118 ? welem[51] : _GEN_500; // @[Execute.scala 117:10]
  assign _GEN_502 = 6'h34 == _T_118 ? welem[52] : _GEN_501; // @[Execute.scala 117:10]
  assign _GEN_503 = 6'h35 == _T_118 ? welem[53] : _GEN_502; // @[Execute.scala 117:10]
  assign _GEN_504 = 6'h36 == _T_118 ? welem[54] : _GEN_503; // @[Execute.scala 117:10]
  assign _GEN_505 = 6'h37 == _T_118 ? welem[55] : _GEN_504; // @[Execute.scala 117:10]
  assign _GEN_506 = 6'h38 == _T_118 ? welem[56] : _GEN_505; // @[Execute.scala 117:10]
  assign _GEN_507 = 6'h39 == _T_118 ? welem[57] : _GEN_506; // @[Execute.scala 117:10]
  assign _GEN_508 = 6'h3a == _T_118 ? welem[58] : _GEN_507; // @[Execute.scala 117:10]
  assign _GEN_509 = 6'h3b == _T_118 ? welem[59] : _GEN_508; // @[Execute.scala 117:10]
  assign _GEN_510 = 6'h3c == _T_118 ? welem[60] : _GEN_509; // @[Execute.scala 117:10]
  assign _GEN_511 = 6'h3d == _T_118 ? welem[61] : _GEN_510; // @[Execute.scala 117:10]
  assign _GEN_512 = 6'h3e == _T_118 ? welem[62] : _GEN_511; // @[Execute.scala 117:10]
  assign _GEN_513 = 6'h3f == _T_118 ? welem[63] : _GEN_512; // @[Execute.scala 117:10]
  assign _T_121 = _T_112 ? _GEN_449 : _GEN_513; // @[Execute.scala 117:10]
  assign _T_122 = r < 6'h3d; // @[Execute.scala 117:15]
  assign _T_124 = r - 6'h3d; // @[Execute.scala 117:37]
  assign _T_128 = 6'h3 + r; // @[Execute.scala 117:60]
  assign _GEN_515 = 6'h1 == _T_124 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_516 = 6'h2 == _T_124 ? welem[2] : _GEN_515; // @[Execute.scala 117:10]
  assign _GEN_517 = 6'h3 == _T_124 ? welem[3] : _GEN_516; // @[Execute.scala 117:10]
  assign _GEN_518 = 6'h4 == _T_124 ? welem[4] : _GEN_517; // @[Execute.scala 117:10]
  assign _GEN_519 = 6'h5 == _T_124 ? welem[5] : _GEN_518; // @[Execute.scala 117:10]
  assign _GEN_520 = 6'h6 == _T_124 ? welem[6] : _GEN_519; // @[Execute.scala 117:10]
  assign _GEN_521 = 6'h7 == _T_124 ? welem[7] : _GEN_520; // @[Execute.scala 117:10]
  assign _GEN_522 = 6'h8 == _T_124 ? welem[8] : _GEN_521; // @[Execute.scala 117:10]
  assign _GEN_523 = 6'h9 == _T_124 ? welem[9] : _GEN_522; // @[Execute.scala 117:10]
  assign _GEN_524 = 6'ha == _T_124 ? welem[10] : _GEN_523; // @[Execute.scala 117:10]
  assign _GEN_525 = 6'hb == _T_124 ? welem[11] : _GEN_524; // @[Execute.scala 117:10]
  assign _GEN_526 = 6'hc == _T_124 ? welem[12] : _GEN_525; // @[Execute.scala 117:10]
  assign _GEN_527 = 6'hd == _T_124 ? welem[13] : _GEN_526; // @[Execute.scala 117:10]
  assign _GEN_528 = 6'he == _T_124 ? welem[14] : _GEN_527; // @[Execute.scala 117:10]
  assign _GEN_529 = 6'hf == _T_124 ? welem[15] : _GEN_528; // @[Execute.scala 117:10]
  assign _GEN_530 = 6'h10 == _T_124 ? welem[16] : _GEN_529; // @[Execute.scala 117:10]
  assign _GEN_531 = 6'h11 == _T_124 ? welem[17] : _GEN_530; // @[Execute.scala 117:10]
  assign _GEN_532 = 6'h12 == _T_124 ? welem[18] : _GEN_531; // @[Execute.scala 117:10]
  assign _GEN_533 = 6'h13 == _T_124 ? welem[19] : _GEN_532; // @[Execute.scala 117:10]
  assign _GEN_534 = 6'h14 == _T_124 ? welem[20] : _GEN_533; // @[Execute.scala 117:10]
  assign _GEN_535 = 6'h15 == _T_124 ? welem[21] : _GEN_534; // @[Execute.scala 117:10]
  assign _GEN_536 = 6'h16 == _T_124 ? welem[22] : _GEN_535; // @[Execute.scala 117:10]
  assign _GEN_537 = 6'h17 == _T_124 ? welem[23] : _GEN_536; // @[Execute.scala 117:10]
  assign _GEN_538 = 6'h18 == _T_124 ? welem[24] : _GEN_537; // @[Execute.scala 117:10]
  assign _GEN_539 = 6'h19 == _T_124 ? welem[25] : _GEN_538; // @[Execute.scala 117:10]
  assign _GEN_540 = 6'h1a == _T_124 ? welem[26] : _GEN_539; // @[Execute.scala 117:10]
  assign _GEN_541 = 6'h1b == _T_124 ? welem[27] : _GEN_540; // @[Execute.scala 117:10]
  assign _GEN_542 = 6'h1c == _T_124 ? welem[28] : _GEN_541; // @[Execute.scala 117:10]
  assign _GEN_543 = 6'h1d == _T_124 ? welem[29] : _GEN_542; // @[Execute.scala 117:10]
  assign _GEN_544 = 6'h1e == _T_124 ? welem[30] : _GEN_543; // @[Execute.scala 117:10]
  assign _GEN_545 = 6'h1f == _T_124 ? welem[31] : _GEN_544; // @[Execute.scala 117:10]
  assign _GEN_546 = 6'h20 == _T_124 ? welem[32] : _GEN_545; // @[Execute.scala 117:10]
  assign _GEN_547 = 6'h21 == _T_124 ? welem[33] : _GEN_546; // @[Execute.scala 117:10]
  assign _GEN_548 = 6'h22 == _T_124 ? welem[34] : _GEN_547; // @[Execute.scala 117:10]
  assign _GEN_549 = 6'h23 == _T_124 ? welem[35] : _GEN_548; // @[Execute.scala 117:10]
  assign _GEN_550 = 6'h24 == _T_124 ? welem[36] : _GEN_549; // @[Execute.scala 117:10]
  assign _GEN_551 = 6'h25 == _T_124 ? welem[37] : _GEN_550; // @[Execute.scala 117:10]
  assign _GEN_552 = 6'h26 == _T_124 ? welem[38] : _GEN_551; // @[Execute.scala 117:10]
  assign _GEN_553 = 6'h27 == _T_124 ? welem[39] : _GEN_552; // @[Execute.scala 117:10]
  assign _GEN_554 = 6'h28 == _T_124 ? welem[40] : _GEN_553; // @[Execute.scala 117:10]
  assign _GEN_555 = 6'h29 == _T_124 ? welem[41] : _GEN_554; // @[Execute.scala 117:10]
  assign _GEN_556 = 6'h2a == _T_124 ? welem[42] : _GEN_555; // @[Execute.scala 117:10]
  assign _GEN_557 = 6'h2b == _T_124 ? welem[43] : _GEN_556; // @[Execute.scala 117:10]
  assign _GEN_558 = 6'h2c == _T_124 ? welem[44] : _GEN_557; // @[Execute.scala 117:10]
  assign _GEN_559 = 6'h2d == _T_124 ? welem[45] : _GEN_558; // @[Execute.scala 117:10]
  assign _GEN_560 = 6'h2e == _T_124 ? welem[46] : _GEN_559; // @[Execute.scala 117:10]
  assign _GEN_561 = 6'h2f == _T_124 ? welem[47] : _GEN_560; // @[Execute.scala 117:10]
  assign _GEN_562 = 6'h30 == _T_124 ? welem[48] : _GEN_561; // @[Execute.scala 117:10]
  assign _GEN_563 = 6'h31 == _T_124 ? welem[49] : _GEN_562; // @[Execute.scala 117:10]
  assign _GEN_564 = 6'h32 == _T_124 ? welem[50] : _GEN_563; // @[Execute.scala 117:10]
  assign _GEN_565 = 6'h33 == _T_124 ? welem[51] : _GEN_564; // @[Execute.scala 117:10]
  assign _GEN_566 = 6'h34 == _T_124 ? welem[52] : _GEN_565; // @[Execute.scala 117:10]
  assign _GEN_567 = 6'h35 == _T_124 ? welem[53] : _GEN_566; // @[Execute.scala 117:10]
  assign _GEN_568 = 6'h36 == _T_124 ? welem[54] : _GEN_567; // @[Execute.scala 117:10]
  assign _GEN_569 = 6'h37 == _T_124 ? welem[55] : _GEN_568; // @[Execute.scala 117:10]
  assign _GEN_570 = 6'h38 == _T_124 ? welem[56] : _GEN_569; // @[Execute.scala 117:10]
  assign _GEN_571 = 6'h39 == _T_124 ? welem[57] : _GEN_570; // @[Execute.scala 117:10]
  assign _GEN_572 = 6'h3a == _T_124 ? welem[58] : _GEN_571; // @[Execute.scala 117:10]
  assign _GEN_573 = 6'h3b == _T_124 ? welem[59] : _GEN_572; // @[Execute.scala 117:10]
  assign _GEN_574 = 6'h3c == _T_124 ? welem[60] : _GEN_573; // @[Execute.scala 117:10]
  assign _GEN_575 = 6'h3d == _T_124 ? welem[61] : _GEN_574; // @[Execute.scala 117:10]
  assign _GEN_576 = 6'h3e == _T_124 ? welem[62] : _GEN_575; // @[Execute.scala 117:10]
  assign _GEN_577 = 6'h3f == _T_124 ? welem[63] : _GEN_576; // @[Execute.scala 117:10]
  assign _GEN_579 = 6'h1 == _T_128 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_580 = 6'h2 == _T_128 ? welem[2] : _GEN_579; // @[Execute.scala 117:10]
  assign _GEN_581 = 6'h3 == _T_128 ? welem[3] : _GEN_580; // @[Execute.scala 117:10]
  assign _GEN_582 = 6'h4 == _T_128 ? welem[4] : _GEN_581; // @[Execute.scala 117:10]
  assign _GEN_583 = 6'h5 == _T_128 ? welem[5] : _GEN_582; // @[Execute.scala 117:10]
  assign _GEN_584 = 6'h6 == _T_128 ? welem[6] : _GEN_583; // @[Execute.scala 117:10]
  assign _GEN_585 = 6'h7 == _T_128 ? welem[7] : _GEN_584; // @[Execute.scala 117:10]
  assign _GEN_586 = 6'h8 == _T_128 ? welem[8] : _GEN_585; // @[Execute.scala 117:10]
  assign _GEN_587 = 6'h9 == _T_128 ? welem[9] : _GEN_586; // @[Execute.scala 117:10]
  assign _GEN_588 = 6'ha == _T_128 ? welem[10] : _GEN_587; // @[Execute.scala 117:10]
  assign _GEN_589 = 6'hb == _T_128 ? welem[11] : _GEN_588; // @[Execute.scala 117:10]
  assign _GEN_590 = 6'hc == _T_128 ? welem[12] : _GEN_589; // @[Execute.scala 117:10]
  assign _GEN_591 = 6'hd == _T_128 ? welem[13] : _GEN_590; // @[Execute.scala 117:10]
  assign _GEN_592 = 6'he == _T_128 ? welem[14] : _GEN_591; // @[Execute.scala 117:10]
  assign _GEN_593 = 6'hf == _T_128 ? welem[15] : _GEN_592; // @[Execute.scala 117:10]
  assign _GEN_594 = 6'h10 == _T_128 ? welem[16] : _GEN_593; // @[Execute.scala 117:10]
  assign _GEN_595 = 6'h11 == _T_128 ? welem[17] : _GEN_594; // @[Execute.scala 117:10]
  assign _GEN_596 = 6'h12 == _T_128 ? welem[18] : _GEN_595; // @[Execute.scala 117:10]
  assign _GEN_597 = 6'h13 == _T_128 ? welem[19] : _GEN_596; // @[Execute.scala 117:10]
  assign _GEN_598 = 6'h14 == _T_128 ? welem[20] : _GEN_597; // @[Execute.scala 117:10]
  assign _GEN_599 = 6'h15 == _T_128 ? welem[21] : _GEN_598; // @[Execute.scala 117:10]
  assign _GEN_600 = 6'h16 == _T_128 ? welem[22] : _GEN_599; // @[Execute.scala 117:10]
  assign _GEN_601 = 6'h17 == _T_128 ? welem[23] : _GEN_600; // @[Execute.scala 117:10]
  assign _GEN_602 = 6'h18 == _T_128 ? welem[24] : _GEN_601; // @[Execute.scala 117:10]
  assign _GEN_603 = 6'h19 == _T_128 ? welem[25] : _GEN_602; // @[Execute.scala 117:10]
  assign _GEN_604 = 6'h1a == _T_128 ? welem[26] : _GEN_603; // @[Execute.scala 117:10]
  assign _GEN_605 = 6'h1b == _T_128 ? welem[27] : _GEN_604; // @[Execute.scala 117:10]
  assign _GEN_606 = 6'h1c == _T_128 ? welem[28] : _GEN_605; // @[Execute.scala 117:10]
  assign _GEN_607 = 6'h1d == _T_128 ? welem[29] : _GEN_606; // @[Execute.scala 117:10]
  assign _GEN_608 = 6'h1e == _T_128 ? welem[30] : _GEN_607; // @[Execute.scala 117:10]
  assign _GEN_609 = 6'h1f == _T_128 ? welem[31] : _GEN_608; // @[Execute.scala 117:10]
  assign _GEN_610 = 6'h20 == _T_128 ? welem[32] : _GEN_609; // @[Execute.scala 117:10]
  assign _GEN_611 = 6'h21 == _T_128 ? welem[33] : _GEN_610; // @[Execute.scala 117:10]
  assign _GEN_612 = 6'h22 == _T_128 ? welem[34] : _GEN_611; // @[Execute.scala 117:10]
  assign _GEN_613 = 6'h23 == _T_128 ? welem[35] : _GEN_612; // @[Execute.scala 117:10]
  assign _GEN_614 = 6'h24 == _T_128 ? welem[36] : _GEN_613; // @[Execute.scala 117:10]
  assign _GEN_615 = 6'h25 == _T_128 ? welem[37] : _GEN_614; // @[Execute.scala 117:10]
  assign _GEN_616 = 6'h26 == _T_128 ? welem[38] : _GEN_615; // @[Execute.scala 117:10]
  assign _GEN_617 = 6'h27 == _T_128 ? welem[39] : _GEN_616; // @[Execute.scala 117:10]
  assign _GEN_618 = 6'h28 == _T_128 ? welem[40] : _GEN_617; // @[Execute.scala 117:10]
  assign _GEN_619 = 6'h29 == _T_128 ? welem[41] : _GEN_618; // @[Execute.scala 117:10]
  assign _GEN_620 = 6'h2a == _T_128 ? welem[42] : _GEN_619; // @[Execute.scala 117:10]
  assign _GEN_621 = 6'h2b == _T_128 ? welem[43] : _GEN_620; // @[Execute.scala 117:10]
  assign _GEN_622 = 6'h2c == _T_128 ? welem[44] : _GEN_621; // @[Execute.scala 117:10]
  assign _GEN_623 = 6'h2d == _T_128 ? welem[45] : _GEN_622; // @[Execute.scala 117:10]
  assign _GEN_624 = 6'h2e == _T_128 ? welem[46] : _GEN_623; // @[Execute.scala 117:10]
  assign _GEN_625 = 6'h2f == _T_128 ? welem[47] : _GEN_624; // @[Execute.scala 117:10]
  assign _GEN_626 = 6'h30 == _T_128 ? welem[48] : _GEN_625; // @[Execute.scala 117:10]
  assign _GEN_627 = 6'h31 == _T_128 ? welem[49] : _GEN_626; // @[Execute.scala 117:10]
  assign _GEN_628 = 6'h32 == _T_128 ? welem[50] : _GEN_627; // @[Execute.scala 117:10]
  assign _GEN_629 = 6'h33 == _T_128 ? welem[51] : _GEN_628; // @[Execute.scala 117:10]
  assign _GEN_630 = 6'h34 == _T_128 ? welem[52] : _GEN_629; // @[Execute.scala 117:10]
  assign _GEN_631 = 6'h35 == _T_128 ? welem[53] : _GEN_630; // @[Execute.scala 117:10]
  assign _GEN_632 = 6'h36 == _T_128 ? welem[54] : _GEN_631; // @[Execute.scala 117:10]
  assign _GEN_633 = 6'h37 == _T_128 ? welem[55] : _GEN_632; // @[Execute.scala 117:10]
  assign _GEN_634 = 6'h38 == _T_128 ? welem[56] : _GEN_633; // @[Execute.scala 117:10]
  assign _GEN_635 = 6'h39 == _T_128 ? welem[57] : _GEN_634; // @[Execute.scala 117:10]
  assign _GEN_636 = 6'h3a == _T_128 ? welem[58] : _GEN_635; // @[Execute.scala 117:10]
  assign _GEN_637 = 6'h3b == _T_128 ? welem[59] : _GEN_636; // @[Execute.scala 117:10]
  assign _GEN_638 = 6'h3c == _T_128 ? welem[60] : _GEN_637; // @[Execute.scala 117:10]
  assign _GEN_639 = 6'h3d == _T_128 ? welem[61] : _GEN_638; // @[Execute.scala 117:10]
  assign _GEN_640 = 6'h3e == _T_128 ? welem[62] : _GEN_639; // @[Execute.scala 117:10]
  assign _GEN_641 = 6'h3f == _T_128 ? welem[63] : _GEN_640; // @[Execute.scala 117:10]
  assign _T_131 = _T_122 ? _GEN_577 : _GEN_641; // @[Execute.scala 117:10]
  assign _T_132 = r < 6'h3c; // @[Execute.scala 117:15]
  assign _T_134 = r - 6'h3c; // @[Execute.scala 117:37]
  assign _T_138 = 6'h4 + r; // @[Execute.scala 117:60]
  assign _GEN_643 = 6'h1 == _T_134 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_644 = 6'h2 == _T_134 ? welem[2] : _GEN_643; // @[Execute.scala 117:10]
  assign _GEN_645 = 6'h3 == _T_134 ? welem[3] : _GEN_644; // @[Execute.scala 117:10]
  assign _GEN_646 = 6'h4 == _T_134 ? welem[4] : _GEN_645; // @[Execute.scala 117:10]
  assign _GEN_647 = 6'h5 == _T_134 ? welem[5] : _GEN_646; // @[Execute.scala 117:10]
  assign _GEN_648 = 6'h6 == _T_134 ? welem[6] : _GEN_647; // @[Execute.scala 117:10]
  assign _GEN_649 = 6'h7 == _T_134 ? welem[7] : _GEN_648; // @[Execute.scala 117:10]
  assign _GEN_650 = 6'h8 == _T_134 ? welem[8] : _GEN_649; // @[Execute.scala 117:10]
  assign _GEN_651 = 6'h9 == _T_134 ? welem[9] : _GEN_650; // @[Execute.scala 117:10]
  assign _GEN_652 = 6'ha == _T_134 ? welem[10] : _GEN_651; // @[Execute.scala 117:10]
  assign _GEN_653 = 6'hb == _T_134 ? welem[11] : _GEN_652; // @[Execute.scala 117:10]
  assign _GEN_654 = 6'hc == _T_134 ? welem[12] : _GEN_653; // @[Execute.scala 117:10]
  assign _GEN_655 = 6'hd == _T_134 ? welem[13] : _GEN_654; // @[Execute.scala 117:10]
  assign _GEN_656 = 6'he == _T_134 ? welem[14] : _GEN_655; // @[Execute.scala 117:10]
  assign _GEN_657 = 6'hf == _T_134 ? welem[15] : _GEN_656; // @[Execute.scala 117:10]
  assign _GEN_658 = 6'h10 == _T_134 ? welem[16] : _GEN_657; // @[Execute.scala 117:10]
  assign _GEN_659 = 6'h11 == _T_134 ? welem[17] : _GEN_658; // @[Execute.scala 117:10]
  assign _GEN_660 = 6'h12 == _T_134 ? welem[18] : _GEN_659; // @[Execute.scala 117:10]
  assign _GEN_661 = 6'h13 == _T_134 ? welem[19] : _GEN_660; // @[Execute.scala 117:10]
  assign _GEN_662 = 6'h14 == _T_134 ? welem[20] : _GEN_661; // @[Execute.scala 117:10]
  assign _GEN_663 = 6'h15 == _T_134 ? welem[21] : _GEN_662; // @[Execute.scala 117:10]
  assign _GEN_664 = 6'h16 == _T_134 ? welem[22] : _GEN_663; // @[Execute.scala 117:10]
  assign _GEN_665 = 6'h17 == _T_134 ? welem[23] : _GEN_664; // @[Execute.scala 117:10]
  assign _GEN_666 = 6'h18 == _T_134 ? welem[24] : _GEN_665; // @[Execute.scala 117:10]
  assign _GEN_667 = 6'h19 == _T_134 ? welem[25] : _GEN_666; // @[Execute.scala 117:10]
  assign _GEN_668 = 6'h1a == _T_134 ? welem[26] : _GEN_667; // @[Execute.scala 117:10]
  assign _GEN_669 = 6'h1b == _T_134 ? welem[27] : _GEN_668; // @[Execute.scala 117:10]
  assign _GEN_670 = 6'h1c == _T_134 ? welem[28] : _GEN_669; // @[Execute.scala 117:10]
  assign _GEN_671 = 6'h1d == _T_134 ? welem[29] : _GEN_670; // @[Execute.scala 117:10]
  assign _GEN_672 = 6'h1e == _T_134 ? welem[30] : _GEN_671; // @[Execute.scala 117:10]
  assign _GEN_673 = 6'h1f == _T_134 ? welem[31] : _GEN_672; // @[Execute.scala 117:10]
  assign _GEN_674 = 6'h20 == _T_134 ? welem[32] : _GEN_673; // @[Execute.scala 117:10]
  assign _GEN_675 = 6'h21 == _T_134 ? welem[33] : _GEN_674; // @[Execute.scala 117:10]
  assign _GEN_676 = 6'h22 == _T_134 ? welem[34] : _GEN_675; // @[Execute.scala 117:10]
  assign _GEN_677 = 6'h23 == _T_134 ? welem[35] : _GEN_676; // @[Execute.scala 117:10]
  assign _GEN_678 = 6'h24 == _T_134 ? welem[36] : _GEN_677; // @[Execute.scala 117:10]
  assign _GEN_679 = 6'h25 == _T_134 ? welem[37] : _GEN_678; // @[Execute.scala 117:10]
  assign _GEN_680 = 6'h26 == _T_134 ? welem[38] : _GEN_679; // @[Execute.scala 117:10]
  assign _GEN_681 = 6'h27 == _T_134 ? welem[39] : _GEN_680; // @[Execute.scala 117:10]
  assign _GEN_682 = 6'h28 == _T_134 ? welem[40] : _GEN_681; // @[Execute.scala 117:10]
  assign _GEN_683 = 6'h29 == _T_134 ? welem[41] : _GEN_682; // @[Execute.scala 117:10]
  assign _GEN_684 = 6'h2a == _T_134 ? welem[42] : _GEN_683; // @[Execute.scala 117:10]
  assign _GEN_685 = 6'h2b == _T_134 ? welem[43] : _GEN_684; // @[Execute.scala 117:10]
  assign _GEN_686 = 6'h2c == _T_134 ? welem[44] : _GEN_685; // @[Execute.scala 117:10]
  assign _GEN_687 = 6'h2d == _T_134 ? welem[45] : _GEN_686; // @[Execute.scala 117:10]
  assign _GEN_688 = 6'h2e == _T_134 ? welem[46] : _GEN_687; // @[Execute.scala 117:10]
  assign _GEN_689 = 6'h2f == _T_134 ? welem[47] : _GEN_688; // @[Execute.scala 117:10]
  assign _GEN_690 = 6'h30 == _T_134 ? welem[48] : _GEN_689; // @[Execute.scala 117:10]
  assign _GEN_691 = 6'h31 == _T_134 ? welem[49] : _GEN_690; // @[Execute.scala 117:10]
  assign _GEN_692 = 6'h32 == _T_134 ? welem[50] : _GEN_691; // @[Execute.scala 117:10]
  assign _GEN_693 = 6'h33 == _T_134 ? welem[51] : _GEN_692; // @[Execute.scala 117:10]
  assign _GEN_694 = 6'h34 == _T_134 ? welem[52] : _GEN_693; // @[Execute.scala 117:10]
  assign _GEN_695 = 6'h35 == _T_134 ? welem[53] : _GEN_694; // @[Execute.scala 117:10]
  assign _GEN_696 = 6'h36 == _T_134 ? welem[54] : _GEN_695; // @[Execute.scala 117:10]
  assign _GEN_697 = 6'h37 == _T_134 ? welem[55] : _GEN_696; // @[Execute.scala 117:10]
  assign _GEN_698 = 6'h38 == _T_134 ? welem[56] : _GEN_697; // @[Execute.scala 117:10]
  assign _GEN_699 = 6'h39 == _T_134 ? welem[57] : _GEN_698; // @[Execute.scala 117:10]
  assign _GEN_700 = 6'h3a == _T_134 ? welem[58] : _GEN_699; // @[Execute.scala 117:10]
  assign _GEN_701 = 6'h3b == _T_134 ? welem[59] : _GEN_700; // @[Execute.scala 117:10]
  assign _GEN_702 = 6'h3c == _T_134 ? welem[60] : _GEN_701; // @[Execute.scala 117:10]
  assign _GEN_703 = 6'h3d == _T_134 ? welem[61] : _GEN_702; // @[Execute.scala 117:10]
  assign _GEN_704 = 6'h3e == _T_134 ? welem[62] : _GEN_703; // @[Execute.scala 117:10]
  assign _GEN_705 = 6'h3f == _T_134 ? welem[63] : _GEN_704; // @[Execute.scala 117:10]
  assign _GEN_707 = 6'h1 == _T_138 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_708 = 6'h2 == _T_138 ? welem[2] : _GEN_707; // @[Execute.scala 117:10]
  assign _GEN_709 = 6'h3 == _T_138 ? welem[3] : _GEN_708; // @[Execute.scala 117:10]
  assign _GEN_710 = 6'h4 == _T_138 ? welem[4] : _GEN_709; // @[Execute.scala 117:10]
  assign _GEN_711 = 6'h5 == _T_138 ? welem[5] : _GEN_710; // @[Execute.scala 117:10]
  assign _GEN_712 = 6'h6 == _T_138 ? welem[6] : _GEN_711; // @[Execute.scala 117:10]
  assign _GEN_713 = 6'h7 == _T_138 ? welem[7] : _GEN_712; // @[Execute.scala 117:10]
  assign _GEN_714 = 6'h8 == _T_138 ? welem[8] : _GEN_713; // @[Execute.scala 117:10]
  assign _GEN_715 = 6'h9 == _T_138 ? welem[9] : _GEN_714; // @[Execute.scala 117:10]
  assign _GEN_716 = 6'ha == _T_138 ? welem[10] : _GEN_715; // @[Execute.scala 117:10]
  assign _GEN_717 = 6'hb == _T_138 ? welem[11] : _GEN_716; // @[Execute.scala 117:10]
  assign _GEN_718 = 6'hc == _T_138 ? welem[12] : _GEN_717; // @[Execute.scala 117:10]
  assign _GEN_719 = 6'hd == _T_138 ? welem[13] : _GEN_718; // @[Execute.scala 117:10]
  assign _GEN_720 = 6'he == _T_138 ? welem[14] : _GEN_719; // @[Execute.scala 117:10]
  assign _GEN_721 = 6'hf == _T_138 ? welem[15] : _GEN_720; // @[Execute.scala 117:10]
  assign _GEN_722 = 6'h10 == _T_138 ? welem[16] : _GEN_721; // @[Execute.scala 117:10]
  assign _GEN_723 = 6'h11 == _T_138 ? welem[17] : _GEN_722; // @[Execute.scala 117:10]
  assign _GEN_724 = 6'h12 == _T_138 ? welem[18] : _GEN_723; // @[Execute.scala 117:10]
  assign _GEN_725 = 6'h13 == _T_138 ? welem[19] : _GEN_724; // @[Execute.scala 117:10]
  assign _GEN_726 = 6'h14 == _T_138 ? welem[20] : _GEN_725; // @[Execute.scala 117:10]
  assign _GEN_727 = 6'h15 == _T_138 ? welem[21] : _GEN_726; // @[Execute.scala 117:10]
  assign _GEN_728 = 6'h16 == _T_138 ? welem[22] : _GEN_727; // @[Execute.scala 117:10]
  assign _GEN_729 = 6'h17 == _T_138 ? welem[23] : _GEN_728; // @[Execute.scala 117:10]
  assign _GEN_730 = 6'h18 == _T_138 ? welem[24] : _GEN_729; // @[Execute.scala 117:10]
  assign _GEN_731 = 6'h19 == _T_138 ? welem[25] : _GEN_730; // @[Execute.scala 117:10]
  assign _GEN_732 = 6'h1a == _T_138 ? welem[26] : _GEN_731; // @[Execute.scala 117:10]
  assign _GEN_733 = 6'h1b == _T_138 ? welem[27] : _GEN_732; // @[Execute.scala 117:10]
  assign _GEN_734 = 6'h1c == _T_138 ? welem[28] : _GEN_733; // @[Execute.scala 117:10]
  assign _GEN_735 = 6'h1d == _T_138 ? welem[29] : _GEN_734; // @[Execute.scala 117:10]
  assign _GEN_736 = 6'h1e == _T_138 ? welem[30] : _GEN_735; // @[Execute.scala 117:10]
  assign _GEN_737 = 6'h1f == _T_138 ? welem[31] : _GEN_736; // @[Execute.scala 117:10]
  assign _GEN_738 = 6'h20 == _T_138 ? welem[32] : _GEN_737; // @[Execute.scala 117:10]
  assign _GEN_739 = 6'h21 == _T_138 ? welem[33] : _GEN_738; // @[Execute.scala 117:10]
  assign _GEN_740 = 6'h22 == _T_138 ? welem[34] : _GEN_739; // @[Execute.scala 117:10]
  assign _GEN_741 = 6'h23 == _T_138 ? welem[35] : _GEN_740; // @[Execute.scala 117:10]
  assign _GEN_742 = 6'h24 == _T_138 ? welem[36] : _GEN_741; // @[Execute.scala 117:10]
  assign _GEN_743 = 6'h25 == _T_138 ? welem[37] : _GEN_742; // @[Execute.scala 117:10]
  assign _GEN_744 = 6'h26 == _T_138 ? welem[38] : _GEN_743; // @[Execute.scala 117:10]
  assign _GEN_745 = 6'h27 == _T_138 ? welem[39] : _GEN_744; // @[Execute.scala 117:10]
  assign _GEN_746 = 6'h28 == _T_138 ? welem[40] : _GEN_745; // @[Execute.scala 117:10]
  assign _GEN_747 = 6'h29 == _T_138 ? welem[41] : _GEN_746; // @[Execute.scala 117:10]
  assign _GEN_748 = 6'h2a == _T_138 ? welem[42] : _GEN_747; // @[Execute.scala 117:10]
  assign _GEN_749 = 6'h2b == _T_138 ? welem[43] : _GEN_748; // @[Execute.scala 117:10]
  assign _GEN_750 = 6'h2c == _T_138 ? welem[44] : _GEN_749; // @[Execute.scala 117:10]
  assign _GEN_751 = 6'h2d == _T_138 ? welem[45] : _GEN_750; // @[Execute.scala 117:10]
  assign _GEN_752 = 6'h2e == _T_138 ? welem[46] : _GEN_751; // @[Execute.scala 117:10]
  assign _GEN_753 = 6'h2f == _T_138 ? welem[47] : _GEN_752; // @[Execute.scala 117:10]
  assign _GEN_754 = 6'h30 == _T_138 ? welem[48] : _GEN_753; // @[Execute.scala 117:10]
  assign _GEN_755 = 6'h31 == _T_138 ? welem[49] : _GEN_754; // @[Execute.scala 117:10]
  assign _GEN_756 = 6'h32 == _T_138 ? welem[50] : _GEN_755; // @[Execute.scala 117:10]
  assign _GEN_757 = 6'h33 == _T_138 ? welem[51] : _GEN_756; // @[Execute.scala 117:10]
  assign _GEN_758 = 6'h34 == _T_138 ? welem[52] : _GEN_757; // @[Execute.scala 117:10]
  assign _GEN_759 = 6'h35 == _T_138 ? welem[53] : _GEN_758; // @[Execute.scala 117:10]
  assign _GEN_760 = 6'h36 == _T_138 ? welem[54] : _GEN_759; // @[Execute.scala 117:10]
  assign _GEN_761 = 6'h37 == _T_138 ? welem[55] : _GEN_760; // @[Execute.scala 117:10]
  assign _GEN_762 = 6'h38 == _T_138 ? welem[56] : _GEN_761; // @[Execute.scala 117:10]
  assign _GEN_763 = 6'h39 == _T_138 ? welem[57] : _GEN_762; // @[Execute.scala 117:10]
  assign _GEN_764 = 6'h3a == _T_138 ? welem[58] : _GEN_763; // @[Execute.scala 117:10]
  assign _GEN_765 = 6'h3b == _T_138 ? welem[59] : _GEN_764; // @[Execute.scala 117:10]
  assign _GEN_766 = 6'h3c == _T_138 ? welem[60] : _GEN_765; // @[Execute.scala 117:10]
  assign _GEN_767 = 6'h3d == _T_138 ? welem[61] : _GEN_766; // @[Execute.scala 117:10]
  assign _GEN_768 = 6'h3e == _T_138 ? welem[62] : _GEN_767; // @[Execute.scala 117:10]
  assign _GEN_769 = 6'h3f == _T_138 ? welem[63] : _GEN_768; // @[Execute.scala 117:10]
  assign _T_141 = _T_132 ? _GEN_705 : _GEN_769; // @[Execute.scala 117:10]
  assign _T_142 = r < 6'h3b; // @[Execute.scala 117:15]
  assign _T_144 = r - 6'h3b; // @[Execute.scala 117:37]
  assign _T_148 = 6'h5 + r; // @[Execute.scala 117:60]
  assign _GEN_771 = 6'h1 == _T_144 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_772 = 6'h2 == _T_144 ? welem[2] : _GEN_771; // @[Execute.scala 117:10]
  assign _GEN_773 = 6'h3 == _T_144 ? welem[3] : _GEN_772; // @[Execute.scala 117:10]
  assign _GEN_774 = 6'h4 == _T_144 ? welem[4] : _GEN_773; // @[Execute.scala 117:10]
  assign _GEN_775 = 6'h5 == _T_144 ? welem[5] : _GEN_774; // @[Execute.scala 117:10]
  assign _GEN_776 = 6'h6 == _T_144 ? welem[6] : _GEN_775; // @[Execute.scala 117:10]
  assign _GEN_777 = 6'h7 == _T_144 ? welem[7] : _GEN_776; // @[Execute.scala 117:10]
  assign _GEN_778 = 6'h8 == _T_144 ? welem[8] : _GEN_777; // @[Execute.scala 117:10]
  assign _GEN_779 = 6'h9 == _T_144 ? welem[9] : _GEN_778; // @[Execute.scala 117:10]
  assign _GEN_780 = 6'ha == _T_144 ? welem[10] : _GEN_779; // @[Execute.scala 117:10]
  assign _GEN_781 = 6'hb == _T_144 ? welem[11] : _GEN_780; // @[Execute.scala 117:10]
  assign _GEN_782 = 6'hc == _T_144 ? welem[12] : _GEN_781; // @[Execute.scala 117:10]
  assign _GEN_783 = 6'hd == _T_144 ? welem[13] : _GEN_782; // @[Execute.scala 117:10]
  assign _GEN_784 = 6'he == _T_144 ? welem[14] : _GEN_783; // @[Execute.scala 117:10]
  assign _GEN_785 = 6'hf == _T_144 ? welem[15] : _GEN_784; // @[Execute.scala 117:10]
  assign _GEN_786 = 6'h10 == _T_144 ? welem[16] : _GEN_785; // @[Execute.scala 117:10]
  assign _GEN_787 = 6'h11 == _T_144 ? welem[17] : _GEN_786; // @[Execute.scala 117:10]
  assign _GEN_788 = 6'h12 == _T_144 ? welem[18] : _GEN_787; // @[Execute.scala 117:10]
  assign _GEN_789 = 6'h13 == _T_144 ? welem[19] : _GEN_788; // @[Execute.scala 117:10]
  assign _GEN_790 = 6'h14 == _T_144 ? welem[20] : _GEN_789; // @[Execute.scala 117:10]
  assign _GEN_791 = 6'h15 == _T_144 ? welem[21] : _GEN_790; // @[Execute.scala 117:10]
  assign _GEN_792 = 6'h16 == _T_144 ? welem[22] : _GEN_791; // @[Execute.scala 117:10]
  assign _GEN_793 = 6'h17 == _T_144 ? welem[23] : _GEN_792; // @[Execute.scala 117:10]
  assign _GEN_794 = 6'h18 == _T_144 ? welem[24] : _GEN_793; // @[Execute.scala 117:10]
  assign _GEN_795 = 6'h19 == _T_144 ? welem[25] : _GEN_794; // @[Execute.scala 117:10]
  assign _GEN_796 = 6'h1a == _T_144 ? welem[26] : _GEN_795; // @[Execute.scala 117:10]
  assign _GEN_797 = 6'h1b == _T_144 ? welem[27] : _GEN_796; // @[Execute.scala 117:10]
  assign _GEN_798 = 6'h1c == _T_144 ? welem[28] : _GEN_797; // @[Execute.scala 117:10]
  assign _GEN_799 = 6'h1d == _T_144 ? welem[29] : _GEN_798; // @[Execute.scala 117:10]
  assign _GEN_800 = 6'h1e == _T_144 ? welem[30] : _GEN_799; // @[Execute.scala 117:10]
  assign _GEN_801 = 6'h1f == _T_144 ? welem[31] : _GEN_800; // @[Execute.scala 117:10]
  assign _GEN_802 = 6'h20 == _T_144 ? welem[32] : _GEN_801; // @[Execute.scala 117:10]
  assign _GEN_803 = 6'h21 == _T_144 ? welem[33] : _GEN_802; // @[Execute.scala 117:10]
  assign _GEN_804 = 6'h22 == _T_144 ? welem[34] : _GEN_803; // @[Execute.scala 117:10]
  assign _GEN_805 = 6'h23 == _T_144 ? welem[35] : _GEN_804; // @[Execute.scala 117:10]
  assign _GEN_806 = 6'h24 == _T_144 ? welem[36] : _GEN_805; // @[Execute.scala 117:10]
  assign _GEN_807 = 6'h25 == _T_144 ? welem[37] : _GEN_806; // @[Execute.scala 117:10]
  assign _GEN_808 = 6'h26 == _T_144 ? welem[38] : _GEN_807; // @[Execute.scala 117:10]
  assign _GEN_809 = 6'h27 == _T_144 ? welem[39] : _GEN_808; // @[Execute.scala 117:10]
  assign _GEN_810 = 6'h28 == _T_144 ? welem[40] : _GEN_809; // @[Execute.scala 117:10]
  assign _GEN_811 = 6'h29 == _T_144 ? welem[41] : _GEN_810; // @[Execute.scala 117:10]
  assign _GEN_812 = 6'h2a == _T_144 ? welem[42] : _GEN_811; // @[Execute.scala 117:10]
  assign _GEN_813 = 6'h2b == _T_144 ? welem[43] : _GEN_812; // @[Execute.scala 117:10]
  assign _GEN_814 = 6'h2c == _T_144 ? welem[44] : _GEN_813; // @[Execute.scala 117:10]
  assign _GEN_815 = 6'h2d == _T_144 ? welem[45] : _GEN_814; // @[Execute.scala 117:10]
  assign _GEN_816 = 6'h2e == _T_144 ? welem[46] : _GEN_815; // @[Execute.scala 117:10]
  assign _GEN_817 = 6'h2f == _T_144 ? welem[47] : _GEN_816; // @[Execute.scala 117:10]
  assign _GEN_818 = 6'h30 == _T_144 ? welem[48] : _GEN_817; // @[Execute.scala 117:10]
  assign _GEN_819 = 6'h31 == _T_144 ? welem[49] : _GEN_818; // @[Execute.scala 117:10]
  assign _GEN_820 = 6'h32 == _T_144 ? welem[50] : _GEN_819; // @[Execute.scala 117:10]
  assign _GEN_821 = 6'h33 == _T_144 ? welem[51] : _GEN_820; // @[Execute.scala 117:10]
  assign _GEN_822 = 6'h34 == _T_144 ? welem[52] : _GEN_821; // @[Execute.scala 117:10]
  assign _GEN_823 = 6'h35 == _T_144 ? welem[53] : _GEN_822; // @[Execute.scala 117:10]
  assign _GEN_824 = 6'h36 == _T_144 ? welem[54] : _GEN_823; // @[Execute.scala 117:10]
  assign _GEN_825 = 6'h37 == _T_144 ? welem[55] : _GEN_824; // @[Execute.scala 117:10]
  assign _GEN_826 = 6'h38 == _T_144 ? welem[56] : _GEN_825; // @[Execute.scala 117:10]
  assign _GEN_827 = 6'h39 == _T_144 ? welem[57] : _GEN_826; // @[Execute.scala 117:10]
  assign _GEN_828 = 6'h3a == _T_144 ? welem[58] : _GEN_827; // @[Execute.scala 117:10]
  assign _GEN_829 = 6'h3b == _T_144 ? welem[59] : _GEN_828; // @[Execute.scala 117:10]
  assign _GEN_830 = 6'h3c == _T_144 ? welem[60] : _GEN_829; // @[Execute.scala 117:10]
  assign _GEN_831 = 6'h3d == _T_144 ? welem[61] : _GEN_830; // @[Execute.scala 117:10]
  assign _GEN_832 = 6'h3e == _T_144 ? welem[62] : _GEN_831; // @[Execute.scala 117:10]
  assign _GEN_833 = 6'h3f == _T_144 ? welem[63] : _GEN_832; // @[Execute.scala 117:10]
  assign _GEN_835 = 6'h1 == _T_148 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_836 = 6'h2 == _T_148 ? welem[2] : _GEN_835; // @[Execute.scala 117:10]
  assign _GEN_837 = 6'h3 == _T_148 ? welem[3] : _GEN_836; // @[Execute.scala 117:10]
  assign _GEN_838 = 6'h4 == _T_148 ? welem[4] : _GEN_837; // @[Execute.scala 117:10]
  assign _GEN_839 = 6'h5 == _T_148 ? welem[5] : _GEN_838; // @[Execute.scala 117:10]
  assign _GEN_840 = 6'h6 == _T_148 ? welem[6] : _GEN_839; // @[Execute.scala 117:10]
  assign _GEN_841 = 6'h7 == _T_148 ? welem[7] : _GEN_840; // @[Execute.scala 117:10]
  assign _GEN_842 = 6'h8 == _T_148 ? welem[8] : _GEN_841; // @[Execute.scala 117:10]
  assign _GEN_843 = 6'h9 == _T_148 ? welem[9] : _GEN_842; // @[Execute.scala 117:10]
  assign _GEN_844 = 6'ha == _T_148 ? welem[10] : _GEN_843; // @[Execute.scala 117:10]
  assign _GEN_845 = 6'hb == _T_148 ? welem[11] : _GEN_844; // @[Execute.scala 117:10]
  assign _GEN_846 = 6'hc == _T_148 ? welem[12] : _GEN_845; // @[Execute.scala 117:10]
  assign _GEN_847 = 6'hd == _T_148 ? welem[13] : _GEN_846; // @[Execute.scala 117:10]
  assign _GEN_848 = 6'he == _T_148 ? welem[14] : _GEN_847; // @[Execute.scala 117:10]
  assign _GEN_849 = 6'hf == _T_148 ? welem[15] : _GEN_848; // @[Execute.scala 117:10]
  assign _GEN_850 = 6'h10 == _T_148 ? welem[16] : _GEN_849; // @[Execute.scala 117:10]
  assign _GEN_851 = 6'h11 == _T_148 ? welem[17] : _GEN_850; // @[Execute.scala 117:10]
  assign _GEN_852 = 6'h12 == _T_148 ? welem[18] : _GEN_851; // @[Execute.scala 117:10]
  assign _GEN_853 = 6'h13 == _T_148 ? welem[19] : _GEN_852; // @[Execute.scala 117:10]
  assign _GEN_854 = 6'h14 == _T_148 ? welem[20] : _GEN_853; // @[Execute.scala 117:10]
  assign _GEN_855 = 6'h15 == _T_148 ? welem[21] : _GEN_854; // @[Execute.scala 117:10]
  assign _GEN_856 = 6'h16 == _T_148 ? welem[22] : _GEN_855; // @[Execute.scala 117:10]
  assign _GEN_857 = 6'h17 == _T_148 ? welem[23] : _GEN_856; // @[Execute.scala 117:10]
  assign _GEN_858 = 6'h18 == _T_148 ? welem[24] : _GEN_857; // @[Execute.scala 117:10]
  assign _GEN_859 = 6'h19 == _T_148 ? welem[25] : _GEN_858; // @[Execute.scala 117:10]
  assign _GEN_860 = 6'h1a == _T_148 ? welem[26] : _GEN_859; // @[Execute.scala 117:10]
  assign _GEN_861 = 6'h1b == _T_148 ? welem[27] : _GEN_860; // @[Execute.scala 117:10]
  assign _GEN_862 = 6'h1c == _T_148 ? welem[28] : _GEN_861; // @[Execute.scala 117:10]
  assign _GEN_863 = 6'h1d == _T_148 ? welem[29] : _GEN_862; // @[Execute.scala 117:10]
  assign _GEN_864 = 6'h1e == _T_148 ? welem[30] : _GEN_863; // @[Execute.scala 117:10]
  assign _GEN_865 = 6'h1f == _T_148 ? welem[31] : _GEN_864; // @[Execute.scala 117:10]
  assign _GEN_866 = 6'h20 == _T_148 ? welem[32] : _GEN_865; // @[Execute.scala 117:10]
  assign _GEN_867 = 6'h21 == _T_148 ? welem[33] : _GEN_866; // @[Execute.scala 117:10]
  assign _GEN_868 = 6'h22 == _T_148 ? welem[34] : _GEN_867; // @[Execute.scala 117:10]
  assign _GEN_869 = 6'h23 == _T_148 ? welem[35] : _GEN_868; // @[Execute.scala 117:10]
  assign _GEN_870 = 6'h24 == _T_148 ? welem[36] : _GEN_869; // @[Execute.scala 117:10]
  assign _GEN_871 = 6'h25 == _T_148 ? welem[37] : _GEN_870; // @[Execute.scala 117:10]
  assign _GEN_872 = 6'h26 == _T_148 ? welem[38] : _GEN_871; // @[Execute.scala 117:10]
  assign _GEN_873 = 6'h27 == _T_148 ? welem[39] : _GEN_872; // @[Execute.scala 117:10]
  assign _GEN_874 = 6'h28 == _T_148 ? welem[40] : _GEN_873; // @[Execute.scala 117:10]
  assign _GEN_875 = 6'h29 == _T_148 ? welem[41] : _GEN_874; // @[Execute.scala 117:10]
  assign _GEN_876 = 6'h2a == _T_148 ? welem[42] : _GEN_875; // @[Execute.scala 117:10]
  assign _GEN_877 = 6'h2b == _T_148 ? welem[43] : _GEN_876; // @[Execute.scala 117:10]
  assign _GEN_878 = 6'h2c == _T_148 ? welem[44] : _GEN_877; // @[Execute.scala 117:10]
  assign _GEN_879 = 6'h2d == _T_148 ? welem[45] : _GEN_878; // @[Execute.scala 117:10]
  assign _GEN_880 = 6'h2e == _T_148 ? welem[46] : _GEN_879; // @[Execute.scala 117:10]
  assign _GEN_881 = 6'h2f == _T_148 ? welem[47] : _GEN_880; // @[Execute.scala 117:10]
  assign _GEN_882 = 6'h30 == _T_148 ? welem[48] : _GEN_881; // @[Execute.scala 117:10]
  assign _GEN_883 = 6'h31 == _T_148 ? welem[49] : _GEN_882; // @[Execute.scala 117:10]
  assign _GEN_884 = 6'h32 == _T_148 ? welem[50] : _GEN_883; // @[Execute.scala 117:10]
  assign _GEN_885 = 6'h33 == _T_148 ? welem[51] : _GEN_884; // @[Execute.scala 117:10]
  assign _GEN_886 = 6'h34 == _T_148 ? welem[52] : _GEN_885; // @[Execute.scala 117:10]
  assign _GEN_887 = 6'h35 == _T_148 ? welem[53] : _GEN_886; // @[Execute.scala 117:10]
  assign _GEN_888 = 6'h36 == _T_148 ? welem[54] : _GEN_887; // @[Execute.scala 117:10]
  assign _GEN_889 = 6'h37 == _T_148 ? welem[55] : _GEN_888; // @[Execute.scala 117:10]
  assign _GEN_890 = 6'h38 == _T_148 ? welem[56] : _GEN_889; // @[Execute.scala 117:10]
  assign _GEN_891 = 6'h39 == _T_148 ? welem[57] : _GEN_890; // @[Execute.scala 117:10]
  assign _GEN_892 = 6'h3a == _T_148 ? welem[58] : _GEN_891; // @[Execute.scala 117:10]
  assign _GEN_893 = 6'h3b == _T_148 ? welem[59] : _GEN_892; // @[Execute.scala 117:10]
  assign _GEN_894 = 6'h3c == _T_148 ? welem[60] : _GEN_893; // @[Execute.scala 117:10]
  assign _GEN_895 = 6'h3d == _T_148 ? welem[61] : _GEN_894; // @[Execute.scala 117:10]
  assign _GEN_896 = 6'h3e == _T_148 ? welem[62] : _GEN_895; // @[Execute.scala 117:10]
  assign _GEN_897 = 6'h3f == _T_148 ? welem[63] : _GEN_896; // @[Execute.scala 117:10]
  assign _T_151 = _T_142 ? _GEN_833 : _GEN_897; // @[Execute.scala 117:10]
  assign _T_152 = r < 6'h3a; // @[Execute.scala 117:15]
  assign _T_154 = r - 6'h3a; // @[Execute.scala 117:37]
  assign _T_158 = 6'h6 + r; // @[Execute.scala 117:60]
  assign _GEN_899 = 6'h1 == _T_154 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_900 = 6'h2 == _T_154 ? welem[2] : _GEN_899; // @[Execute.scala 117:10]
  assign _GEN_901 = 6'h3 == _T_154 ? welem[3] : _GEN_900; // @[Execute.scala 117:10]
  assign _GEN_902 = 6'h4 == _T_154 ? welem[4] : _GEN_901; // @[Execute.scala 117:10]
  assign _GEN_903 = 6'h5 == _T_154 ? welem[5] : _GEN_902; // @[Execute.scala 117:10]
  assign _GEN_904 = 6'h6 == _T_154 ? welem[6] : _GEN_903; // @[Execute.scala 117:10]
  assign _GEN_905 = 6'h7 == _T_154 ? welem[7] : _GEN_904; // @[Execute.scala 117:10]
  assign _GEN_906 = 6'h8 == _T_154 ? welem[8] : _GEN_905; // @[Execute.scala 117:10]
  assign _GEN_907 = 6'h9 == _T_154 ? welem[9] : _GEN_906; // @[Execute.scala 117:10]
  assign _GEN_908 = 6'ha == _T_154 ? welem[10] : _GEN_907; // @[Execute.scala 117:10]
  assign _GEN_909 = 6'hb == _T_154 ? welem[11] : _GEN_908; // @[Execute.scala 117:10]
  assign _GEN_910 = 6'hc == _T_154 ? welem[12] : _GEN_909; // @[Execute.scala 117:10]
  assign _GEN_911 = 6'hd == _T_154 ? welem[13] : _GEN_910; // @[Execute.scala 117:10]
  assign _GEN_912 = 6'he == _T_154 ? welem[14] : _GEN_911; // @[Execute.scala 117:10]
  assign _GEN_913 = 6'hf == _T_154 ? welem[15] : _GEN_912; // @[Execute.scala 117:10]
  assign _GEN_914 = 6'h10 == _T_154 ? welem[16] : _GEN_913; // @[Execute.scala 117:10]
  assign _GEN_915 = 6'h11 == _T_154 ? welem[17] : _GEN_914; // @[Execute.scala 117:10]
  assign _GEN_916 = 6'h12 == _T_154 ? welem[18] : _GEN_915; // @[Execute.scala 117:10]
  assign _GEN_917 = 6'h13 == _T_154 ? welem[19] : _GEN_916; // @[Execute.scala 117:10]
  assign _GEN_918 = 6'h14 == _T_154 ? welem[20] : _GEN_917; // @[Execute.scala 117:10]
  assign _GEN_919 = 6'h15 == _T_154 ? welem[21] : _GEN_918; // @[Execute.scala 117:10]
  assign _GEN_920 = 6'h16 == _T_154 ? welem[22] : _GEN_919; // @[Execute.scala 117:10]
  assign _GEN_921 = 6'h17 == _T_154 ? welem[23] : _GEN_920; // @[Execute.scala 117:10]
  assign _GEN_922 = 6'h18 == _T_154 ? welem[24] : _GEN_921; // @[Execute.scala 117:10]
  assign _GEN_923 = 6'h19 == _T_154 ? welem[25] : _GEN_922; // @[Execute.scala 117:10]
  assign _GEN_924 = 6'h1a == _T_154 ? welem[26] : _GEN_923; // @[Execute.scala 117:10]
  assign _GEN_925 = 6'h1b == _T_154 ? welem[27] : _GEN_924; // @[Execute.scala 117:10]
  assign _GEN_926 = 6'h1c == _T_154 ? welem[28] : _GEN_925; // @[Execute.scala 117:10]
  assign _GEN_927 = 6'h1d == _T_154 ? welem[29] : _GEN_926; // @[Execute.scala 117:10]
  assign _GEN_928 = 6'h1e == _T_154 ? welem[30] : _GEN_927; // @[Execute.scala 117:10]
  assign _GEN_929 = 6'h1f == _T_154 ? welem[31] : _GEN_928; // @[Execute.scala 117:10]
  assign _GEN_930 = 6'h20 == _T_154 ? welem[32] : _GEN_929; // @[Execute.scala 117:10]
  assign _GEN_931 = 6'h21 == _T_154 ? welem[33] : _GEN_930; // @[Execute.scala 117:10]
  assign _GEN_932 = 6'h22 == _T_154 ? welem[34] : _GEN_931; // @[Execute.scala 117:10]
  assign _GEN_933 = 6'h23 == _T_154 ? welem[35] : _GEN_932; // @[Execute.scala 117:10]
  assign _GEN_934 = 6'h24 == _T_154 ? welem[36] : _GEN_933; // @[Execute.scala 117:10]
  assign _GEN_935 = 6'h25 == _T_154 ? welem[37] : _GEN_934; // @[Execute.scala 117:10]
  assign _GEN_936 = 6'h26 == _T_154 ? welem[38] : _GEN_935; // @[Execute.scala 117:10]
  assign _GEN_937 = 6'h27 == _T_154 ? welem[39] : _GEN_936; // @[Execute.scala 117:10]
  assign _GEN_938 = 6'h28 == _T_154 ? welem[40] : _GEN_937; // @[Execute.scala 117:10]
  assign _GEN_939 = 6'h29 == _T_154 ? welem[41] : _GEN_938; // @[Execute.scala 117:10]
  assign _GEN_940 = 6'h2a == _T_154 ? welem[42] : _GEN_939; // @[Execute.scala 117:10]
  assign _GEN_941 = 6'h2b == _T_154 ? welem[43] : _GEN_940; // @[Execute.scala 117:10]
  assign _GEN_942 = 6'h2c == _T_154 ? welem[44] : _GEN_941; // @[Execute.scala 117:10]
  assign _GEN_943 = 6'h2d == _T_154 ? welem[45] : _GEN_942; // @[Execute.scala 117:10]
  assign _GEN_944 = 6'h2e == _T_154 ? welem[46] : _GEN_943; // @[Execute.scala 117:10]
  assign _GEN_945 = 6'h2f == _T_154 ? welem[47] : _GEN_944; // @[Execute.scala 117:10]
  assign _GEN_946 = 6'h30 == _T_154 ? welem[48] : _GEN_945; // @[Execute.scala 117:10]
  assign _GEN_947 = 6'h31 == _T_154 ? welem[49] : _GEN_946; // @[Execute.scala 117:10]
  assign _GEN_948 = 6'h32 == _T_154 ? welem[50] : _GEN_947; // @[Execute.scala 117:10]
  assign _GEN_949 = 6'h33 == _T_154 ? welem[51] : _GEN_948; // @[Execute.scala 117:10]
  assign _GEN_950 = 6'h34 == _T_154 ? welem[52] : _GEN_949; // @[Execute.scala 117:10]
  assign _GEN_951 = 6'h35 == _T_154 ? welem[53] : _GEN_950; // @[Execute.scala 117:10]
  assign _GEN_952 = 6'h36 == _T_154 ? welem[54] : _GEN_951; // @[Execute.scala 117:10]
  assign _GEN_953 = 6'h37 == _T_154 ? welem[55] : _GEN_952; // @[Execute.scala 117:10]
  assign _GEN_954 = 6'h38 == _T_154 ? welem[56] : _GEN_953; // @[Execute.scala 117:10]
  assign _GEN_955 = 6'h39 == _T_154 ? welem[57] : _GEN_954; // @[Execute.scala 117:10]
  assign _GEN_956 = 6'h3a == _T_154 ? welem[58] : _GEN_955; // @[Execute.scala 117:10]
  assign _GEN_957 = 6'h3b == _T_154 ? welem[59] : _GEN_956; // @[Execute.scala 117:10]
  assign _GEN_958 = 6'h3c == _T_154 ? welem[60] : _GEN_957; // @[Execute.scala 117:10]
  assign _GEN_959 = 6'h3d == _T_154 ? welem[61] : _GEN_958; // @[Execute.scala 117:10]
  assign _GEN_960 = 6'h3e == _T_154 ? welem[62] : _GEN_959; // @[Execute.scala 117:10]
  assign _GEN_961 = 6'h3f == _T_154 ? welem[63] : _GEN_960; // @[Execute.scala 117:10]
  assign _GEN_963 = 6'h1 == _T_158 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_964 = 6'h2 == _T_158 ? welem[2] : _GEN_963; // @[Execute.scala 117:10]
  assign _GEN_965 = 6'h3 == _T_158 ? welem[3] : _GEN_964; // @[Execute.scala 117:10]
  assign _GEN_966 = 6'h4 == _T_158 ? welem[4] : _GEN_965; // @[Execute.scala 117:10]
  assign _GEN_967 = 6'h5 == _T_158 ? welem[5] : _GEN_966; // @[Execute.scala 117:10]
  assign _GEN_968 = 6'h6 == _T_158 ? welem[6] : _GEN_967; // @[Execute.scala 117:10]
  assign _GEN_969 = 6'h7 == _T_158 ? welem[7] : _GEN_968; // @[Execute.scala 117:10]
  assign _GEN_970 = 6'h8 == _T_158 ? welem[8] : _GEN_969; // @[Execute.scala 117:10]
  assign _GEN_971 = 6'h9 == _T_158 ? welem[9] : _GEN_970; // @[Execute.scala 117:10]
  assign _GEN_972 = 6'ha == _T_158 ? welem[10] : _GEN_971; // @[Execute.scala 117:10]
  assign _GEN_973 = 6'hb == _T_158 ? welem[11] : _GEN_972; // @[Execute.scala 117:10]
  assign _GEN_974 = 6'hc == _T_158 ? welem[12] : _GEN_973; // @[Execute.scala 117:10]
  assign _GEN_975 = 6'hd == _T_158 ? welem[13] : _GEN_974; // @[Execute.scala 117:10]
  assign _GEN_976 = 6'he == _T_158 ? welem[14] : _GEN_975; // @[Execute.scala 117:10]
  assign _GEN_977 = 6'hf == _T_158 ? welem[15] : _GEN_976; // @[Execute.scala 117:10]
  assign _GEN_978 = 6'h10 == _T_158 ? welem[16] : _GEN_977; // @[Execute.scala 117:10]
  assign _GEN_979 = 6'h11 == _T_158 ? welem[17] : _GEN_978; // @[Execute.scala 117:10]
  assign _GEN_980 = 6'h12 == _T_158 ? welem[18] : _GEN_979; // @[Execute.scala 117:10]
  assign _GEN_981 = 6'h13 == _T_158 ? welem[19] : _GEN_980; // @[Execute.scala 117:10]
  assign _GEN_982 = 6'h14 == _T_158 ? welem[20] : _GEN_981; // @[Execute.scala 117:10]
  assign _GEN_983 = 6'h15 == _T_158 ? welem[21] : _GEN_982; // @[Execute.scala 117:10]
  assign _GEN_984 = 6'h16 == _T_158 ? welem[22] : _GEN_983; // @[Execute.scala 117:10]
  assign _GEN_985 = 6'h17 == _T_158 ? welem[23] : _GEN_984; // @[Execute.scala 117:10]
  assign _GEN_986 = 6'h18 == _T_158 ? welem[24] : _GEN_985; // @[Execute.scala 117:10]
  assign _GEN_987 = 6'h19 == _T_158 ? welem[25] : _GEN_986; // @[Execute.scala 117:10]
  assign _GEN_988 = 6'h1a == _T_158 ? welem[26] : _GEN_987; // @[Execute.scala 117:10]
  assign _GEN_989 = 6'h1b == _T_158 ? welem[27] : _GEN_988; // @[Execute.scala 117:10]
  assign _GEN_990 = 6'h1c == _T_158 ? welem[28] : _GEN_989; // @[Execute.scala 117:10]
  assign _GEN_991 = 6'h1d == _T_158 ? welem[29] : _GEN_990; // @[Execute.scala 117:10]
  assign _GEN_992 = 6'h1e == _T_158 ? welem[30] : _GEN_991; // @[Execute.scala 117:10]
  assign _GEN_993 = 6'h1f == _T_158 ? welem[31] : _GEN_992; // @[Execute.scala 117:10]
  assign _GEN_994 = 6'h20 == _T_158 ? welem[32] : _GEN_993; // @[Execute.scala 117:10]
  assign _GEN_995 = 6'h21 == _T_158 ? welem[33] : _GEN_994; // @[Execute.scala 117:10]
  assign _GEN_996 = 6'h22 == _T_158 ? welem[34] : _GEN_995; // @[Execute.scala 117:10]
  assign _GEN_997 = 6'h23 == _T_158 ? welem[35] : _GEN_996; // @[Execute.scala 117:10]
  assign _GEN_998 = 6'h24 == _T_158 ? welem[36] : _GEN_997; // @[Execute.scala 117:10]
  assign _GEN_999 = 6'h25 == _T_158 ? welem[37] : _GEN_998; // @[Execute.scala 117:10]
  assign _GEN_1000 = 6'h26 == _T_158 ? welem[38] : _GEN_999; // @[Execute.scala 117:10]
  assign _GEN_1001 = 6'h27 == _T_158 ? welem[39] : _GEN_1000; // @[Execute.scala 117:10]
  assign _GEN_1002 = 6'h28 == _T_158 ? welem[40] : _GEN_1001; // @[Execute.scala 117:10]
  assign _GEN_1003 = 6'h29 == _T_158 ? welem[41] : _GEN_1002; // @[Execute.scala 117:10]
  assign _GEN_1004 = 6'h2a == _T_158 ? welem[42] : _GEN_1003; // @[Execute.scala 117:10]
  assign _GEN_1005 = 6'h2b == _T_158 ? welem[43] : _GEN_1004; // @[Execute.scala 117:10]
  assign _GEN_1006 = 6'h2c == _T_158 ? welem[44] : _GEN_1005; // @[Execute.scala 117:10]
  assign _GEN_1007 = 6'h2d == _T_158 ? welem[45] : _GEN_1006; // @[Execute.scala 117:10]
  assign _GEN_1008 = 6'h2e == _T_158 ? welem[46] : _GEN_1007; // @[Execute.scala 117:10]
  assign _GEN_1009 = 6'h2f == _T_158 ? welem[47] : _GEN_1008; // @[Execute.scala 117:10]
  assign _GEN_1010 = 6'h30 == _T_158 ? welem[48] : _GEN_1009; // @[Execute.scala 117:10]
  assign _GEN_1011 = 6'h31 == _T_158 ? welem[49] : _GEN_1010; // @[Execute.scala 117:10]
  assign _GEN_1012 = 6'h32 == _T_158 ? welem[50] : _GEN_1011; // @[Execute.scala 117:10]
  assign _GEN_1013 = 6'h33 == _T_158 ? welem[51] : _GEN_1012; // @[Execute.scala 117:10]
  assign _GEN_1014 = 6'h34 == _T_158 ? welem[52] : _GEN_1013; // @[Execute.scala 117:10]
  assign _GEN_1015 = 6'h35 == _T_158 ? welem[53] : _GEN_1014; // @[Execute.scala 117:10]
  assign _GEN_1016 = 6'h36 == _T_158 ? welem[54] : _GEN_1015; // @[Execute.scala 117:10]
  assign _GEN_1017 = 6'h37 == _T_158 ? welem[55] : _GEN_1016; // @[Execute.scala 117:10]
  assign _GEN_1018 = 6'h38 == _T_158 ? welem[56] : _GEN_1017; // @[Execute.scala 117:10]
  assign _GEN_1019 = 6'h39 == _T_158 ? welem[57] : _GEN_1018; // @[Execute.scala 117:10]
  assign _GEN_1020 = 6'h3a == _T_158 ? welem[58] : _GEN_1019; // @[Execute.scala 117:10]
  assign _GEN_1021 = 6'h3b == _T_158 ? welem[59] : _GEN_1020; // @[Execute.scala 117:10]
  assign _GEN_1022 = 6'h3c == _T_158 ? welem[60] : _GEN_1021; // @[Execute.scala 117:10]
  assign _GEN_1023 = 6'h3d == _T_158 ? welem[61] : _GEN_1022; // @[Execute.scala 117:10]
  assign _GEN_1024 = 6'h3e == _T_158 ? welem[62] : _GEN_1023; // @[Execute.scala 117:10]
  assign _GEN_1025 = 6'h3f == _T_158 ? welem[63] : _GEN_1024; // @[Execute.scala 117:10]
  assign _T_161 = _T_152 ? _GEN_961 : _GEN_1025; // @[Execute.scala 117:10]
  assign _T_162 = r < 6'h39; // @[Execute.scala 117:15]
  assign _T_164 = r - 6'h39; // @[Execute.scala 117:37]
  assign _T_168 = 6'h7 + r; // @[Execute.scala 117:60]
  assign _GEN_1027 = 6'h1 == _T_164 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1028 = 6'h2 == _T_164 ? welem[2] : _GEN_1027; // @[Execute.scala 117:10]
  assign _GEN_1029 = 6'h3 == _T_164 ? welem[3] : _GEN_1028; // @[Execute.scala 117:10]
  assign _GEN_1030 = 6'h4 == _T_164 ? welem[4] : _GEN_1029; // @[Execute.scala 117:10]
  assign _GEN_1031 = 6'h5 == _T_164 ? welem[5] : _GEN_1030; // @[Execute.scala 117:10]
  assign _GEN_1032 = 6'h6 == _T_164 ? welem[6] : _GEN_1031; // @[Execute.scala 117:10]
  assign _GEN_1033 = 6'h7 == _T_164 ? welem[7] : _GEN_1032; // @[Execute.scala 117:10]
  assign _GEN_1034 = 6'h8 == _T_164 ? welem[8] : _GEN_1033; // @[Execute.scala 117:10]
  assign _GEN_1035 = 6'h9 == _T_164 ? welem[9] : _GEN_1034; // @[Execute.scala 117:10]
  assign _GEN_1036 = 6'ha == _T_164 ? welem[10] : _GEN_1035; // @[Execute.scala 117:10]
  assign _GEN_1037 = 6'hb == _T_164 ? welem[11] : _GEN_1036; // @[Execute.scala 117:10]
  assign _GEN_1038 = 6'hc == _T_164 ? welem[12] : _GEN_1037; // @[Execute.scala 117:10]
  assign _GEN_1039 = 6'hd == _T_164 ? welem[13] : _GEN_1038; // @[Execute.scala 117:10]
  assign _GEN_1040 = 6'he == _T_164 ? welem[14] : _GEN_1039; // @[Execute.scala 117:10]
  assign _GEN_1041 = 6'hf == _T_164 ? welem[15] : _GEN_1040; // @[Execute.scala 117:10]
  assign _GEN_1042 = 6'h10 == _T_164 ? welem[16] : _GEN_1041; // @[Execute.scala 117:10]
  assign _GEN_1043 = 6'h11 == _T_164 ? welem[17] : _GEN_1042; // @[Execute.scala 117:10]
  assign _GEN_1044 = 6'h12 == _T_164 ? welem[18] : _GEN_1043; // @[Execute.scala 117:10]
  assign _GEN_1045 = 6'h13 == _T_164 ? welem[19] : _GEN_1044; // @[Execute.scala 117:10]
  assign _GEN_1046 = 6'h14 == _T_164 ? welem[20] : _GEN_1045; // @[Execute.scala 117:10]
  assign _GEN_1047 = 6'h15 == _T_164 ? welem[21] : _GEN_1046; // @[Execute.scala 117:10]
  assign _GEN_1048 = 6'h16 == _T_164 ? welem[22] : _GEN_1047; // @[Execute.scala 117:10]
  assign _GEN_1049 = 6'h17 == _T_164 ? welem[23] : _GEN_1048; // @[Execute.scala 117:10]
  assign _GEN_1050 = 6'h18 == _T_164 ? welem[24] : _GEN_1049; // @[Execute.scala 117:10]
  assign _GEN_1051 = 6'h19 == _T_164 ? welem[25] : _GEN_1050; // @[Execute.scala 117:10]
  assign _GEN_1052 = 6'h1a == _T_164 ? welem[26] : _GEN_1051; // @[Execute.scala 117:10]
  assign _GEN_1053 = 6'h1b == _T_164 ? welem[27] : _GEN_1052; // @[Execute.scala 117:10]
  assign _GEN_1054 = 6'h1c == _T_164 ? welem[28] : _GEN_1053; // @[Execute.scala 117:10]
  assign _GEN_1055 = 6'h1d == _T_164 ? welem[29] : _GEN_1054; // @[Execute.scala 117:10]
  assign _GEN_1056 = 6'h1e == _T_164 ? welem[30] : _GEN_1055; // @[Execute.scala 117:10]
  assign _GEN_1057 = 6'h1f == _T_164 ? welem[31] : _GEN_1056; // @[Execute.scala 117:10]
  assign _GEN_1058 = 6'h20 == _T_164 ? welem[32] : _GEN_1057; // @[Execute.scala 117:10]
  assign _GEN_1059 = 6'h21 == _T_164 ? welem[33] : _GEN_1058; // @[Execute.scala 117:10]
  assign _GEN_1060 = 6'h22 == _T_164 ? welem[34] : _GEN_1059; // @[Execute.scala 117:10]
  assign _GEN_1061 = 6'h23 == _T_164 ? welem[35] : _GEN_1060; // @[Execute.scala 117:10]
  assign _GEN_1062 = 6'h24 == _T_164 ? welem[36] : _GEN_1061; // @[Execute.scala 117:10]
  assign _GEN_1063 = 6'h25 == _T_164 ? welem[37] : _GEN_1062; // @[Execute.scala 117:10]
  assign _GEN_1064 = 6'h26 == _T_164 ? welem[38] : _GEN_1063; // @[Execute.scala 117:10]
  assign _GEN_1065 = 6'h27 == _T_164 ? welem[39] : _GEN_1064; // @[Execute.scala 117:10]
  assign _GEN_1066 = 6'h28 == _T_164 ? welem[40] : _GEN_1065; // @[Execute.scala 117:10]
  assign _GEN_1067 = 6'h29 == _T_164 ? welem[41] : _GEN_1066; // @[Execute.scala 117:10]
  assign _GEN_1068 = 6'h2a == _T_164 ? welem[42] : _GEN_1067; // @[Execute.scala 117:10]
  assign _GEN_1069 = 6'h2b == _T_164 ? welem[43] : _GEN_1068; // @[Execute.scala 117:10]
  assign _GEN_1070 = 6'h2c == _T_164 ? welem[44] : _GEN_1069; // @[Execute.scala 117:10]
  assign _GEN_1071 = 6'h2d == _T_164 ? welem[45] : _GEN_1070; // @[Execute.scala 117:10]
  assign _GEN_1072 = 6'h2e == _T_164 ? welem[46] : _GEN_1071; // @[Execute.scala 117:10]
  assign _GEN_1073 = 6'h2f == _T_164 ? welem[47] : _GEN_1072; // @[Execute.scala 117:10]
  assign _GEN_1074 = 6'h30 == _T_164 ? welem[48] : _GEN_1073; // @[Execute.scala 117:10]
  assign _GEN_1075 = 6'h31 == _T_164 ? welem[49] : _GEN_1074; // @[Execute.scala 117:10]
  assign _GEN_1076 = 6'h32 == _T_164 ? welem[50] : _GEN_1075; // @[Execute.scala 117:10]
  assign _GEN_1077 = 6'h33 == _T_164 ? welem[51] : _GEN_1076; // @[Execute.scala 117:10]
  assign _GEN_1078 = 6'h34 == _T_164 ? welem[52] : _GEN_1077; // @[Execute.scala 117:10]
  assign _GEN_1079 = 6'h35 == _T_164 ? welem[53] : _GEN_1078; // @[Execute.scala 117:10]
  assign _GEN_1080 = 6'h36 == _T_164 ? welem[54] : _GEN_1079; // @[Execute.scala 117:10]
  assign _GEN_1081 = 6'h37 == _T_164 ? welem[55] : _GEN_1080; // @[Execute.scala 117:10]
  assign _GEN_1082 = 6'h38 == _T_164 ? welem[56] : _GEN_1081; // @[Execute.scala 117:10]
  assign _GEN_1083 = 6'h39 == _T_164 ? welem[57] : _GEN_1082; // @[Execute.scala 117:10]
  assign _GEN_1084 = 6'h3a == _T_164 ? welem[58] : _GEN_1083; // @[Execute.scala 117:10]
  assign _GEN_1085 = 6'h3b == _T_164 ? welem[59] : _GEN_1084; // @[Execute.scala 117:10]
  assign _GEN_1086 = 6'h3c == _T_164 ? welem[60] : _GEN_1085; // @[Execute.scala 117:10]
  assign _GEN_1087 = 6'h3d == _T_164 ? welem[61] : _GEN_1086; // @[Execute.scala 117:10]
  assign _GEN_1088 = 6'h3e == _T_164 ? welem[62] : _GEN_1087; // @[Execute.scala 117:10]
  assign _GEN_1089 = 6'h3f == _T_164 ? welem[63] : _GEN_1088; // @[Execute.scala 117:10]
  assign _GEN_1091 = 6'h1 == _T_168 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1092 = 6'h2 == _T_168 ? welem[2] : _GEN_1091; // @[Execute.scala 117:10]
  assign _GEN_1093 = 6'h3 == _T_168 ? welem[3] : _GEN_1092; // @[Execute.scala 117:10]
  assign _GEN_1094 = 6'h4 == _T_168 ? welem[4] : _GEN_1093; // @[Execute.scala 117:10]
  assign _GEN_1095 = 6'h5 == _T_168 ? welem[5] : _GEN_1094; // @[Execute.scala 117:10]
  assign _GEN_1096 = 6'h6 == _T_168 ? welem[6] : _GEN_1095; // @[Execute.scala 117:10]
  assign _GEN_1097 = 6'h7 == _T_168 ? welem[7] : _GEN_1096; // @[Execute.scala 117:10]
  assign _GEN_1098 = 6'h8 == _T_168 ? welem[8] : _GEN_1097; // @[Execute.scala 117:10]
  assign _GEN_1099 = 6'h9 == _T_168 ? welem[9] : _GEN_1098; // @[Execute.scala 117:10]
  assign _GEN_1100 = 6'ha == _T_168 ? welem[10] : _GEN_1099; // @[Execute.scala 117:10]
  assign _GEN_1101 = 6'hb == _T_168 ? welem[11] : _GEN_1100; // @[Execute.scala 117:10]
  assign _GEN_1102 = 6'hc == _T_168 ? welem[12] : _GEN_1101; // @[Execute.scala 117:10]
  assign _GEN_1103 = 6'hd == _T_168 ? welem[13] : _GEN_1102; // @[Execute.scala 117:10]
  assign _GEN_1104 = 6'he == _T_168 ? welem[14] : _GEN_1103; // @[Execute.scala 117:10]
  assign _GEN_1105 = 6'hf == _T_168 ? welem[15] : _GEN_1104; // @[Execute.scala 117:10]
  assign _GEN_1106 = 6'h10 == _T_168 ? welem[16] : _GEN_1105; // @[Execute.scala 117:10]
  assign _GEN_1107 = 6'h11 == _T_168 ? welem[17] : _GEN_1106; // @[Execute.scala 117:10]
  assign _GEN_1108 = 6'h12 == _T_168 ? welem[18] : _GEN_1107; // @[Execute.scala 117:10]
  assign _GEN_1109 = 6'h13 == _T_168 ? welem[19] : _GEN_1108; // @[Execute.scala 117:10]
  assign _GEN_1110 = 6'h14 == _T_168 ? welem[20] : _GEN_1109; // @[Execute.scala 117:10]
  assign _GEN_1111 = 6'h15 == _T_168 ? welem[21] : _GEN_1110; // @[Execute.scala 117:10]
  assign _GEN_1112 = 6'h16 == _T_168 ? welem[22] : _GEN_1111; // @[Execute.scala 117:10]
  assign _GEN_1113 = 6'h17 == _T_168 ? welem[23] : _GEN_1112; // @[Execute.scala 117:10]
  assign _GEN_1114 = 6'h18 == _T_168 ? welem[24] : _GEN_1113; // @[Execute.scala 117:10]
  assign _GEN_1115 = 6'h19 == _T_168 ? welem[25] : _GEN_1114; // @[Execute.scala 117:10]
  assign _GEN_1116 = 6'h1a == _T_168 ? welem[26] : _GEN_1115; // @[Execute.scala 117:10]
  assign _GEN_1117 = 6'h1b == _T_168 ? welem[27] : _GEN_1116; // @[Execute.scala 117:10]
  assign _GEN_1118 = 6'h1c == _T_168 ? welem[28] : _GEN_1117; // @[Execute.scala 117:10]
  assign _GEN_1119 = 6'h1d == _T_168 ? welem[29] : _GEN_1118; // @[Execute.scala 117:10]
  assign _GEN_1120 = 6'h1e == _T_168 ? welem[30] : _GEN_1119; // @[Execute.scala 117:10]
  assign _GEN_1121 = 6'h1f == _T_168 ? welem[31] : _GEN_1120; // @[Execute.scala 117:10]
  assign _GEN_1122 = 6'h20 == _T_168 ? welem[32] : _GEN_1121; // @[Execute.scala 117:10]
  assign _GEN_1123 = 6'h21 == _T_168 ? welem[33] : _GEN_1122; // @[Execute.scala 117:10]
  assign _GEN_1124 = 6'h22 == _T_168 ? welem[34] : _GEN_1123; // @[Execute.scala 117:10]
  assign _GEN_1125 = 6'h23 == _T_168 ? welem[35] : _GEN_1124; // @[Execute.scala 117:10]
  assign _GEN_1126 = 6'h24 == _T_168 ? welem[36] : _GEN_1125; // @[Execute.scala 117:10]
  assign _GEN_1127 = 6'h25 == _T_168 ? welem[37] : _GEN_1126; // @[Execute.scala 117:10]
  assign _GEN_1128 = 6'h26 == _T_168 ? welem[38] : _GEN_1127; // @[Execute.scala 117:10]
  assign _GEN_1129 = 6'h27 == _T_168 ? welem[39] : _GEN_1128; // @[Execute.scala 117:10]
  assign _GEN_1130 = 6'h28 == _T_168 ? welem[40] : _GEN_1129; // @[Execute.scala 117:10]
  assign _GEN_1131 = 6'h29 == _T_168 ? welem[41] : _GEN_1130; // @[Execute.scala 117:10]
  assign _GEN_1132 = 6'h2a == _T_168 ? welem[42] : _GEN_1131; // @[Execute.scala 117:10]
  assign _GEN_1133 = 6'h2b == _T_168 ? welem[43] : _GEN_1132; // @[Execute.scala 117:10]
  assign _GEN_1134 = 6'h2c == _T_168 ? welem[44] : _GEN_1133; // @[Execute.scala 117:10]
  assign _GEN_1135 = 6'h2d == _T_168 ? welem[45] : _GEN_1134; // @[Execute.scala 117:10]
  assign _GEN_1136 = 6'h2e == _T_168 ? welem[46] : _GEN_1135; // @[Execute.scala 117:10]
  assign _GEN_1137 = 6'h2f == _T_168 ? welem[47] : _GEN_1136; // @[Execute.scala 117:10]
  assign _GEN_1138 = 6'h30 == _T_168 ? welem[48] : _GEN_1137; // @[Execute.scala 117:10]
  assign _GEN_1139 = 6'h31 == _T_168 ? welem[49] : _GEN_1138; // @[Execute.scala 117:10]
  assign _GEN_1140 = 6'h32 == _T_168 ? welem[50] : _GEN_1139; // @[Execute.scala 117:10]
  assign _GEN_1141 = 6'h33 == _T_168 ? welem[51] : _GEN_1140; // @[Execute.scala 117:10]
  assign _GEN_1142 = 6'h34 == _T_168 ? welem[52] : _GEN_1141; // @[Execute.scala 117:10]
  assign _GEN_1143 = 6'h35 == _T_168 ? welem[53] : _GEN_1142; // @[Execute.scala 117:10]
  assign _GEN_1144 = 6'h36 == _T_168 ? welem[54] : _GEN_1143; // @[Execute.scala 117:10]
  assign _GEN_1145 = 6'h37 == _T_168 ? welem[55] : _GEN_1144; // @[Execute.scala 117:10]
  assign _GEN_1146 = 6'h38 == _T_168 ? welem[56] : _GEN_1145; // @[Execute.scala 117:10]
  assign _GEN_1147 = 6'h39 == _T_168 ? welem[57] : _GEN_1146; // @[Execute.scala 117:10]
  assign _GEN_1148 = 6'h3a == _T_168 ? welem[58] : _GEN_1147; // @[Execute.scala 117:10]
  assign _GEN_1149 = 6'h3b == _T_168 ? welem[59] : _GEN_1148; // @[Execute.scala 117:10]
  assign _GEN_1150 = 6'h3c == _T_168 ? welem[60] : _GEN_1149; // @[Execute.scala 117:10]
  assign _GEN_1151 = 6'h3d == _T_168 ? welem[61] : _GEN_1150; // @[Execute.scala 117:10]
  assign _GEN_1152 = 6'h3e == _T_168 ? welem[62] : _GEN_1151; // @[Execute.scala 117:10]
  assign _GEN_1153 = 6'h3f == _T_168 ? welem[63] : _GEN_1152; // @[Execute.scala 117:10]
  assign _T_171 = _T_162 ? _GEN_1089 : _GEN_1153; // @[Execute.scala 117:10]
  assign _T_172 = r < 6'h38; // @[Execute.scala 117:15]
  assign _T_174 = r - 6'h38; // @[Execute.scala 117:37]
  assign _T_178 = 6'h8 + r; // @[Execute.scala 117:60]
  assign _GEN_1155 = 6'h1 == _T_174 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1156 = 6'h2 == _T_174 ? welem[2] : _GEN_1155; // @[Execute.scala 117:10]
  assign _GEN_1157 = 6'h3 == _T_174 ? welem[3] : _GEN_1156; // @[Execute.scala 117:10]
  assign _GEN_1158 = 6'h4 == _T_174 ? welem[4] : _GEN_1157; // @[Execute.scala 117:10]
  assign _GEN_1159 = 6'h5 == _T_174 ? welem[5] : _GEN_1158; // @[Execute.scala 117:10]
  assign _GEN_1160 = 6'h6 == _T_174 ? welem[6] : _GEN_1159; // @[Execute.scala 117:10]
  assign _GEN_1161 = 6'h7 == _T_174 ? welem[7] : _GEN_1160; // @[Execute.scala 117:10]
  assign _GEN_1162 = 6'h8 == _T_174 ? welem[8] : _GEN_1161; // @[Execute.scala 117:10]
  assign _GEN_1163 = 6'h9 == _T_174 ? welem[9] : _GEN_1162; // @[Execute.scala 117:10]
  assign _GEN_1164 = 6'ha == _T_174 ? welem[10] : _GEN_1163; // @[Execute.scala 117:10]
  assign _GEN_1165 = 6'hb == _T_174 ? welem[11] : _GEN_1164; // @[Execute.scala 117:10]
  assign _GEN_1166 = 6'hc == _T_174 ? welem[12] : _GEN_1165; // @[Execute.scala 117:10]
  assign _GEN_1167 = 6'hd == _T_174 ? welem[13] : _GEN_1166; // @[Execute.scala 117:10]
  assign _GEN_1168 = 6'he == _T_174 ? welem[14] : _GEN_1167; // @[Execute.scala 117:10]
  assign _GEN_1169 = 6'hf == _T_174 ? welem[15] : _GEN_1168; // @[Execute.scala 117:10]
  assign _GEN_1170 = 6'h10 == _T_174 ? welem[16] : _GEN_1169; // @[Execute.scala 117:10]
  assign _GEN_1171 = 6'h11 == _T_174 ? welem[17] : _GEN_1170; // @[Execute.scala 117:10]
  assign _GEN_1172 = 6'h12 == _T_174 ? welem[18] : _GEN_1171; // @[Execute.scala 117:10]
  assign _GEN_1173 = 6'h13 == _T_174 ? welem[19] : _GEN_1172; // @[Execute.scala 117:10]
  assign _GEN_1174 = 6'h14 == _T_174 ? welem[20] : _GEN_1173; // @[Execute.scala 117:10]
  assign _GEN_1175 = 6'h15 == _T_174 ? welem[21] : _GEN_1174; // @[Execute.scala 117:10]
  assign _GEN_1176 = 6'h16 == _T_174 ? welem[22] : _GEN_1175; // @[Execute.scala 117:10]
  assign _GEN_1177 = 6'h17 == _T_174 ? welem[23] : _GEN_1176; // @[Execute.scala 117:10]
  assign _GEN_1178 = 6'h18 == _T_174 ? welem[24] : _GEN_1177; // @[Execute.scala 117:10]
  assign _GEN_1179 = 6'h19 == _T_174 ? welem[25] : _GEN_1178; // @[Execute.scala 117:10]
  assign _GEN_1180 = 6'h1a == _T_174 ? welem[26] : _GEN_1179; // @[Execute.scala 117:10]
  assign _GEN_1181 = 6'h1b == _T_174 ? welem[27] : _GEN_1180; // @[Execute.scala 117:10]
  assign _GEN_1182 = 6'h1c == _T_174 ? welem[28] : _GEN_1181; // @[Execute.scala 117:10]
  assign _GEN_1183 = 6'h1d == _T_174 ? welem[29] : _GEN_1182; // @[Execute.scala 117:10]
  assign _GEN_1184 = 6'h1e == _T_174 ? welem[30] : _GEN_1183; // @[Execute.scala 117:10]
  assign _GEN_1185 = 6'h1f == _T_174 ? welem[31] : _GEN_1184; // @[Execute.scala 117:10]
  assign _GEN_1186 = 6'h20 == _T_174 ? welem[32] : _GEN_1185; // @[Execute.scala 117:10]
  assign _GEN_1187 = 6'h21 == _T_174 ? welem[33] : _GEN_1186; // @[Execute.scala 117:10]
  assign _GEN_1188 = 6'h22 == _T_174 ? welem[34] : _GEN_1187; // @[Execute.scala 117:10]
  assign _GEN_1189 = 6'h23 == _T_174 ? welem[35] : _GEN_1188; // @[Execute.scala 117:10]
  assign _GEN_1190 = 6'h24 == _T_174 ? welem[36] : _GEN_1189; // @[Execute.scala 117:10]
  assign _GEN_1191 = 6'h25 == _T_174 ? welem[37] : _GEN_1190; // @[Execute.scala 117:10]
  assign _GEN_1192 = 6'h26 == _T_174 ? welem[38] : _GEN_1191; // @[Execute.scala 117:10]
  assign _GEN_1193 = 6'h27 == _T_174 ? welem[39] : _GEN_1192; // @[Execute.scala 117:10]
  assign _GEN_1194 = 6'h28 == _T_174 ? welem[40] : _GEN_1193; // @[Execute.scala 117:10]
  assign _GEN_1195 = 6'h29 == _T_174 ? welem[41] : _GEN_1194; // @[Execute.scala 117:10]
  assign _GEN_1196 = 6'h2a == _T_174 ? welem[42] : _GEN_1195; // @[Execute.scala 117:10]
  assign _GEN_1197 = 6'h2b == _T_174 ? welem[43] : _GEN_1196; // @[Execute.scala 117:10]
  assign _GEN_1198 = 6'h2c == _T_174 ? welem[44] : _GEN_1197; // @[Execute.scala 117:10]
  assign _GEN_1199 = 6'h2d == _T_174 ? welem[45] : _GEN_1198; // @[Execute.scala 117:10]
  assign _GEN_1200 = 6'h2e == _T_174 ? welem[46] : _GEN_1199; // @[Execute.scala 117:10]
  assign _GEN_1201 = 6'h2f == _T_174 ? welem[47] : _GEN_1200; // @[Execute.scala 117:10]
  assign _GEN_1202 = 6'h30 == _T_174 ? welem[48] : _GEN_1201; // @[Execute.scala 117:10]
  assign _GEN_1203 = 6'h31 == _T_174 ? welem[49] : _GEN_1202; // @[Execute.scala 117:10]
  assign _GEN_1204 = 6'h32 == _T_174 ? welem[50] : _GEN_1203; // @[Execute.scala 117:10]
  assign _GEN_1205 = 6'h33 == _T_174 ? welem[51] : _GEN_1204; // @[Execute.scala 117:10]
  assign _GEN_1206 = 6'h34 == _T_174 ? welem[52] : _GEN_1205; // @[Execute.scala 117:10]
  assign _GEN_1207 = 6'h35 == _T_174 ? welem[53] : _GEN_1206; // @[Execute.scala 117:10]
  assign _GEN_1208 = 6'h36 == _T_174 ? welem[54] : _GEN_1207; // @[Execute.scala 117:10]
  assign _GEN_1209 = 6'h37 == _T_174 ? welem[55] : _GEN_1208; // @[Execute.scala 117:10]
  assign _GEN_1210 = 6'h38 == _T_174 ? welem[56] : _GEN_1209; // @[Execute.scala 117:10]
  assign _GEN_1211 = 6'h39 == _T_174 ? welem[57] : _GEN_1210; // @[Execute.scala 117:10]
  assign _GEN_1212 = 6'h3a == _T_174 ? welem[58] : _GEN_1211; // @[Execute.scala 117:10]
  assign _GEN_1213 = 6'h3b == _T_174 ? welem[59] : _GEN_1212; // @[Execute.scala 117:10]
  assign _GEN_1214 = 6'h3c == _T_174 ? welem[60] : _GEN_1213; // @[Execute.scala 117:10]
  assign _GEN_1215 = 6'h3d == _T_174 ? welem[61] : _GEN_1214; // @[Execute.scala 117:10]
  assign _GEN_1216 = 6'h3e == _T_174 ? welem[62] : _GEN_1215; // @[Execute.scala 117:10]
  assign _GEN_1217 = 6'h3f == _T_174 ? welem[63] : _GEN_1216; // @[Execute.scala 117:10]
  assign _GEN_1219 = 6'h1 == _T_178 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1220 = 6'h2 == _T_178 ? welem[2] : _GEN_1219; // @[Execute.scala 117:10]
  assign _GEN_1221 = 6'h3 == _T_178 ? welem[3] : _GEN_1220; // @[Execute.scala 117:10]
  assign _GEN_1222 = 6'h4 == _T_178 ? welem[4] : _GEN_1221; // @[Execute.scala 117:10]
  assign _GEN_1223 = 6'h5 == _T_178 ? welem[5] : _GEN_1222; // @[Execute.scala 117:10]
  assign _GEN_1224 = 6'h6 == _T_178 ? welem[6] : _GEN_1223; // @[Execute.scala 117:10]
  assign _GEN_1225 = 6'h7 == _T_178 ? welem[7] : _GEN_1224; // @[Execute.scala 117:10]
  assign _GEN_1226 = 6'h8 == _T_178 ? welem[8] : _GEN_1225; // @[Execute.scala 117:10]
  assign _GEN_1227 = 6'h9 == _T_178 ? welem[9] : _GEN_1226; // @[Execute.scala 117:10]
  assign _GEN_1228 = 6'ha == _T_178 ? welem[10] : _GEN_1227; // @[Execute.scala 117:10]
  assign _GEN_1229 = 6'hb == _T_178 ? welem[11] : _GEN_1228; // @[Execute.scala 117:10]
  assign _GEN_1230 = 6'hc == _T_178 ? welem[12] : _GEN_1229; // @[Execute.scala 117:10]
  assign _GEN_1231 = 6'hd == _T_178 ? welem[13] : _GEN_1230; // @[Execute.scala 117:10]
  assign _GEN_1232 = 6'he == _T_178 ? welem[14] : _GEN_1231; // @[Execute.scala 117:10]
  assign _GEN_1233 = 6'hf == _T_178 ? welem[15] : _GEN_1232; // @[Execute.scala 117:10]
  assign _GEN_1234 = 6'h10 == _T_178 ? welem[16] : _GEN_1233; // @[Execute.scala 117:10]
  assign _GEN_1235 = 6'h11 == _T_178 ? welem[17] : _GEN_1234; // @[Execute.scala 117:10]
  assign _GEN_1236 = 6'h12 == _T_178 ? welem[18] : _GEN_1235; // @[Execute.scala 117:10]
  assign _GEN_1237 = 6'h13 == _T_178 ? welem[19] : _GEN_1236; // @[Execute.scala 117:10]
  assign _GEN_1238 = 6'h14 == _T_178 ? welem[20] : _GEN_1237; // @[Execute.scala 117:10]
  assign _GEN_1239 = 6'h15 == _T_178 ? welem[21] : _GEN_1238; // @[Execute.scala 117:10]
  assign _GEN_1240 = 6'h16 == _T_178 ? welem[22] : _GEN_1239; // @[Execute.scala 117:10]
  assign _GEN_1241 = 6'h17 == _T_178 ? welem[23] : _GEN_1240; // @[Execute.scala 117:10]
  assign _GEN_1242 = 6'h18 == _T_178 ? welem[24] : _GEN_1241; // @[Execute.scala 117:10]
  assign _GEN_1243 = 6'h19 == _T_178 ? welem[25] : _GEN_1242; // @[Execute.scala 117:10]
  assign _GEN_1244 = 6'h1a == _T_178 ? welem[26] : _GEN_1243; // @[Execute.scala 117:10]
  assign _GEN_1245 = 6'h1b == _T_178 ? welem[27] : _GEN_1244; // @[Execute.scala 117:10]
  assign _GEN_1246 = 6'h1c == _T_178 ? welem[28] : _GEN_1245; // @[Execute.scala 117:10]
  assign _GEN_1247 = 6'h1d == _T_178 ? welem[29] : _GEN_1246; // @[Execute.scala 117:10]
  assign _GEN_1248 = 6'h1e == _T_178 ? welem[30] : _GEN_1247; // @[Execute.scala 117:10]
  assign _GEN_1249 = 6'h1f == _T_178 ? welem[31] : _GEN_1248; // @[Execute.scala 117:10]
  assign _GEN_1250 = 6'h20 == _T_178 ? welem[32] : _GEN_1249; // @[Execute.scala 117:10]
  assign _GEN_1251 = 6'h21 == _T_178 ? welem[33] : _GEN_1250; // @[Execute.scala 117:10]
  assign _GEN_1252 = 6'h22 == _T_178 ? welem[34] : _GEN_1251; // @[Execute.scala 117:10]
  assign _GEN_1253 = 6'h23 == _T_178 ? welem[35] : _GEN_1252; // @[Execute.scala 117:10]
  assign _GEN_1254 = 6'h24 == _T_178 ? welem[36] : _GEN_1253; // @[Execute.scala 117:10]
  assign _GEN_1255 = 6'h25 == _T_178 ? welem[37] : _GEN_1254; // @[Execute.scala 117:10]
  assign _GEN_1256 = 6'h26 == _T_178 ? welem[38] : _GEN_1255; // @[Execute.scala 117:10]
  assign _GEN_1257 = 6'h27 == _T_178 ? welem[39] : _GEN_1256; // @[Execute.scala 117:10]
  assign _GEN_1258 = 6'h28 == _T_178 ? welem[40] : _GEN_1257; // @[Execute.scala 117:10]
  assign _GEN_1259 = 6'h29 == _T_178 ? welem[41] : _GEN_1258; // @[Execute.scala 117:10]
  assign _GEN_1260 = 6'h2a == _T_178 ? welem[42] : _GEN_1259; // @[Execute.scala 117:10]
  assign _GEN_1261 = 6'h2b == _T_178 ? welem[43] : _GEN_1260; // @[Execute.scala 117:10]
  assign _GEN_1262 = 6'h2c == _T_178 ? welem[44] : _GEN_1261; // @[Execute.scala 117:10]
  assign _GEN_1263 = 6'h2d == _T_178 ? welem[45] : _GEN_1262; // @[Execute.scala 117:10]
  assign _GEN_1264 = 6'h2e == _T_178 ? welem[46] : _GEN_1263; // @[Execute.scala 117:10]
  assign _GEN_1265 = 6'h2f == _T_178 ? welem[47] : _GEN_1264; // @[Execute.scala 117:10]
  assign _GEN_1266 = 6'h30 == _T_178 ? welem[48] : _GEN_1265; // @[Execute.scala 117:10]
  assign _GEN_1267 = 6'h31 == _T_178 ? welem[49] : _GEN_1266; // @[Execute.scala 117:10]
  assign _GEN_1268 = 6'h32 == _T_178 ? welem[50] : _GEN_1267; // @[Execute.scala 117:10]
  assign _GEN_1269 = 6'h33 == _T_178 ? welem[51] : _GEN_1268; // @[Execute.scala 117:10]
  assign _GEN_1270 = 6'h34 == _T_178 ? welem[52] : _GEN_1269; // @[Execute.scala 117:10]
  assign _GEN_1271 = 6'h35 == _T_178 ? welem[53] : _GEN_1270; // @[Execute.scala 117:10]
  assign _GEN_1272 = 6'h36 == _T_178 ? welem[54] : _GEN_1271; // @[Execute.scala 117:10]
  assign _GEN_1273 = 6'h37 == _T_178 ? welem[55] : _GEN_1272; // @[Execute.scala 117:10]
  assign _GEN_1274 = 6'h38 == _T_178 ? welem[56] : _GEN_1273; // @[Execute.scala 117:10]
  assign _GEN_1275 = 6'h39 == _T_178 ? welem[57] : _GEN_1274; // @[Execute.scala 117:10]
  assign _GEN_1276 = 6'h3a == _T_178 ? welem[58] : _GEN_1275; // @[Execute.scala 117:10]
  assign _GEN_1277 = 6'h3b == _T_178 ? welem[59] : _GEN_1276; // @[Execute.scala 117:10]
  assign _GEN_1278 = 6'h3c == _T_178 ? welem[60] : _GEN_1277; // @[Execute.scala 117:10]
  assign _GEN_1279 = 6'h3d == _T_178 ? welem[61] : _GEN_1278; // @[Execute.scala 117:10]
  assign _GEN_1280 = 6'h3e == _T_178 ? welem[62] : _GEN_1279; // @[Execute.scala 117:10]
  assign _GEN_1281 = 6'h3f == _T_178 ? welem[63] : _GEN_1280; // @[Execute.scala 117:10]
  assign _T_181 = _T_172 ? _GEN_1217 : _GEN_1281; // @[Execute.scala 117:10]
  assign _T_182 = r < 6'h37; // @[Execute.scala 117:15]
  assign _T_184 = r - 6'h37; // @[Execute.scala 117:37]
  assign _T_188 = 6'h9 + r; // @[Execute.scala 117:60]
  assign _GEN_1283 = 6'h1 == _T_184 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1284 = 6'h2 == _T_184 ? welem[2] : _GEN_1283; // @[Execute.scala 117:10]
  assign _GEN_1285 = 6'h3 == _T_184 ? welem[3] : _GEN_1284; // @[Execute.scala 117:10]
  assign _GEN_1286 = 6'h4 == _T_184 ? welem[4] : _GEN_1285; // @[Execute.scala 117:10]
  assign _GEN_1287 = 6'h5 == _T_184 ? welem[5] : _GEN_1286; // @[Execute.scala 117:10]
  assign _GEN_1288 = 6'h6 == _T_184 ? welem[6] : _GEN_1287; // @[Execute.scala 117:10]
  assign _GEN_1289 = 6'h7 == _T_184 ? welem[7] : _GEN_1288; // @[Execute.scala 117:10]
  assign _GEN_1290 = 6'h8 == _T_184 ? welem[8] : _GEN_1289; // @[Execute.scala 117:10]
  assign _GEN_1291 = 6'h9 == _T_184 ? welem[9] : _GEN_1290; // @[Execute.scala 117:10]
  assign _GEN_1292 = 6'ha == _T_184 ? welem[10] : _GEN_1291; // @[Execute.scala 117:10]
  assign _GEN_1293 = 6'hb == _T_184 ? welem[11] : _GEN_1292; // @[Execute.scala 117:10]
  assign _GEN_1294 = 6'hc == _T_184 ? welem[12] : _GEN_1293; // @[Execute.scala 117:10]
  assign _GEN_1295 = 6'hd == _T_184 ? welem[13] : _GEN_1294; // @[Execute.scala 117:10]
  assign _GEN_1296 = 6'he == _T_184 ? welem[14] : _GEN_1295; // @[Execute.scala 117:10]
  assign _GEN_1297 = 6'hf == _T_184 ? welem[15] : _GEN_1296; // @[Execute.scala 117:10]
  assign _GEN_1298 = 6'h10 == _T_184 ? welem[16] : _GEN_1297; // @[Execute.scala 117:10]
  assign _GEN_1299 = 6'h11 == _T_184 ? welem[17] : _GEN_1298; // @[Execute.scala 117:10]
  assign _GEN_1300 = 6'h12 == _T_184 ? welem[18] : _GEN_1299; // @[Execute.scala 117:10]
  assign _GEN_1301 = 6'h13 == _T_184 ? welem[19] : _GEN_1300; // @[Execute.scala 117:10]
  assign _GEN_1302 = 6'h14 == _T_184 ? welem[20] : _GEN_1301; // @[Execute.scala 117:10]
  assign _GEN_1303 = 6'h15 == _T_184 ? welem[21] : _GEN_1302; // @[Execute.scala 117:10]
  assign _GEN_1304 = 6'h16 == _T_184 ? welem[22] : _GEN_1303; // @[Execute.scala 117:10]
  assign _GEN_1305 = 6'h17 == _T_184 ? welem[23] : _GEN_1304; // @[Execute.scala 117:10]
  assign _GEN_1306 = 6'h18 == _T_184 ? welem[24] : _GEN_1305; // @[Execute.scala 117:10]
  assign _GEN_1307 = 6'h19 == _T_184 ? welem[25] : _GEN_1306; // @[Execute.scala 117:10]
  assign _GEN_1308 = 6'h1a == _T_184 ? welem[26] : _GEN_1307; // @[Execute.scala 117:10]
  assign _GEN_1309 = 6'h1b == _T_184 ? welem[27] : _GEN_1308; // @[Execute.scala 117:10]
  assign _GEN_1310 = 6'h1c == _T_184 ? welem[28] : _GEN_1309; // @[Execute.scala 117:10]
  assign _GEN_1311 = 6'h1d == _T_184 ? welem[29] : _GEN_1310; // @[Execute.scala 117:10]
  assign _GEN_1312 = 6'h1e == _T_184 ? welem[30] : _GEN_1311; // @[Execute.scala 117:10]
  assign _GEN_1313 = 6'h1f == _T_184 ? welem[31] : _GEN_1312; // @[Execute.scala 117:10]
  assign _GEN_1314 = 6'h20 == _T_184 ? welem[32] : _GEN_1313; // @[Execute.scala 117:10]
  assign _GEN_1315 = 6'h21 == _T_184 ? welem[33] : _GEN_1314; // @[Execute.scala 117:10]
  assign _GEN_1316 = 6'h22 == _T_184 ? welem[34] : _GEN_1315; // @[Execute.scala 117:10]
  assign _GEN_1317 = 6'h23 == _T_184 ? welem[35] : _GEN_1316; // @[Execute.scala 117:10]
  assign _GEN_1318 = 6'h24 == _T_184 ? welem[36] : _GEN_1317; // @[Execute.scala 117:10]
  assign _GEN_1319 = 6'h25 == _T_184 ? welem[37] : _GEN_1318; // @[Execute.scala 117:10]
  assign _GEN_1320 = 6'h26 == _T_184 ? welem[38] : _GEN_1319; // @[Execute.scala 117:10]
  assign _GEN_1321 = 6'h27 == _T_184 ? welem[39] : _GEN_1320; // @[Execute.scala 117:10]
  assign _GEN_1322 = 6'h28 == _T_184 ? welem[40] : _GEN_1321; // @[Execute.scala 117:10]
  assign _GEN_1323 = 6'h29 == _T_184 ? welem[41] : _GEN_1322; // @[Execute.scala 117:10]
  assign _GEN_1324 = 6'h2a == _T_184 ? welem[42] : _GEN_1323; // @[Execute.scala 117:10]
  assign _GEN_1325 = 6'h2b == _T_184 ? welem[43] : _GEN_1324; // @[Execute.scala 117:10]
  assign _GEN_1326 = 6'h2c == _T_184 ? welem[44] : _GEN_1325; // @[Execute.scala 117:10]
  assign _GEN_1327 = 6'h2d == _T_184 ? welem[45] : _GEN_1326; // @[Execute.scala 117:10]
  assign _GEN_1328 = 6'h2e == _T_184 ? welem[46] : _GEN_1327; // @[Execute.scala 117:10]
  assign _GEN_1329 = 6'h2f == _T_184 ? welem[47] : _GEN_1328; // @[Execute.scala 117:10]
  assign _GEN_1330 = 6'h30 == _T_184 ? welem[48] : _GEN_1329; // @[Execute.scala 117:10]
  assign _GEN_1331 = 6'h31 == _T_184 ? welem[49] : _GEN_1330; // @[Execute.scala 117:10]
  assign _GEN_1332 = 6'h32 == _T_184 ? welem[50] : _GEN_1331; // @[Execute.scala 117:10]
  assign _GEN_1333 = 6'h33 == _T_184 ? welem[51] : _GEN_1332; // @[Execute.scala 117:10]
  assign _GEN_1334 = 6'h34 == _T_184 ? welem[52] : _GEN_1333; // @[Execute.scala 117:10]
  assign _GEN_1335 = 6'h35 == _T_184 ? welem[53] : _GEN_1334; // @[Execute.scala 117:10]
  assign _GEN_1336 = 6'h36 == _T_184 ? welem[54] : _GEN_1335; // @[Execute.scala 117:10]
  assign _GEN_1337 = 6'h37 == _T_184 ? welem[55] : _GEN_1336; // @[Execute.scala 117:10]
  assign _GEN_1338 = 6'h38 == _T_184 ? welem[56] : _GEN_1337; // @[Execute.scala 117:10]
  assign _GEN_1339 = 6'h39 == _T_184 ? welem[57] : _GEN_1338; // @[Execute.scala 117:10]
  assign _GEN_1340 = 6'h3a == _T_184 ? welem[58] : _GEN_1339; // @[Execute.scala 117:10]
  assign _GEN_1341 = 6'h3b == _T_184 ? welem[59] : _GEN_1340; // @[Execute.scala 117:10]
  assign _GEN_1342 = 6'h3c == _T_184 ? welem[60] : _GEN_1341; // @[Execute.scala 117:10]
  assign _GEN_1343 = 6'h3d == _T_184 ? welem[61] : _GEN_1342; // @[Execute.scala 117:10]
  assign _GEN_1344 = 6'h3e == _T_184 ? welem[62] : _GEN_1343; // @[Execute.scala 117:10]
  assign _GEN_1345 = 6'h3f == _T_184 ? welem[63] : _GEN_1344; // @[Execute.scala 117:10]
  assign _GEN_1347 = 6'h1 == _T_188 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1348 = 6'h2 == _T_188 ? welem[2] : _GEN_1347; // @[Execute.scala 117:10]
  assign _GEN_1349 = 6'h3 == _T_188 ? welem[3] : _GEN_1348; // @[Execute.scala 117:10]
  assign _GEN_1350 = 6'h4 == _T_188 ? welem[4] : _GEN_1349; // @[Execute.scala 117:10]
  assign _GEN_1351 = 6'h5 == _T_188 ? welem[5] : _GEN_1350; // @[Execute.scala 117:10]
  assign _GEN_1352 = 6'h6 == _T_188 ? welem[6] : _GEN_1351; // @[Execute.scala 117:10]
  assign _GEN_1353 = 6'h7 == _T_188 ? welem[7] : _GEN_1352; // @[Execute.scala 117:10]
  assign _GEN_1354 = 6'h8 == _T_188 ? welem[8] : _GEN_1353; // @[Execute.scala 117:10]
  assign _GEN_1355 = 6'h9 == _T_188 ? welem[9] : _GEN_1354; // @[Execute.scala 117:10]
  assign _GEN_1356 = 6'ha == _T_188 ? welem[10] : _GEN_1355; // @[Execute.scala 117:10]
  assign _GEN_1357 = 6'hb == _T_188 ? welem[11] : _GEN_1356; // @[Execute.scala 117:10]
  assign _GEN_1358 = 6'hc == _T_188 ? welem[12] : _GEN_1357; // @[Execute.scala 117:10]
  assign _GEN_1359 = 6'hd == _T_188 ? welem[13] : _GEN_1358; // @[Execute.scala 117:10]
  assign _GEN_1360 = 6'he == _T_188 ? welem[14] : _GEN_1359; // @[Execute.scala 117:10]
  assign _GEN_1361 = 6'hf == _T_188 ? welem[15] : _GEN_1360; // @[Execute.scala 117:10]
  assign _GEN_1362 = 6'h10 == _T_188 ? welem[16] : _GEN_1361; // @[Execute.scala 117:10]
  assign _GEN_1363 = 6'h11 == _T_188 ? welem[17] : _GEN_1362; // @[Execute.scala 117:10]
  assign _GEN_1364 = 6'h12 == _T_188 ? welem[18] : _GEN_1363; // @[Execute.scala 117:10]
  assign _GEN_1365 = 6'h13 == _T_188 ? welem[19] : _GEN_1364; // @[Execute.scala 117:10]
  assign _GEN_1366 = 6'h14 == _T_188 ? welem[20] : _GEN_1365; // @[Execute.scala 117:10]
  assign _GEN_1367 = 6'h15 == _T_188 ? welem[21] : _GEN_1366; // @[Execute.scala 117:10]
  assign _GEN_1368 = 6'h16 == _T_188 ? welem[22] : _GEN_1367; // @[Execute.scala 117:10]
  assign _GEN_1369 = 6'h17 == _T_188 ? welem[23] : _GEN_1368; // @[Execute.scala 117:10]
  assign _GEN_1370 = 6'h18 == _T_188 ? welem[24] : _GEN_1369; // @[Execute.scala 117:10]
  assign _GEN_1371 = 6'h19 == _T_188 ? welem[25] : _GEN_1370; // @[Execute.scala 117:10]
  assign _GEN_1372 = 6'h1a == _T_188 ? welem[26] : _GEN_1371; // @[Execute.scala 117:10]
  assign _GEN_1373 = 6'h1b == _T_188 ? welem[27] : _GEN_1372; // @[Execute.scala 117:10]
  assign _GEN_1374 = 6'h1c == _T_188 ? welem[28] : _GEN_1373; // @[Execute.scala 117:10]
  assign _GEN_1375 = 6'h1d == _T_188 ? welem[29] : _GEN_1374; // @[Execute.scala 117:10]
  assign _GEN_1376 = 6'h1e == _T_188 ? welem[30] : _GEN_1375; // @[Execute.scala 117:10]
  assign _GEN_1377 = 6'h1f == _T_188 ? welem[31] : _GEN_1376; // @[Execute.scala 117:10]
  assign _GEN_1378 = 6'h20 == _T_188 ? welem[32] : _GEN_1377; // @[Execute.scala 117:10]
  assign _GEN_1379 = 6'h21 == _T_188 ? welem[33] : _GEN_1378; // @[Execute.scala 117:10]
  assign _GEN_1380 = 6'h22 == _T_188 ? welem[34] : _GEN_1379; // @[Execute.scala 117:10]
  assign _GEN_1381 = 6'h23 == _T_188 ? welem[35] : _GEN_1380; // @[Execute.scala 117:10]
  assign _GEN_1382 = 6'h24 == _T_188 ? welem[36] : _GEN_1381; // @[Execute.scala 117:10]
  assign _GEN_1383 = 6'h25 == _T_188 ? welem[37] : _GEN_1382; // @[Execute.scala 117:10]
  assign _GEN_1384 = 6'h26 == _T_188 ? welem[38] : _GEN_1383; // @[Execute.scala 117:10]
  assign _GEN_1385 = 6'h27 == _T_188 ? welem[39] : _GEN_1384; // @[Execute.scala 117:10]
  assign _GEN_1386 = 6'h28 == _T_188 ? welem[40] : _GEN_1385; // @[Execute.scala 117:10]
  assign _GEN_1387 = 6'h29 == _T_188 ? welem[41] : _GEN_1386; // @[Execute.scala 117:10]
  assign _GEN_1388 = 6'h2a == _T_188 ? welem[42] : _GEN_1387; // @[Execute.scala 117:10]
  assign _GEN_1389 = 6'h2b == _T_188 ? welem[43] : _GEN_1388; // @[Execute.scala 117:10]
  assign _GEN_1390 = 6'h2c == _T_188 ? welem[44] : _GEN_1389; // @[Execute.scala 117:10]
  assign _GEN_1391 = 6'h2d == _T_188 ? welem[45] : _GEN_1390; // @[Execute.scala 117:10]
  assign _GEN_1392 = 6'h2e == _T_188 ? welem[46] : _GEN_1391; // @[Execute.scala 117:10]
  assign _GEN_1393 = 6'h2f == _T_188 ? welem[47] : _GEN_1392; // @[Execute.scala 117:10]
  assign _GEN_1394 = 6'h30 == _T_188 ? welem[48] : _GEN_1393; // @[Execute.scala 117:10]
  assign _GEN_1395 = 6'h31 == _T_188 ? welem[49] : _GEN_1394; // @[Execute.scala 117:10]
  assign _GEN_1396 = 6'h32 == _T_188 ? welem[50] : _GEN_1395; // @[Execute.scala 117:10]
  assign _GEN_1397 = 6'h33 == _T_188 ? welem[51] : _GEN_1396; // @[Execute.scala 117:10]
  assign _GEN_1398 = 6'h34 == _T_188 ? welem[52] : _GEN_1397; // @[Execute.scala 117:10]
  assign _GEN_1399 = 6'h35 == _T_188 ? welem[53] : _GEN_1398; // @[Execute.scala 117:10]
  assign _GEN_1400 = 6'h36 == _T_188 ? welem[54] : _GEN_1399; // @[Execute.scala 117:10]
  assign _GEN_1401 = 6'h37 == _T_188 ? welem[55] : _GEN_1400; // @[Execute.scala 117:10]
  assign _GEN_1402 = 6'h38 == _T_188 ? welem[56] : _GEN_1401; // @[Execute.scala 117:10]
  assign _GEN_1403 = 6'h39 == _T_188 ? welem[57] : _GEN_1402; // @[Execute.scala 117:10]
  assign _GEN_1404 = 6'h3a == _T_188 ? welem[58] : _GEN_1403; // @[Execute.scala 117:10]
  assign _GEN_1405 = 6'h3b == _T_188 ? welem[59] : _GEN_1404; // @[Execute.scala 117:10]
  assign _GEN_1406 = 6'h3c == _T_188 ? welem[60] : _GEN_1405; // @[Execute.scala 117:10]
  assign _GEN_1407 = 6'h3d == _T_188 ? welem[61] : _GEN_1406; // @[Execute.scala 117:10]
  assign _GEN_1408 = 6'h3e == _T_188 ? welem[62] : _GEN_1407; // @[Execute.scala 117:10]
  assign _GEN_1409 = 6'h3f == _T_188 ? welem[63] : _GEN_1408; // @[Execute.scala 117:10]
  assign _T_191 = _T_182 ? _GEN_1345 : _GEN_1409; // @[Execute.scala 117:10]
  assign _T_192 = r < 6'h36; // @[Execute.scala 117:15]
  assign _T_194 = r - 6'h36; // @[Execute.scala 117:37]
  assign _T_198 = 6'ha + r; // @[Execute.scala 117:60]
  assign _GEN_1411 = 6'h1 == _T_194 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1412 = 6'h2 == _T_194 ? welem[2] : _GEN_1411; // @[Execute.scala 117:10]
  assign _GEN_1413 = 6'h3 == _T_194 ? welem[3] : _GEN_1412; // @[Execute.scala 117:10]
  assign _GEN_1414 = 6'h4 == _T_194 ? welem[4] : _GEN_1413; // @[Execute.scala 117:10]
  assign _GEN_1415 = 6'h5 == _T_194 ? welem[5] : _GEN_1414; // @[Execute.scala 117:10]
  assign _GEN_1416 = 6'h6 == _T_194 ? welem[6] : _GEN_1415; // @[Execute.scala 117:10]
  assign _GEN_1417 = 6'h7 == _T_194 ? welem[7] : _GEN_1416; // @[Execute.scala 117:10]
  assign _GEN_1418 = 6'h8 == _T_194 ? welem[8] : _GEN_1417; // @[Execute.scala 117:10]
  assign _GEN_1419 = 6'h9 == _T_194 ? welem[9] : _GEN_1418; // @[Execute.scala 117:10]
  assign _GEN_1420 = 6'ha == _T_194 ? welem[10] : _GEN_1419; // @[Execute.scala 117:10]
  assign _GEN_1421 = 6'hb == _T_194 ? welem[11] : _GEN_1420; // @[Execute.scala 117:10]
  assign _GEN_1422 = 6'hc == _T_194 ? welem[12] : _GEN_1421; // @[Execute.scala 117:10]
  assign _GEN_1423 = 6'hd == _T_194 ? welem[13] : _GEN_1422; // @[Execute.scala 117:10]
  assign _GEN_1424 = 6'he == _T_194 ? welem[14] : _GEN_1423; // @[Execute.scala 117:10]
  assign _GEN_1425 = 6'hf == _T_194 ? welem[15] : _GEN_1424; // @[Execute.scala 117:10]
  assign _GEN_1426 = 6'h10 == _T_194 ? welem[16] : _GEN_1425; // @[Execute.scala 117:10]
  assign _GEN_1427 = 6'h11 == _T_194 ? welem[17] : _GEN_1426; // @[Execute.scala 117:10]
  assign _GEN_1428 = 6'h12 == _T_194 ? welem[18] : _GEN_1427; // @[Execute.scala 117:10]
  assign _GEN_1429 = 6'h13 == _T_194 ? welem[19] : _GEN_1428; // @[Execute.scala 117:10]
  assign _GEN_1430 = 6'h14 == _T_194 ? welem[20] : _GEN_1429; // @[Execute.scala 117:10]
  assign _GEN_1431 = 6'h15 == _T_194 ? welem[21] : _GEN_1430; // @[Execute.scala 117:10]
  assign _GEN_1432 = 6'h16 == _T_194 ? welem[22] : _GEN_1431; // @[Execute.scala 117:10]
  assign _GEN_1433 = 6'h17 == _T_194 ? welem[23] : _GEN_1432; // @[Execute.scala 117:10]
  assign _GEN_1434 = 6'h18 == _T_194 ? welem[24] : _GEN_1433; // @[Execute.scala 117:10]
  assign _GEN_1435 = 6'h19 == _T_194 ? welem[25] : _GEN_1434; // @[Execute.scala 117:10]
  assign _GEN_1436 = 6'h1a == _T_194 ? welem[26] : _GEN_1435; // @[Execute.scala 117:10]
  assign _GEN_1437 = 6'h1b == _T_194 ? welem[27] : _GEN_1436; // @[Execute.scala 117:10]
  assign _GEN_1438 = 6'h1c == _T_194 ? welem[28] : _GEN_1437; // @[Execute.scala 117:10]
  assign _GEN_1439 = 6'h1d == _T_194 ? welem[29] : _GEN_1438; // @[Execute.scala 117:10]
  assign _GEN_1440 = 6'h1e == _T_194 ? welem[30] : _GEN_1439; // @[Execute.scala 117:10]
  assign _GEN_1441 = 6'h1f == _T_194 ? welem[31] : _GEN_1440; // @[Execute.scala 117:10]
  assign _GEN_1442 = 6'h20 == _T_194 ? welem[32] : _GEN_1441; // @[Execute.scala 117:10]
  assign _GEN_1443 = 6'h21 == _T_194 ? welem[33] : _GEN_1442; // @[Execute.scala 117:10]
  assign _GEN_1444 = 6'h22 == _T_194 ? welem[34] : _GEN_1443; // @[Execute.scala 117:10]
  assign _GEN_1445 = 6'h23 == _T_194 ? welem[35] : _GEN_1444; // @[Execute.scala 117:10]
  assign _GEN_1446 = 6'h24 == _T_194 ? welem[36] : _GEN_1445; // @[Execute.scala 117:10]
  assign _GEN_1447 = 6'h25 == _T_194 ? welem[37] : _GEN_1446; // @[Execute.scala 117:10]
  assign _GEN_1448 = 6'h26 == _T_194 ? welem[38] : _GEN_1447; // @[Execute.scala 117:10]
  assign _GEN_1449 = 6'h27 == _T_194 ? welem[39] : _GEN_1448; // @[Execute.scala 117:10]
  assign _GEN_1450 = 6'h28 == _T_194 ? welem[40] : _GEN_1449; // @[Execute.scala 117:10]
  assign _GEN_1451 = 6'h29 == _T_194 ? welem[41] : _GEN_1450; // @[Execute.scala 117:10]
  assign _GEN_1452 = 6'h2a == _T_194 ? welem[42] : _GEN_1451; // @[Execute.scala 117:10]
  assign _GEN_1453 = 6'h2b == _T_194 ? welem[43] : _GEN_1452; // @[Execute.scala 117:10]
  assign _GEN_1454 = 6'h2c == _T_194 ? welem[44] : _GEN_1453; // @[Execute.scala 117:10]
  assign _GEN_1455 = 6'h2d == _T_194 ? welem[45] : _GEN_1454; // @[Execute.scala 117:10]
  assign _GEN_1456 = 6'h2e == _T_194 ? welem[46] : _GEN_1455; // @[Execute.scala 117:10]
  assign _GEN_1457 = 6'h2f == _T_194 ? welem[47] : _GEN_1456; // @[Execute.scala 117:10]
  assign _GEN_1458 = 6'h30 == _T_194 ? welem[48] : _GEN_1457; // @[Execute.scala 117:10]
  assign _GEN_1459 = 6'h31 == _T_194 ? welem[49] : _GEN_1458; // @[Execute.scala 117:10]
  assign _GEN_1460 = 6'h32 == _T_194 ? welem[50] : _GEN_1459; // @[Execute.scala 117:10]
  assign _GEN_1461 = 6'h33 == _T_194 ? welem[51] : _GEN_1460; // @[Execute.scala 117:10]
  assign _GEN_1462 = 6'h34 == _T_194 ? welem[52] : _GEN_1461; // @[Execute.scala 117:10]
  assign _GEN_1463 = 6'h35 == _T_194 ? welem[53] : _GEN_1462; // @[Execute.scala 117:10]
  assign _GEN_1464 = 6'h36 == _T_194 ? welem[54] : _GEN_1463; // @[Execute.scala 117:10]
  assign _GEN_1465 = 6'h37 == _T_194 ? welem[55] : _GEN_1464; // @[Execute.scala 117:10]
  assign _GEN_1466 = 6'h38 == _T_194 ? welem[56] : _GEN_1465; // @[Execute.scala 117:10]
  assign _GEN_1467 = 6'h39 == _T_194 ? welem[57] : _GEN_1466; // @[Execute.scala 117:10]
  assign _GEN_1468 = 6'h3a == _T_194 ? welem[58] : _GEN_1467; // @[Execute.scala 117:10]
  assign _GEN_1469 = 6'h3b == _T_194 ? welem[59] : _GEN_1468; // @[Execute.scala 117:10]
  assign _GEN_1470 = 6'h3c == _T_194 ? welem[60] : _GEN_1469; // @[Execute.scala 117:10]
  assign _GEN_1471 = 6'h3d == _T_194 ? welem[61] : _GEN_1470; // @[Execute.scala 117:10]
  assign _GEN_1472 = 6'h3e == _T_194 ? welem[62] : _GEN_1471; // @[Execute.scala 117:10]
  assign _GEN_1473 = 6'h3f == _T_194 ? welem[63] : _GEN_1472; // @[Execute.scala 117:10]
  assign _GEN_1475 = 6'h1 == _T_198 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1476 = 6'h2 == _T_198 ? welem[2] : _GEN_1475; // @[Execute.scala 117:10]
  assign _GEN_1477 = 6'h3 == _T_198 ? welem[3] : _GEN_1476; // @[Execute.scala 117:10]
  assign _GEN_1478 = 6'h4 == _T_198 ? welem[4] : _GEN_1477; // @[Execute.scala 117:10]
  assign _GEN_1479 = 6'h5 == _T_198 ? welem[5] : _GEN_1478; // @[Execute.scala 117:10]
  assign _GEN_1480 = 6'h6 == _T_198 ? welem[6] : _GEN_1479; // @[Execute.scala 117:10]
  assign _GEN_1481 = 6'h7 == _T_198 ? welem[7] : _GEN_1480; // @[Execute.scala 117:10]
  assign _GEN_1482 = 6'h8 == _T_198 ? welem[8] : _GEN_1481; // @[Execute.scala 117:10]
  assign _GEN_1483 = 6'h9 == _T_198 ? welem[9] : _GEN_1482; // @[Execute.scala 117:10]
  assign _GEN_1484 = 6'ha == _T_198 ? welem[10] : _GEN_1483; // @[Execute.scala 117:10]
  assign _GEN_1485 = 6'hb == _T_198 ? welem[11] : _GEN_1484; // @[Execute.scala 117:10]
  assign _GEN_1486 = 6'hc == _T_198 ? welem[12] : _GEN_1485; // @[Execute.scala 117:10]
  assign _GEN_1487 = 6'hd == _T_198 ? welem[13] : _GEN_1486; // @[Execute.scala 117:10]
  assign _GEN_1488 = 6'he == _T_198 ? welem[14] : _GEN_1487; // @[Execute.scala 117:10]
  assign _GEN_1489 = 6'hf == _T_198 ? welem[15] : _GEN_1488; // @[Execute.scala 117:10]
  assign _GEN_1490 = 6'h10 == _T_198 ? welem[16] : _GEN_1489; // @[Execute.scala 117:10]
  assign _GEN_1491 = 6'h11 == _T_198 ? welem[17] : _GEN_1490; // @[Execute.scala 117:10]
  assign _GEN_1492 = 6'h12 == _T_198 ? welem[18] : _GEN_1491; // @[Execute.scala 117:10]
  assign _GEN_1493 = 6'h13 == _T_198 ? welem[19] : _GEN_1492; // @[Execute.scala 117:10]
  assign _GEN_1494 = 6'h14 == _T_198 ? welem[20] : _GEN_1493; // @[Execute.scala 117:10]
  assign _GEN_1495 = 6'h15 == _T_198 ? welem[21] : _GEN_1494; // @[Execute.scala 117:10]
  assign _GEN_1496 = 6'h16 == _T_198 ? welem[22] : _GEN_1495; // @[Execute.scala 117:10]
  assign _GEN_1497 = 6'h17 == _T_198 ? welem[23] : _GEN_1496; // @[Execute.scala 117:10]
  assign _GEN_1498 = 6'h18 == _T_198 ? welem[24] : _GEN_1497; // @[Execute.scala 117:10]
  assign _GEN_1499 = 6'h19 == _T_198 ? welem[25] : _GEN_1498; // @[Execute.scala 117:10]
  assign _GEN_1500 = 6'h1a == _T_198 ? welem[26] : _GEN_1499; // @[Execute.scala 117:10]
  assign _GEN_1501 = 6'h1b == _T_198 ? welem[27] : _GEN_1500; // @[Execute.scala 117:10]
  assign _GEN_1502 = 6'h1c == _T_198 ? welem[28] : _GEN_1501; // @[Execute.scala 117:10]
  assign _GEN_1503 = 6'h1d == _T_198 ? welem[29] : _GEN_1502; // @[Execute.scala 117:10]
  assign _GEN_1504 = 6'h1e == _T_198 ? welem[30] : _GEN_1503; // @[Execute.scala 117:10]
  assign _GEN_1505 = 6'h1f == _T_198 ? welem[31] : _GEN_1504; // @[Execute.scala 117:10]
  assign _GEN_1506 = 6'h20 == _T_198 ? welem[32] : _GEN_1505; // @[Execute.scala 117:10]
  assign _GEN_1507 = 6'h21 == _T_198 ? welem[33] : _GEN_1506; // @[Execute.scala 117:10]
  assign _GEN_1508 = 6'h22 == _T_198 ? welem[34] : _GEN_1507; // @[Execute.scala 117:10]
  assign _GEN_1509 = 6'h23 == _T_198 ? welem[35] : _GEN_1508; // @[Execute.scala 117:10]
  assign _GEN_1510 = 6'h24 == _T_198 ? welem[36] : _GEN_1509; // @[Execute.scala 117:10]
  assign _GEN_1511 = 6'h25 == _T_198 ? welem[37] : _GEN_1510; // @[Execute.scala 117:10]
  assign _GEN_1512 = 6'h26 == _T_198 ? welem[38] : _GEN_1511; // @[Execute.scala 117:10]
  assign _GEN_1513 = 6'h27 == _T_198 ? welem[39] : _GEN_1512; // @[Execute.scala 117:10]
  assign _GEN_1514 = 6'h28 == _T_198 ? welem[40] : _GEN_1513; // @[Execute.scala 117:10]
  assign _GEN_1515 = 6'h29 == _T_198 ? welem[41] : _GEN_1514; // @[Execute.scala 117:10]
  assign _GEN_1516 = 6'h2a == _T_198 ? welem[42] : _GEN_1515; // @[Execute.scala 117:10]
  assign _GEN_1517 = 6'h2b == _T_198 ? welem[43] : _GEN_1516; // @[Execute.scala 117:10]
  assign _GEN_1518 = 6'h2c == _T_198 ? welem[44] : _GEN_1517; // @[Execute.scala 117:10]
  assign _GEN_1519 = 6'h2d == _T_198 ? welem[45] : _GEN_1518; // @[Execute.scala 117:10]
  assign _GEN_1520 = 6'h2e == _T_198 ? welem[46] : _GEN_1519; // @[Execute.scala 117:10]
  assign _GEN_1521 = 6'h2f == _T_198 ? welem[47] : _GEN_1520; // @[Execute.scala 117:10]
  assign _GEN_1522 = 6'h30 == _T_198 ? welem[48] : _GEN_1521; // @[Execute.scala 117:10]
  assign _GEN_1523 = 6'h31 == _T_198 ? welem[49] : _GEN_1522; // @[Execute.scala 117:10]
  assign _GEN_1524 = 6'h32 == _T_198 ? welem[50] : _GEN_1523; // @[Execute.scala 117:10]
  assign _GEN_1525 = 6'h33 == _T_198 ? welem[51] : _GEN_1524; // @[Execute.scala 117:10]
  assign _GEN_1526 = 6'h34 == _T_198 ? welem[52] : _GEN_1525; // @[Execute.scala 117:10]
  assign _GEN_1527 = 6'h35 == _T_198 ? welem[53] : _GEN_1526; // @[Execute.scala 117:10]
  assign _GEN_1528 = 6'h36 == _T_198 ? welem[54] : _GEN_1527; // @[Execute.scala 117:10]
  assign _GEN_1529 = 6'h37 == _T_198 ? welem[55] : _GEN_1528; // @[Execute.scala 117:10]
  assign _GEN_1530 = 6'h38 == _T_198 ? welem[56] : _GEN_1529; // @[Execute.scala 117:10]
  assign _GEN_1531 = 6'h39 == _T_198 ? welem[57] : _GEN_1530; // @[Execute.scala 117:10]
  assign _GEN_1532 = 6'h3a == _T_198 ? welem[58] : _GEN_1531; // @[Execute.scala 117:10]
  assign _GEN_1533 = 6'h3b == _T_198 ? welem[59] : _GEN_1532; // @[Execute.scala 117:10]
  assign _GEN_1534 = 6'h3c == _T_198 ? welem[60] : _GEN_1533; // @[Execute.scala 117:10]
  assign _GEN_1535 = 6'h3d == _T_198 ? welem[61] : _GEN_1534; // @[Execute.scala 117:10]
  assign _GEN_1536 = 6'h3e == _T_198 ? welem[62] : _GEN_1535; // @[Execute.scala 117:10]
  assign _GEN_1537 = 6'h3f == _T_198 ? welem[63] : _GEN_1536; // @[Execute.scala 117:10]
  assign _T_201 = _T_192 ? _GEN_1473 : _GEN_1537; // @[Execute.scala 117:10]
  assign _T_202 = r < 6'h35; // @[Execute.scala 117:15]
  assign _T_204 = r - 6'h35; // @[Execute.scala 117:37]
  assign _T_208 = 6'hb + r; // @[Execute.scala 117:60]
  assign _GEN_1539 = 6'h1 == _T_204 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1540 = 6'h2 == _T_204 ? welem[2] : _GEN_1539; // @[Execute.scala 117:10]
  assign _GEN_1541 = 6'h3 == _T_204 ? welem[3] : _GEN_1540; // @[Execute.scala 117:10]
  assign _GEN_1542 = 6'h4 == _T_204 ? welem[4] : _GEN_1541; // @[Execute.scala 117:10]
  assign _GEN_1543 = 6'h5 == _T_204 ? welem[5] : _GEN_1542; // @[Execute.scala 117:10]
  assign _GEN_1544 = 6'h6 == _T_204 ? welem[6] : _GEN_1543; // @[Execute.scala 117:10]
  assign _GEN_1545 = 6'h7 == _T_204 ? welem[7] : _GEN_1544; // @[Execute.scala 117:10]
  assign _GEN_1546 = 6'h8 == _T_204 ? welem[8] : _GEN_1545; // @[Execute.scala 117:10]
  assign _GEN_1547 = 6'h9 == _T_204 ? welem[9] : _GEN_1546; // @[Execute.scala 117:10]
  assign _GEN_1548 = 6'ha == _T_204 ? welem[10] : _GEN_1547; // @[Execute.scala 117:10]
  assign _GEN_1549 = 6'hb == _T_204 ? welem[11] : _GEN_1548; // @[Execute.scala 117:10]
  assign _GEN_1550 = 6'hc == _T_204 ? welem[12] : _GEN_1549; // @[Execute.scala 117:10]
  assign _GEN_1551 = 6'hd == _T_204 ? welem[13] : _GEN_1550; // @[Execute.scala 117:10]
  assign _GEN_1552 = 6'he == _T_204 ? welem[14] : _GEN_1551; // @[Execute.scala 117:10]
  assign _GEN_1553 = 6'hf == _T_204 ? welem[15] : _GEN_1552; // @[Execute.scala 117:10]
  assign _GEN_1554 = 6'h10 == _T_204 ? welem[16] : _GEN_1553; // @[Execute.scala 117:10]
  assign _GEN_1555 = 6'h11 == _T_204 ? welem[17] : _GEN_1554; // @[Execute.scala 117:10]
  assign _GEN_1556 = 6'h12 == _T_204 ? welem[18] : _GEN_1555; // @[Execute.scala 117:10]
  assign _GEN_1557 = 6'h13 == _T_204 ? welem[19] : _GEN_1556; // @[Execute.scala 117:10]
  assign _GEN_1558 = 6'h14 == _T_204 ? welem[20] : _GEN_1557; // @[Execute.scala 117:10]
  assign _GEN_1559 = 6'h15 == _T_204 ? welem[21] : _GEN_1558; // @[Execute.scala 117:10]
  assign _GEN_1560 = 6'h16 == _T_204 ? welem[22] : _GEN_1559; // @[Execute.scala 117:10]
  assign _GEN_1561 = 6'h17 == _T_204 ? welem[23] : _GEN_1560; // @[Execute.scala 117:10]
  assign _GEN_1562 = 6'h18 == _T_204 ? welem[24] : _GEN_1561; // @[Execute.scala 117:10]
  assign _GEN_1563 = 6'h19 == _T_204 ? welem[25] : _GEN_1562; // @[Execute.scala 117:10]
  assign _GEN_1564 = 6'h1a == _T_204 ? welem[26] : _GEN_1563; // @[Execute.scala 117:10]
  assign _GEN_1565 = 6'h1b == _T_204 ? welem[27] : _GEN_1564; // @[Execute.scala 117:10]
  assign _GEN_1566 = 6'h1c == _T_204 ? welem[28] : _GEN_1565; // @[Execute.scala 117:10]
  assign _GEN_1567 = 6'h1d == _T_204 ? welem[29] : _GEN_1566; // @[Execute.scala 117:10]
  assign _GEN_1568 = 6'h1e == _T_204 ? welem[30] : _GEN_1567; // @[Execute.scala 117:10]
  assign _GEN_1569 = 6'h1f == _T_204 ? welem[31] : _GEN_1568; // @[Execute.scala 117:10]
  assign _GEN_1570 = 6'h20 == _T_204 ? welem[32] : _GEN_1569; // @[Execute.scala 117:10]
  assign _GEN_1571 = 6'h21 == _T_204 ? welem[33] : _GEN_1570; // @[Execute.scala 117:10]
  assign _GEN_1572 = 6'h22 == _T_204 ? welem[34] : _GEN_1571; // @[Execute.scala 117:10]
  assign _GEN_1573 = 6'h23 == _T_204 ? welem[35] : _GEN_1572; // @[Execute.scala 117:10]
  assign _GEN_1574 = 6'h24 == _T_204 ? welem[36] : _GEN_1573; // @[Execute.scala 117:10]
  assign _GEN_1575 = 6'h25 == _T_204 ? welem[37] : _GEN_1574; // @[Execute.scala 117:10]
  assign _GEN_1576 = 6'h26 == _T_204 ? welem[38] : _GEN_1575; // @[Execute.scala 117:10]
  assign _GEN_1577 = 6'h27 == _T_204 ? welem[39] : _GEN_1576; // @[Execute.scala 117:10]
  assign _GEN_1578 = 6'h28 == _T_204 ? welem[40] : _GEN_1577; // @[Execute.scala 117:10]
  assign _GEN_1579 = 6'h29 == _T_204 ? welem[41] : _GEN_1578; // @[Execute.scala 117:10]
  assign _GEN_1580 = 6'h2a == _T_204 ? welem[42] : _GEN_1579; // @[Execute.scala 117:10]
  assign _GEN_1581 = 6'h2b == _T_204 ? welem[43] : _GEN_1580; // @[Execute.scala 117:10]
  assign _GEN_1582 = 6'h2c == _T_204 ? welem[44] : _GEN_1581; // @[Execute.scala 117:10]
  assign _GEN_1583 = 6'h2d == _T_204 ? welem[45] : _GEN_1582; // @[Execute.scala 117:10]
  assign _GEN_1584 = 6'h2e == _T_204 ? welem[46] : _GEN_1583; // @[Execute.scala 117:10]
  assign _GEN_1585 = 6'h2f == _T_204 ? welem[47] : _GEN_1584; // @[Execute.scala 117:10]
  assign _GEN_1586 = 6'h30 == _T_204 ? welem[48] : _GEN_1585; // @[Execute.scala 117:10]
  assign _GEN_1587 = 6'h31 == _T_204 ? welem[49] : _GEN_1586; // @[Execute.scala 117:10]
  assign _GEN_1588 = 6'h32 == _T_204 ? welem[50] : _GEN_1587; // @[Execute.scala 117:10]
  assign _GEN_1589 = 6'h33 == _T_204 ? welem[51] : _GEN_1588; // @[Execute.scala 117:10]
  assign _GEN_1590 = 6'h34 == _T_204 ? welem[52] : _GEN_1589; // @[Execute.scala 117:10]
  assign _GEN_1591 = 6'h35 == _T_204 ? welem[53] : _GEN_1590; // @[Execute.scala 117:10]
  assign _GEN_1592 = 6'h36 == _T_204 ? welem[54] : _GEN_1591; // @[Execute.scala 117:10]
  assign _GEN_1593 = 6'h37 == _T_204 ? welem[55] : _GEN_1592; // @[Execute.scala 117:10]
  assign _GEN_1594 = 6'h38 == _T_204 ? welem[56] : _GEN_1593; // @[Execute.scala 117:10]
  assign _GEN_1595 = 6'h39 == _T_204 ? welem[57] : _GEN_1594; // @[Execute.scala 117:10]
  assign _GEN_1596 = 6'h3a == _T_204 ? welem[58] : _GEN_1595; // @[Execute.scala 117:10]
  assign _GEN_1597 = 6'h3b == _T_204 ? welem[59] : _GEN_1596; // @[Execute.scala 117:10]
  assign _GEN_1598 = 6'h3c == _T_204 ? welem[60] : _GEN_1597; // @[Execute.scala 117:10]
  assign _GEN_1599 = 6'h3d == _T_204 ? welem[61] : _GEN_1598; // @[Execute.scala 117:10]
  assign _GEN_1600 = 6'h3e == _T_204 ? welem[62] : _GEN_1599; // @[Execute.scala 117:10]
  assign _GEN_1601 = 6'h3f == _T_204 ? welem[63] : _GEN_1600; // @[Execute.scala 117:10]
  assign _GEN_1603 = 6'h1 == _T_208 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1604 = 6'h2 == _T_208 ? welem[2] : _GEN_1603; // @[Execute.scala 117:10]
  assign _GEN_1605 = 6'h3 == _T_208 ? welem[3] : _GEN_1604; // @[Execute.scala 117:10]
  assign _GEN_1606 = 6'h4 == _T_208 ? welem[4] : _GEN_1605; // @[Execute.scala 117:10]
  assign _GEN_1607 = 6'h5 == _T_208 ? welem[5] : _GEN_1606; // @[Execute.scala 117:10]
  assign _GEN_1608 = 6'h6 == _T_208 ? welem[6] : _GEN_1607; // @[Execute.scala 117:10]
  assign _GEN_1609 = 6'h7 == _T_208 ? welem[7] : _GEN_1608; // @[Execute.scala 117:10]
  assign _GEN_1610 = 6'h8 == _T_208 ? welem[8] : _GEN_1609; // @[Execute.scala 117:10]
  assign _GEN_1611 = 6'h9 == _T_208 ? welem[9] : _GEN_1610; // @[Execute.scala 117:10]
  assign _GEN_1612 = 6'ha == _T_208 ? welem[10] : _GEN_1611; // @[Execute.scala 117:10]
  assign _GEN_1613 = 6'hb == _T_208 ? welem[11] : _GEN_1612; // @[Execute.scala 117:10]
  assign _GEN_1614 = 6'hc == _T_208 ? welem[12] : _GEN_1613; // @[Execute.scala 117:10]
  assign _GEN_1615 = 6'hd == _T_208 ? welem[13] : _GEN_1614; // @[Execute.scala 117:10]
  assign _GEN_1616 = 6'he == _T_208 ? welem[14] : _GEN_1615; // @[Execute.scala 117:10]
  assign _GEN_1617 = 6'hf == _T_208 ? welem[15] : _GEN_1616; // @[Execute.scala 117:10]
  assign _GEN_1618 = 6'h10 == _T_208 ? welem[16] : _GEN_1617; // @[Execute.scala 117:10]
  assign _GEN_1619 = 6'h11 == _T_208 ? welem[17] : _GEN_1618; // @[Execute.scala 117:10]
  assign _GEN_1620 = 6'h12 == _T_208 ? welem[18] : _GEN_1619; // @[Execute.scala 117:10]
  assign _GEN_1621 = 6'h13 == _T_208 ? welem[19] : _GEN_1620; // @[Execute.scala 117:10]
  assign _GEN_1622 = 6'h14 == _T_208 ? welem[20] : _GEN_1621; // @[Execute.scala 117:10]
  assign _GEN_1623 = 6'h15 == _T_208 ? welem[21] : _GEN_1622; // @[Execute.scala 117:10]
  assign _GEN_1624 = 6'h16 == _T_208 ? welem[22] : _GEN_1623; // @[Execute.scala 117:10]
  assign _GEN_1625 = 6'h17 == _T_208 ? welem[23] : _GEN_1624; // @[Execute.scala 117:10]
  assign _GEN_1626 = 6'h18 == _T_208 ? welem[24] : _GEN_1625; // @[Execute.scala 117:10]
  assign _GEN_1627 = 6'h19 == _T_208 ? welem[25] : _GEN_1626; // @[Execute.scala 117:10]
  assign _GEN_1628 = 6'h1a == _T_208 ? welem[26] : _GEN_1627; // @[Execute.scala 117:10]
  assign _GEN_1629 = 6'h1b == _T_208 ? welem[27] : _GEN_1628; // @[Execute.scala 117:10]
  assign _GEN_1630 = 6'h1c == _T_208 ? welem[28] : _GEN_1629; // @[Execute.scala 117:10]
  assign _GEN_1631 = 6'h1d == _T_208 ? welem[29] : _GEN_1630; // @[Execute.scala 117:10]
  assign _GEN_1632 = 6'h1e == _T_208 ? welem[30] : _GEN_1631; // @[Execute.scala 117:10]
  assign _GEN_1633 = 6'h1f == _T_208 ? welem[31] : _GEN_1632; // @[Execute.scala 117:10]
  assign _GEN_1634 = 6'h20 == _T_208 ? welem[32] : _GEN_1633; // @[Execute.scala 117:10]
  assign _GEN_1635 = 6'h21 == _T_208 ? welem[33] : _GEN_1634; // @[Execute.scala 117:10]
  assign _GEN_1636 = 6'h22 == _T_208 ? welem[34] : _GEN_1635; // @[Execute.scala 117:10]
  assign _GEN_1637 = 6'h23 == _T_208 ? welem[35] : _GEN_1636; // @[Execute.scala 117:10]
  assign _GEN_1638 = 6'h24 == _T_208 ? welem[36] : _GEN_1637; // @[Execute.scala 117:10]
  assign _GEN_1639 = 6'h25 == _T_208 ? welem[37] : _GEN_1638; // @[Execute.scala 117:10]
  assign _GEN_1640 = 6'h26 == _T_208 ? welem[38] : _GEN_1639; // @[Execute.scala 117:10]
  assign _GEN_1641 = 6'h27 == _T_208 ? welem[39] : _GEN_1640; // @[Execute.scala 117:10]
  assign _GEN_1642 = 6'h28 == _T_208 ? welem[40] : _GEN_1641; // @[Execute.scala 117:10]
  assign _GEN_1643 = 6'h29 == _T_208 ? welem[41] : _GEN_1642; // @[Execute.scala 117:10]
  assign _GEN_1644 = 6'h2a == _T_208 ? welem[42] : _GEN_1643; // @[Execute.scala 117:10]
  assign _GEN_1645 = 6'h2b == _T_208 ? welem[43] : _GEN_1644; // @[Execute.scala 117:10]
  assign _GEN_1646 = 6'h2c == _T_208 ? welem[44] : _GEN_1645; // @[Execute.scala 117:10]
  assign _GEN_1647 = 6'h2d == _T_208 ? welem[45] : _GEN_1646; // @[Execute.scala 117:10]
  assign _GEN_1648 = 6'h2e == _T_208 ? welem[46] : _GEN_1647; // @[Execute.scala 117:10]
  assign _GEN_1649 = 6'h2f == _T_208 ? welem[47] : _GEN_1648; // @[Execute.scala 117:10]
  assign _GEN_1650 = 6'h30 == _T_208 ? welem[48] : _GEN_1649; // @[Execute.scala 117:10]
  assign _GEN_1651 = 6'h31 == _T_208 ? welem[49] : _GEN_1650; // @[Execute.scala 117:10]
  assign _GEN_1652 = 6'h32 == _T_208 ? welem[50] : _GEN_1651; // @[Execute.scala 117:10]
  assign _GEN_1653 = 6'h33 == _T_208 ? welem[51] : _GEN_1652; // @[Execute.scala 117:10]
  assign _GEN_1654 = 6'h34 == _T_208 ? welem[52] : _GEN_1653; // @[Execute.scala 117:10]
  assign _GEN_1655 = 6'h35 == _T_208 ? welem[53] : _GEN_1654; // @[Execute.scala 117:10]
  assign _GEN_1656 = 6'h36 == _T_208 ? welem[54] : _GEN_1655; // @[Execute.scala 117:10]
  assign _GEN_1657 = 6'h37 == _T_208 ? welem[55] : _GEN_1656; // @[Execute.scala 117:10]
  assign _GEN_1658 = 6'h38 == _T_208 ? welem[56] : _GEN_1657; // @[Execute.scala 117:10]
  assign _GEN_1659 = 6'h39 == _T_208 ? welem[57] : _GEN_1658; // @[Execute.scala 117:10]
  assign _GEN_1660 = 6'h3a == _T_208 ? welem[58] : _GEN_1659; // @[Execute.scala 117:10]
  assign _GEN_1661 = 6'h3b == _T_208 ? welem[59] : _GEN_1660; // @[Execute.scala 117:10]
  assign _GEN_1662 = 6'h3c == _T_208 ? welem[60] : _GEN_1661; // @[Execute.scala 117:10]
  assign _GEN_1663 = 6'h3d == _T_208 ? welem[61] : _GEN_1662; // @[Execute.scala 117:10]
  assign _GEN_1664 = 6'h3e == _T_208 ? welem[62] : _GEN_1663; // @[Execute.scala 117:10]
  assign _GEN_1665 = 6'h3f == _T_208 ? welem[63] : _GEN_1664; // @[Execute.scala 117:10]
  assign _T_211 = _T_202 ? _GEN_1601 : _GEN_1665; // @[Execute.scala 117:10]
  assign _T_212 = r < 6'h34; // @[Execute.scala 117:15]
  assign _T_214 = r - 6'h34; // @[Execute.scala 117:37]
  assign _T_218 = 6'hc + r; // @[Execute.scala 117:60]
  assign _GEN_1667 = 6'h1 == _T_214 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1668 = 6'h2 == _T_214 ? welem[2] : _GEN_1667; // @[Execute.scala 117:10]
  assign _GEN_1669 = 6'h3 == _T_214 ? welem[3] : _GEN_1668; // @[Execute.scala 117:10]
  assign _GEN_1670 = 6'h4 == _T_214 ? welem[4] : _GEN_1669; // @[Execute.scala 117:10]
  assign _GEN_1671 = 6'h5 == _T_214 ? welem[5] : _GEN_1670; // @[Execute.scala 117:10]
  assign _GEN_1672 = 6'h6 == _T_214 ? welem[6] : _GEN_1671; // @[Execute.scala 117:10]
  assign _GEN_1673 = 6'h7 == _T_214 ? welem[7] : _GEN_1672; // @[Execute.scala 117:10]
  assign _GEN_1674 = 6'h8 == _T_214 ? welem[8] : _GEN_1673; // @[Execute.scala 117:10]
  assign _GEN_1675 = 6'h9 == _T_214 ? welem[9] : _GEN_1674; // @[Execute.scala 117:10]
  assign _GEN_1676 = 6'ha == _T_214 ? welem[10] : _GEN_1675; // @[Execute.scala 117:10]
  assign _GEN_1677 = 6'hb == _T_214 ? welem[11] : _GEN_1676; // @[Execute.scala 117:10]
  assign _GEN_1678 = 6'hc == _T_214 ? welem[12] : _GEN_1677; // @[Execute.scala 117:10]
  assign _GEN_1679 = 6'hd == _T_214 ? welem[13] : _GEN_1678; // @[Execute.scala 117:10]
  assign _GEN_1680 = 6'he == _T_214 ? welem[14] : _GEN_1679; // @[Execute.scala 117:10]
  assign _GEN_1681 = 6'hf == _T_214 ? welem[15] : _GEN_1680; // @[Execute.scala 117:10]
  assign _GEN_1682 = 6'h10 == _T_214 ? welem[16] : _GEN_1681; // @[Execute.scala 117:10]
  assign _GEN_1683 = 6'h11 == _T_214 ? welem[17] : _GEN_1682; // @[Execute.scala 117:10]
  assign _GEN_1684 = 6'h12 == _T_214 ? welem[18] : _GEN_1683; // @[Execute.scala 117:10]
  assign _GEN_1685 = 6'h13 == _T_214 ? welem[19] : _GEN_1684; // @[Execute.scala 117:10]
  assign _GEN_1686 = 6'h14 == _T_214 ? welem[20] : _GEN_1685; // @[Execute.scala 117:10]
  assign _GEN_1687 = 6'h15 == _T_214 ? welem[21] : _GEN_1686; // @[Execute.scala 117:10]
  assign _GEN_1688 = 6'h16 == _T_214 ? welem[22] : _GEN_1687; // @[Execute.scala 117:10]
  assign _GEN_1689 = 6'h17 == _T_214 ? welem[23] : _GEN_1688; // @[Execute.scala 117:10]
  assign _GEN_1690 = 6'h18 == _T_214 ? welem[24] : _GEN_1689; // @[Execute.scala 117:10]
  assign _GEN_1691 = 6'h19 == _T_214 ? welem[25] : _GEN_1690; // @[Execute.scala 117:10]
  assign _GEN_1692 = 6'h1a == _T_214 ? welem[26] : _GEN_1691; // @[Execute.scala 117:10]
  assign _GEN_1693 = 6'h1b == _T_214 ? welem[27] : _GEN_1692; // @[Execute.scala 117:10]
  assign _GEN_1694 = 6'h1c == _T_214 ? welem[28] : _GEN_1693; // @[Execute.scala 117:10]
  assign _GEN_1695 = 6'h1d == _T_214 ? welem[29] : _GEN_1694; // @[Execute.scala 117:10]
  assign _GEN_1696 = 6'h1e == _T_214 ? welem[30] : _GEN_1695; // @[Execute.scala 117:10]
  assign _GEN_1697 = 6'h1f == _T_214 ? welem[31] : _GEN_1696; // @[Execute.scala 117:10]
  assign _GEN_1698 = 6'h20 == _T_214 ? welem[32] : _GEN_1697; // @[Execute.scala 117:10]
  assign _GEN_1699 = 6'h21 == _T_214 ? welem[33] : _GEN_1698; // @[Execute.scala 117:10]
  assign _GEN_1700 = 6'h22 == _T_214 ? welem[34] : _GEN_1699; // @[Execute.scala 117:10]
  assign _GEN_1701 = 6'h23 == _T_214 ? welem[35] : _GEN_1700; // @[Execute.scala 117:10]
  assign _GEN_1702 = 6'h24 == _T_214 ? welem[36] : _GEN_1701; // @[Execute.scala 117:10]
  assign _GEN_1703 = 6'h25 == _T_214 ? welem[37] : _GEN_1702; // @[Execute.scala 117:10]
  assign _GEN_1704 = 6'h26 == _T_214 ? welem[38] : _GEN_1703; // @[Execute.scala 117:10]
  assign _GEN_1705 = 6'h27 == _T_214 ? welem[39] : _GEN_1704; // @[Execute.scala 117:10]
  assign _GEN_1706 = 6'h28 == _T_214 ? welem[40] : _GEN_1705; // @[Execute.scala 117:10]
  assign _GEN_1707 = 6'h29 == _T_214 ? welem[41] : _GEN_1706; // @[Execute.scala 117:10]
  assign _GEN_1708 = 6'h2a == _T_214 ? welem[42] : _GEN_1707; // @[Execute.scala 117:10]
  assign _GEN_1709 = 6'h2b == _T_214 ? welem[43] : _GEN_1708; // @[Execute.scala 117:10]
  assign _GEN_1710 = 6'h2c == _T_214 ? welem[44] : _GEN_1709; // @[Execute.scala 117:10]
  assign _GEN_1711 = 6'h2d == _T_214 ? welem[45] : _GEN_1710; // @[Execute.scala 117:10]
  assign _GEN_1712 = 6'h2e == _T_214 ? welem[46] : _GEN_1711; // @[Execute.scala 117:10]
  assign _GEN_1713 = 6'h2f == _T_214 ? welem[47] : _GEN_1712; // @[Execute.scala 117:10]
  assign _GEN_1714 = 6'h30 == _T_214 ? welem[48] : _GEN_1713; // @[Execute.scala 117:10]
  assign _GEN_1715 = 6'h31 == _T_214 ? welem[49] : _GEN_1714; // @[Execute.scala 117:10]
  assign _GEN_1716 = 6'h32 == _T_214 ? welem[50] : _GEN_1715; // @[Execute.scala 117:10]
  assign _GEN_1717 = 6'h33 == _T_214 ? welem[51] : _GEN_1716; // @[Execute.scala 117:10]
  assign _GEN_1718 = 6'h34 == _T_214 ? welem[52] : _GEN_1717; // @[Execute.scala 117:10]
  assign _GEN_1719 = 6'h35 == _T_214 ? welem[53] : _GEN_1718; // @[Execute.scala 117:10]
  assign _GEN_1720 = 6'h36 == _T_214 ? welem[54] : _GEN_1719; // @[Execute.scala 117:10]
  assign _GEN_1721 = 6'h37 == _T_214 ? welem[55] : _GEN_1720; // @[Execute.scala 117:10]
  assign _GEN_1722 = 6'h38 == _T_214 ? welem[56] : _GEN_1721; // @[Execute.scala 117:10]
  assign _GEN_1723 = 6'h39 == _T_214 ? welem[57] : _GEN_1722; // @[Execute.scala 117:10]
  assign _GEN_1724 = 6'h3a == _T_214 ? welem[58] : _GEN_1723; // @[Execute.scala 117:10]
  assign _GEN_1725 = 6'h3b == _T_214 ? welem[59] : _GEN_1724; // @[Execute.scala 117:10]
  assign _GEN_1726 = 6'h3c == _T_214 ? welem[60] : _GEN_1725; // @[Execute.scala 117:10]
  assign _GEN_1727 = 6'h3d == _T_214 ? welem[61] : _GEN_1726; // @[Execute.scala 117:10]
  assign _GEN_1728 = 6'h3e == _T_214 ? welem[62] : _GEN_1727; // @[Execute.scala 117:10]
  assign _GEN_1729 = 6'h3f == _T_214 ? welem[63] : _GEN_1728; // @[Execute.scala 117:10]
  assign _GEN_1731 = 6'h1 == _T_218 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1732 = 6'h2 == _T_218 ? welem[2] : _GEN_1731; // @[Execute.scala 117:10]
  assign _GEN_1733 = 6'h3 == _T_218 ? welem[3] : _GEN_1732; // @[Execute.scala 117:10]
  assign _GEN_1734 = 6'h4 == _T_218 ? welem[4] : _GEN_1733; // @[Execute.scala 117:10]
  assign _GEN_1735 = 6'h5 == _T_218 ? welem[5] : _GEN_1734; // @[Execute.scala 117:10]
  assign _GEN_1736 = 6'h6 == _T_218 ? welem[6] : _GEN_1735; // @[Execute.scala 117:10]
  assign _GEN_1737 = 6'h7 == _T_218 ? welem[7] : _GEN_1736; // @[Execute.scala 117:10]
  assign _GEN_1738 = 6'h8 == _T_218 ? welem[8] : _GEN_1737; // @[Execute.scala 117:10]
  assign _GEN_1739 = 6'h9 == _T_218 ? welem[9] : _GEN_1738; // @[Execute.scala 117:10]
  assign _GEN_1740 = 6'ha == _T_218 ? welem[10] : _GEN_1739; // @[Execute.scala 117:10]
  assign _GEN_1741 = 6'hb == _T_218 ? welem[11] : _GEN_1740; // @[Execute.scala 117:10]
  assign _GEN_1742 = 6'hc == _T_218 ? welem[12] : _GEN_1741; // @[Execute.scala 117:10]
  assign _GEN_1743 = 6'hd == _T_218 ? welem[13] : _GEN_1742; // @[Execute.scala 117:10]
  assign _GEN_1744 = 6'he == _T_218 ? welem[14] : _GEN_1743; // @[Execute.scala 117:10]
  assign _GEN_1745 = 6'hf == _T_218 ? welem[15] : _GEN_1744; // @[Execute.scala 117:10]
  assign _GEN_1746 = 6'h10 == _T_218 ? welem[16] : _GEN_1745; // @[Execute.scala 117:10]
  assign _GEN_1747 = 6'h11 == _T_218 ? welem[17] : _GEN_1746; // @[Execute.scala 117:10]
  assign _GEN_1748 = 6'h12 == _T_218 ? welem[18] : _GEN_1747; // @[Execute.scala 117:10]
  assign _GEN_1749 = 6'h13 == _T_218 ? welem[19] : _GEN_1748; // @[Execute.scala 117:10]
  assign _GEN_1750 = 6'h14 == _T_218 ? welem[20] : _GEN_1749; // @[Execute.scala 117:10]
  assign _GEN_1751 = 6'h15 == _T_218 ? welem[21] : _GEN_1750; // @[Execute.scala 117:10]
  assign _GEN_1752 = 6'h16 == _T_218 ? welem[22] : _GEN_1751; // @[Execute.scala 117:10]
  assign _GEN_1753 = 6'h17 == _T_218 ? welem[23] : _GEN_1752; // @[Execute.scala 117:10]
  assign _GEN_1754 = 6'h18 == _T_218 ? welem[24] : _GEN_1753; // @[Execute.scala 117:10]
  assign _GEN_1755 = 6'h19 == _T_218 ? welem[25] : _GEN_1754; // @[Execute.scala 117:10]
  assign _GEN_1756 = 6'h1a == _T_218 ? welem[26] : _GEN_1755; // @[Execute.scala 117:10]
  assign _GEN_1757 = 6'h1b == _T_218 ? welem[27] : _GEN_1756; // @[Execute.scala 117:10]
  assign _GEN_1758 = 6'h1c == _T_218 ? welem[28] : _GEN_1757; // @[Execute.scala 117:10]
  assign _GEN_1759 = 6'h1d == _T_218 ? welem[29] : _GEN_1758; // @[Execute.scala 117:10]
  assign _GEN_1760 = 6'h1e == _T_218 ? welem[30] : _GEN_1759; // @[Execute.scala 117:10]
  assign _GEN_1761 = 6'h1f == _T_218 ? welem[31] : _GEN_1760; // @[Execute.scala 117:10]
  assign _GEN_1762 = 6'h20 == _T_218 ? welem[32] : _GEN_1761; // @[Execute.scala 117:10]
  assign _GEN_1763 = 6'h21 == _T_218 ? welem[33] : _GEN_1762; // @[Execute.scala 117:10]
  assign _GEN_1764 = 6'h22 == _T_218 ? welem[34] : _GEN_1763; // @[Execute.scala 117:10]
  assign _GEN_1765 = 6'h23 == _T_218 ? welem[35] : _GEN_1764; // @[Execute.scala 117:10]
  assign _GEN_1766 = 6'h24 == _T_218 ? welem[36] : _GEN_1765; // @[Execute.scala 117:10]
  assign _GEN_1767 = 6'h25 == _T_218 ? welem[37] : _GEN_1766; // @[Execute.scala 117:10]
  assign _GEN_1768 = 6'h26 == _T_218 ? welem[38] : _GEN_1767; // @[Execute.scala 117:10]
  assign _GEN_1769 = 6'h27 == _T_218 ? welem[39] : _GEN_1768; // @[Execute.scala 117:10]
  assign _GEN_1770 = 6'h28 == _T_218 ? welem[40] : _GEN_1769; // @[Execute.scala 117:10]
  assign _GEN_1771 = 6'h29 == _T_218 ? welem[41] : _GEN_1770; // @[Execute.scala 117:10]
  assign _GEN_1772 = 6'h2a == _T_218 ? welem[42] : _GEN_1771; // @[Execute.scala 117:10]
  assign _GEN_1773 = 6'h2b == _T_218 ? welem[43] : _GEN_1772; // @[Execute.scala 117:10]
  assign _GEN_1774 = 6'h2c == _T_218 ? welem[44] : _GEN_1773; // @[Execute.scala 117:10]
  assign _GEN_1775 = 6'h2d == _T_218 ? welem[45] : _GEN_1774; // @[Execute.scala 117:10]
  assign _GEN_1776 = 6'h2e == _T_218 ? welem[46] : _GEN_1775; // @[Execute.scala 117:10]
  assign _GEN_1777 = 6'h2f == _T_218 ? welem[47] : _GEN_1776; // @[Execute.scala 117:10]
  assign _GEN_1778 = 6'h30 == _T_218 ? welem[48] : _GEN_1777; // @[Execute.scala 117:10]
  assign _GEN_1779 = 6'h31 == _T_218 ? welem[49] : _GEN_1778; // @[Execute.scala 117:10]
  assign _GEN_1780 = 6'h32 == _T_218 ? welem[50] : _GEN_1779; // @[Execute.scala 117:10]
  assign _GEN_1781 = 6'h33 == _T_218 ? welem[51] : _GEN_1780; // @[Execute.scala 117:10]
  assign _GEN_1782 = 6'h34 == _T_218 ? welem[52] : _GEN_1781; // @[Execute.scala 117:10]
  assign _GEN_1783 = 6'h35 == _T_218 ? welem[53] : _GEN_1782; // @[Execute.scala 117:10]
  assign _GEN_1784 = 6'h36 == _T_218 ? welem[54] : _GEN_1783; // @[Execute.scala 117:10]
  assign _GEN_1785 = 6'h37 == _T_218 ? welem[55] : _GEN_1784; // @[Execute.scala 117:10]
  assign _GEN_1786 = 6'h38 == _T_218 ? welem[56] : _GEN_1785; // @[Execute.scala 117:10]
  assign _GEN_1787 = 6'h39 == _T_218 ? welem[57] : _GEN_1786; // @[Execute.scala 117:10]
  assign _GEN_1788 = 6'h3a == _T_218 ? welem[58] : _GEN_1787; // @[Execute.scala 117:10]
  assign _GEN_1789 = 6'h3b == _T_218 ? welem[59] : _GEN_1788; // @[Execute.scala 117:10]
  assign _GEN_1790 = 6'h3c == _T_218 ? welem[60] : _GEN_1789; // @[Execute.scala 117:10]
  assign _GEN_1791 = 6'h3d == _T_218 ? welem[61] : _GEN_1790; // @[Execute.scala 117:10]
  assign _GEN_1792 = 6'h3e == _T_218 ? welem[62] : _GEN_1791; // @[Execute.scala 117:10]
  assign _GEN_1793 = 6'h3f == _T_218 ? welem[63] : _GEN_1792; // @[Execute.scala 117:10]
  assign _T_221 = _T_212 ? _GEN_1729 : _GEN_1793; // @[Execute.scala 117:10]
  assign _T_222 = r < 6'h33; // @[Execute.scala 117:15]
  assign _T_224 = r - 6'h33; // @[Execute.scala 117:37]
  assign _T_228 = 6'hd + r; // @[Execute.scala 117:60]
  assign _GEN_1795 = 6'h1 == _T_224 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1796 = 6'h2 == _T_224 ? welem[2] : _GEN_1795; // @[Execute.scala 117:10]
  assign _GEN_1797 = 6'h3 == _T_224 ? welem[3] : _GEN_1796; // @[Execute.scala 117:10]
  assign _GEN_1798 = 6'h4 == _T_224 ? welem[4] : _GEN_1797; // @[Execute.scala 117:10]
  assign _GEN_1799 = 6'h5 == _T_224 ? welem[5] : _GEN_1798; // @[Execute.scala 117:10]
  assign _GEN_1800 = 6'h6 == _T_224 ? welem[6] : _GEN_1799; // @[Execute.scala 117:10]
  assign _GEN_1801 = 6'h7 == _T_224 ? welem[7] : _GEN_1800; // @[Execute.scala 117:10]
  assign _GEN_1802 = 6'h8 == _T_224 ? welem[8] : _GEN_1801; // @[Execute.scala 117:10]
  assign _GEN_1803 = 6'h9 == _T_224 ? welem[9] : _GEN_1802; // @[Execute.scala 117:10]
  assign _GEN_1804 = 6'ha == _T_224 ? welem[10] : _GEN_1803; // @[Execute.scala 117:10]
  assign _GEN_1805 = 6'hb == _T_224 ? welem[11] : _GEN_1804; // @[Execute.scala 117:10]
  assign _GEN_1806 = 6'hc == _T_224 ? welem[12] : _GEN_1805; // @[Execute.scala 117:10]
  assign _GEN_1807 = 6'hd == _T_224 ? welem[13] : _GEN_1806; // @[Execute.scala 117:10]
  assign _GEN_1808 = 6'he == _T_224 ? welem[14] : _GEN_1807; // @[Execute.scala 117:10]
  assign _GEN_1809 = 6'hf == _T_224 ? welem[15] : _GEN_1808; // @[Execute.scala 117:10]
  assign _GEN_1810 = 6'h10 == _T_224 ? welem[16] : _GEN_1809; // @[Execute.scala 117:10]
  assign _GEN_1811 = 6'h11 == _T_224 ? welem[17] : _GEN_1810; // @[Execute.scala 117:10]
  assign _GEN_1812 = 6'h12 == _T_224 ? welem[18] : _GEN_1811; // @[Execute.scala 117:10]
  assign _GEN_1813 = 6'h13 == _T_224 ? welem[19] : _GEN_1812; // @[Execute.scala 117:10]
  assign _GEN_1814 = 6'h14 == _T_224 ? welem[20] : _GEN_1813; // @[Execute.scala 117:10]
  assign _GEN_1815 = 6'h15 == _T_224 ? welem[21] : _GEN_1814; // @[Execute.scala 117:10]
  assign _GEN_1816 = 6'h16 == _T_224 ? welem[22] : _GEN_1815; // @[Execute.scala 117:10]
  assign _GEN_1817 = 6'h17 == _T_224 ? welem[23] : _GEN_1816; // @[Execute.scala 117:10]
  assign _GEN_1818 = 6'h18 == _T_224 ? welem[24] : _GEN_1817; // @[Execute.scala 117:10]
  assign _GEN_1819 = 6'h19 == _T_224 ? welem[25] : _GEN_1818; // @[Execute.scala 117:10]
  assign _GEN_1820 = 6'h1a == _T_224 ? welem[26] : _GEN_1819; // @[Execute.scala 117:10]
  assign _GEN_1821 = 6'h1b == _T_224 ? welem[27] : _GEN_1820; // @[Execute.scala 117:10]
  assign _GEN_1822 = 6'h1c == _T_224 ? welem[28] : _GEN_1821; // @[Execute.scala 117:10]
  assign _GEN_1823 = 6'h1d == _T_224 ? welem[29] : _GEN_1822; // @[Execute.scala 117:10]
  assign _GEN_1824 = 6'h1e == _T_224 ? welem[30] : _GEN_1823; // @[Execute.scala 117:10]
  assign _GEN_1825 = 6'h1f == _T_224 ? welem[31] : _GEN_1824; // @[Execute.scala 117:10]
  assign _GEN_1826 = 6'h20 == _T_224 ? welem[32] : _GEN_1825; // @[Execute.scala 117:10]
  assign _GEN_1827 = 6'h21 == _T_224 ? welem[33] : _GEN_1826; // @[Execute.scala 117:10]
  assign _GEN_1828 = 6'h22 == _T_224 ? welem[34] : _GEN_1827; // @[Execute.scala 117:10]
  assign _GEN_1829 = 6'h23 == _T_224 ? welem[35] : _GEN_1828; // @[Execute.scala 117:10]
  assign _GEN_1830 = 6'h24 == _T_224 ? welem[36] : _GEN_1829; // @[Execute.scala 117:10]
  assign _GEN_1831 = 6'h25 == _T_224 ? welem[37] : _GEN_1830; // @[Execute.scala 117:10]
  assign _GEN_1832 = 6'h26 == _T_224 ? welem[38] : _GEN_1831; // @[Execute.scala 117:10]
  assign _GEN_1833 = 6'h27 == _T_224 ? welem[39] : _GEN_1832; // @[Execute.scala 117:10]
  assign _GEN_1834 = 6'h28 == _T_224 ? welem[40] : _GEN_1833; // @[Execute.scala 117:10]
  assign _GEN_1835 = 6'h29 == _T_224 ? welem[41] : _GEN_1834; // @[Execute.scala 117:10]
  assign _GEN_1836 = 6'h2a == _T_224 ? welem[42] : _GEN_1835; // @[Execute.scala 117:10]
  assign _GEN_1837 = 6'h2b == _T_224 ? welem[43] : _GEN_1836; // @[Execute.scala 117:10]
  assign _GEN_1838 = 6'h2c == _T_224 ? welem[44] : _GEN_1837; // @[Execute.scala 117:10]
  assign _GEN_1839 = 6'h2d == _T_224 ? welem[45] : _GEN_1838; // @[Execute.scala 117:10]
  assign _GEN_1840 = 6'h2e == _T_224 ? welem[46] : _GEN_1839; // @[Execute.scala 117:10]
  assign _GEN_1841 = 6'h2f == _T_224 ? welem[47] : _GEN_1840; // @[Execute.scala 117:10]
  assign _GEN_1842 = 6'h30 == _T_224 ? welem[48] : _GEN_1841; // @[Execute.scala 117:10]
  assign _GEN_1843 = 6'h31 == _T_224 ? welem[49] : _GEN_1842; // @[Execute.scala 117:10]
  assign _GEN_1844 = 6'h32 == _T_224 ? welem[50] : _GEN_1843; // @[Execute.scala 117:10]
  assign _GEN_1845 = 6'h33 == _T_224 ? welem[51] : _GEN_1844; // @[Execute.scala 117:10]
  assign _GEN_1846 = 6'h34 == _T_224 ? welem[52] : _GEN_1845; // @[Execute.scala 117:10]
  assign _GEN_1847 = 6'h35 == _T_224 ? welem[53] : _GEN_1846; // @[Execute.scala 117:10]
  assign _GEN_1848 = 6'h36 == _T_224 ? welem[54] : _GEN_1847; // @[Execute.scala 117:10]
  assign _GEN_1849 = 6'h37 == _T_224 ? welem[55] : _GEN_1848; // @[Execute.scala 117:10]
  assign _GEN_1850 = 6'h38 == _T_224 ? welem[56] : _GEN_1849; // @[Execute.scala 117:10]
  assign _GEN_1851 = 6'h39 == _T_224 ? welem[57] : _GEN_1850; // @[Execute.scala 117:10]
  assign _GEN_1852 = 6'h3a == _T_224 ? welem[58] : _GEN_1851; // @[Execute.scala 117:10]
  assign _GEN_1853 = 6'h3b == _T_224 ? welem[59] : _GEN_1852; // @[Execute.scala 117:10]
  assign _GEN_1854 = 6'h3c == _T_224 ? welem[60] : _GEN_1853; // @[Execute.scala 117:10]
  assign _GEN_1855 = 6'h3d == _T_224 ? welem[61] : _GEN_1854; // @[Execute.scala 117:10]
  assign _GEN_1856 = 6'h3e == _T_224 ? welem[62] : _GEN_1855; // @[Execute.scala 117:10]
  assign _GEN_1857 = 6'h3f == _T_224 ? welem[63] : _GEN_1856; // @[Execute.scala 117:10]
  assign _GEN_1859 = 6'h1 == _T_228 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1860 = 6'h2 == _T_228 ? welem[2] : _GEN_1859; // @[Execute.scala 117:10]
  assign _GEN_1861 = 6'h3 == _T_228 ? welem[3] : _GEN_1860; // @[Execute.scala 117:10]
  assign _GEN_1862 = 6'h4 == _T_228 ? welem[4] : _GEN_1861; // @[Execute.scala 117:10]
  assign _GEN_1863 = 6'h5 == _T_228 ? welem[5] : _GEN_1862; // @[Execute.scala 117:10]
  assign _GEN_1864 = 6'h6 == _T_228 ? welem[6] : _GEN_1863; // @[Execute.scala 117:10]
  assign _GEN_1865 = 6'h7 == _T_228 ? welem[7] : _GEN_1864; // @[Execute.scala 117:10]
  assign _GEN_1866 = 6'h8 == _T_228 ? welem[8] : _GEN_1865; // @[Execute.scala 117:10]
  assign _GEN_1867 = 6'h9 == _T_228 ? welem[9] : _GEN_1866; // @[Execute.scala 117:10]
  assign _GEN_1868 = 6'ha == _T_228 ? welem[10] : _GEN_1867; // @[Execute.scala 117:10]
  assign _GEN_1869 = 6'hb == _T_228 ? welem[11] : _GEN_1868; // @[Execute.scala 117:10]
  assign _GEN_1870 = 6'hc == _T_228 ? welem[12] : _GEN_1869; // @[Execute.scala 117:10]
  assign _GEN_1871 = 6'hd == _T_228 ? welem[13] : _GEN_1870; // @[Execute.scala 117:10]
  assign _GEN_1872 = 6'he == _T_228 ? welem[14] : _GEN_1871; // @[Execute.scala 117:10]
  assign _GEN_1873 = 6'hf == _T_228 ? welem[15] : _GEN_1872; // @[Execute.scala 117:10]
  assign _GEN_1874 = 6'h10 == _T_228 ? welem[16] : _GEN_1873; // @[Execute.scala 117:10]
  assign _GEN_1875 = 6'h11 == _T_228 ? welem[17] : _GEN_1874; // @[Execute.scala 117:10]
  assign _GEN_1876 = 6'h12 == _T_228 ? welem[18] : _GEN_1875; // @[Execute.scala 117:10]
  assign _GEN_1877 = 6'h13 == _T_228 ? welem[19] : _GEN_1876; // @[Execute.scala 117:10]
  assign _GEN_1878 = 6'h14 == _T_228 ? welem[20] : _GEN_1877; // @[Execute.scala 117:10]
  assign _GEN_1879 = 6'h15 == _T_228 ? welem[21] : _GEN_1878; // @[Execute.scala 117:10]
  assign _GEN_1880 = 6'h16 == _T_228 ? welem[22] : _GEN_1879; // @[Execute.scala 117:10]
  assign _GEN_1881 = 6'h17 == _T_228 ? welem[23] : _GEN_1880; // @[Execute.scala 117:10]
  assign _GEN_1882 = 6'h18 == _T_228 ? welem[24] : _GEN_1881; // @[Execute.scala 117:10]
  assign _GEN_1883 = 6'h19 == _T_228 ? welem[25] : _GEN_1882; // @[Execute.scala 117:10]
  assign _GEN_1884 = 6'h1a == _T_228 ? welem[26] : _GEN_1883; // @[Execute.scala 117:10]
  assign _GEN_1885 = 6'h1b == _T_228 ? welem[27] : _GEN_1884; // @[Execute.scala 117:10]
  assign _GEN_1886 = 6'h1c == _T_228 ? welem[28] : _GEN_1885; // @[Execute.scala 117:10]
  assign _GEN_1887 = 6'h1d == _T_228 ? welem[29] : _GEN_1886; // @[Execute.scala 117:10]
  assign _GEN_1888 = 6'h1e == _T_228 ? welem[30] : _GEN_1887; // @[Execute.scala 117:10]
  assign _GEN_1889 = 6'h1f == _T_228 ? welem[31] : _GEN_1888; // @[Execute.scala 117:10]
  assign _GEN_1890 = 6'h20 == _T_228 ? welem[32] : _GEN_1889; // @[Execute.scala 117:10]
  assign _GEN_1891 = 6'h21 == _T_228 ? welem[33] : _GEN_1890; // @[Execute.scala 117:10]
  assign _GEN_1892 = 6'h22 == _T_228 ? welem[34] : _GEN_1891; // @[Execute.scala 117:10]
  assign _GEN_1893 = 6'h23 == _T_228 ? welem[35] : _GEN_1892; // @[Execute.scala 117:10]
  assign _GEN_1894 = 6'h24 == _T_228 ? welem[36] : _GEN_1893; // @[Execute.scala 117:10]
  assign _GEN_1895 = 6'h25 == _T_228 ? welem[37] : _GEN_1894; // @[Execute.scala 117:10]
  assign _GEN_1896 = 6'h26 == _T_228 ? welem[38] : _GEN_1895; // @[Execute.scala 117:10]
  assign _GEN_1897 = 6'h27 == _T_228 ? welem[39] : _GEN_1896; // @[Execute.scala 117:10]
  assign _GEN_1898 = 6'h28 == _T_228 ? welem[40] : _GEN_1897; // @[Execute.scala 117:10]
  assign _GEN_1899 = 6'h29 == _T_228 ? welem[41] : _GEN_1898; // @[Execute.scala 117:10]
  assign _GEN_1900 = 6'h2a == _T_228 ? welem[42] : _GEN_1899; // @[Execute.scala 117:10]
  assign _GEN_1901 = 6'h2b == _T_228 ? welem[43] : _GEN_1900; // @[Execute.scala 117:10]
  assign _GEN_1902 = 6'h2c == _T_228 ? welem[44] : _GEN_1901; // @[Execute.scala 117:10]
  assign _GEN_1903 = 6'h2d == _T_228 ? welem[45] : _GEN_1902; // @[Execute.scala 117:10]
  assign _GEN_1904 = 6'h2e == _T_228 ? welem[46] : _GEN_1903; // @[Execute.scala 117:10]
  assign _GEN_1905 = 6'h2f == _T_228 ? welem[47] : _GEN_1904; // @[Execute.scala 117:10]
  assign _GEN_1906 = 6'h30 == _T_228 ? welem[48] : _GEN_1905; // @[Execute.scala 117:10]
  assign _GEN_1907 = 6'h31 == _T_228 ? welem[49] : _GEN_1906; // @[Execute.scala 117:10]
  assign _GEN_1908 = 6'h32 == _T_228 ? welem[50] : _GEN_1907; // @[Execute.scala 117:10]
  assign _GEN_1909 = 6'h33 == _T_228 ? welem[51] : _GEN_1908; // @[Execute.scala 117:10]
  assign _GEN_1910 = 6'h34 == _T_228 ? welem[52] : _GEN_1909; // @[Execute.scala 117:10]
  assign _GEN_1911 = 6'h35 == _T_228 ? welem[53] : _GEN_1910; // @[Execute.scala 117:10]
  assign _GEN_1912 = 6'h36 == _T_228 ? welem[54] : _GEN_1911; // @[Execute.scala 117:10]
  assign _GEN_1913 = 6'h37 == _T_228 ? welem[55] : _GEN_1912; // @[Execute.scala 117:10]
  assign _GEN_1914 = 6'h38 == _T_228 ? welem[56] : _GEN_1913; // @[Execute.scala 117:10]
  assign _GEN_1915 = 6'h39 == _T_228 ? welem[57] : _GEN_1914; // @[Execute.scala 117:10]
  assign _GEN_1916 = 6'h3a == _T_228 ? welem[58] : _GEN_1915; // @[Execute.scala 117:10]
  assign _GEN_1917 = 6'h3b == _T_228 ? welem[59] : _GEN_1916; // @[Execute.scala 117:10]
  assign _GEN_1918 = 6'h3c == _T_228 ? welem[60] : _GEN_1917; // @[Execute.scala 117:10]
  assign _GEN_1919 = 6'h3d == _T_228 ? welem[61] : _GEN_1918; // @[Execute.scala 117:10]
  assign _GEN_1920 = 6'h3e == _T_228 ? welem[62] : _GEN_1919; // @[Execute.scala 117:10]
  assign _GEN_1921 = 6'h3f == _T_228 ? welem[63] : _GEN_1920; // @[Execute.scala 117:10]
  assign _T_231 = _T_222 ? _GEN_1857 : _GEN_1921; // @[Execute.scala 117:10]
  assign _T_232 = r < 6'h32; // @[Execute.scala 117:15]
  assign _T_234 = r - 6'h32; // @[Execute.scala 117:37]
  assign _T_238 = 6'he + r; // @[Execute.scala 117:60]
  assign _GEN_1923 = 6'h1 == _T_234 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1924 = 6'h2 == _T_234 ? welem[2] : _GEN_1923; // @[Execute.scala 117:10]
  assign _GEN_1925 = 6'h3 == _T_234 ? welem[3] : _GEN_1924; // @[Execute.scala 117:10]
  assign _GEN_1926 = 6'h4 == _T_234 ? welem[4] : _GEN_1925; // @[Execute.scala 117:10]
  assign _GEN_1927 = 6'h5 == _T_234 ? welem[5] : _GEN_1926; // @[Execute.scala 117:10]
  assign _GEN_1928 = 6'h6 == _T_234 ? welem[6] : _GEN_1927; // @[Execute.scala 117:10]
  assign _GEN_1929 = 6'h7 == _T_234 ? welem[7] : _GEN_1928; // @[Execute.scala 117:10]
  assign _GEN_1930 = 6'h8 == _T_234 ? welem[8] : _GEN_1929; // @[Execute.scala 117:10]
  assign _GEN_1931 = 6'h9 == _T_234 ? welem[9] : _GEN_1930; // @[Execute.scala 117:10]
  assign _GEN_1932 = 6'ha == _T_234 ? welem[10] : _GEN_1931; // @[Execute.scala 117:10]
  assign _GEN_1933 = 6'hb == _T_234 ? welem[11] : _GEN_1932; // @[Execute.scala 117:10]
  assign _GEN_1934 = 6'hc == _T_234 ? welem[12] : _GEN_1933; // @[Execute.scala 117:10]
  assign _GEN_1935 = 6'hd == _T_234 ? welem[13] : _GEN_1934; // @[Execute.scala 117:10]
  assign _GEN_1936 = 6'he == _T_234 ? welem[14] : _GEN_1935; // @[Execute.scala 117:10]
  assign _GEN_1937 = 6'hf == _T_234 ? welem[15] : _GEN_1936; // @[Execute.scala 117:10]
  assign _GEN_1938 = 6'h10 == _T_234 ? welem[16] : _GEN_1937; // @[Execute.scala 117:10]
  assign _GEN_1939 = 6'h11 == _T_234 ? welem[17] : _GEN_1938; // @[Execute.scala 117:10]
  assign _GEN_1940 = 6'h12 == _T_234 ? welem[18] : _GEN_1939; // @[Execute.scala 117:10]
  assign _GEN_1941 = 6'h13 == _T_234 ? welem[19] : _GEN_1940; // @[Execute.scala 117:10]
  assign _GEN_1942 = 6'h14 == _T_234 ? welem[20] : _GEN_1941; // @[Execute.scala 117:10]
  assign _GEN_1943 = 6'h15 == _T_234 ? welem[21] : _GEN_1942; // @[Execute.scala 117:10]
  assign _GEN_1944 = 6'h16 == _T_234 ? welem[22] : _GEN_1943; // @[Execute.scala 117:10]
  assign _GEN_1945 = 6'h17 == _T_234 ? welem[23] : _GEN_1944; // @[Execute.scala 117:10]
  assign _GEN_1946 = 6'h18 == _T_234 ? welem[24] : _GEN_1945; // @[Execute.scala 117:10]
  assign _GEN_1947 = 6'h19 == _T_234 ? welem[25] : _GEN_1946; // @[Execute.scala 117:10]
  assign _GEN_1948 = 6'h1a == _T_234 ? welem[26] : _GEN_1947; // @[Execute.scala 117:10]
  assign _GEN_1949 = 6'h1b == _T_234 ? welem[27] : _GEN_1948; // @[Execute.scala 117:10]
  assign _GEN_1950 = 6'h1c == _T_234 ? welem[28] : _GEN_1949; // @[Execute.scala 117:10]
  assign _GEN_1951 = 6'h1d == _T_234 ? welem[29] : _GEN_1950; // @[Execute.scala 117:10]
  assign _GEN_1952 = 6'h1e == _T_234 ? welem[30] : _GEN_1951; // @[Execute.scala 117:10]
  assign _GEN_1953 = 6'h1f == _T_234 ? welem[31] : _GEN_1952; // @[Execute.scala 117:10]
  assign _GEN_1954 = 6'h20 == _T_234 ? welem[32] : _GEN_1953; // @[Execute.scala 117:10]
  assign _GEN_1955 = 6'h21 == _T_234 ? welem[33] : _GEN_1954; // @[Execute.scala 117:10]
  assign _GEN_1956 = 6'h22 == _T_234 ? welem[34] : _GEN_1955; // @[Execute.scala 117:10]
  assign _GEN_1957 = 6'h23 == _T_234 ? welem[35] : _GEN_1956; // @[Execute.scala 117:10]
  assign _GEN_1958 = 6'h24 == _T_234 ? welem[36] : _GEN_1957; // @[Execute.scala 117:10]
  assign _GEN_1959 = 6'h25 == _T_234 ? welem[37] : _GEN_1958; // @[Execute.scala 117:10]
  assign _GEN_1960 = 6'h26 == _T_234 ? welem[38] : _GEN_1959; // @[Execute.scala 117:10]
  assign _GEN_1961 = 6'h27 == _T_234 ? welem[39] : _GEN_1960; // @[Execute.scala 117:10]
  assign _GEN_1962 = 6'h28 == _T_234 ? welem[40] : _GEN_1961; // @[Execute.scala 117:10]
  assign _GEN_1963 = 6'h29 == _T_234 ? welem[41] : _GEN_1962; // @[Execute.scala 117:10]
  assign _GEN_1964 = 6'h2a == _T_234 ? welem[42] : _GEN_1963; // @[Execute.scala 117:10]
  assign _GEN_1965 = 6'h2b == _T_234 ? welem[43] : _GEN_1964; // @[Execute.scala 117:10]
  assign _GEN_1966 = 6'h2c == _T_234 ? welem[44] : _GEN_1965; // @[Execute.scala 117:10]
  assign _GEN_1967 = 6'h2d == _T_234 ? welem[45] : _GEN_1966; // @[Execute.scala 117:10]
  assign _GEN_1968 = 6'h2e == _T_234 ? welem[46] : _GEN_1967; // @[Execute.scala 117:10]
  assign _GEN_1969 = 6'h2f == _T_234 ? welem[47] : _GEN_1968; // @[Execute.scala 117:10]
  assign _GEN_1970 = 6'h30 == _T_234 ? welem[48] : _GEN_1969; // @[Execute.scala 117:10]
  assign _GEN_1971 = 6'h31 == _T_234 ? welem[49] : _GEN_1970; // @[Execute.scala 117:10]
  assign _GEN_1972 = 6'h32 == _T_234 ? welem[50] : _GEN_1971; // @[Execute.scala 117:10]
  assign _GEN_1973 = 6'h33 == _T_234 ? welem[51] : _GEN_1972; // @[Execute.scala 117:10]
  assign _GEN_1974 = 6'h34 == _T_234 ? welem[52] : _GEN_1973; // @[Execute.scala 117:10]
  assign _GEN_1975 = 6'h35 == _T_234 ? welem[53] : _GEN_1974; // @[Execute.scala 117:10]
  assign _GEN_1976 = 6'h36 == _T_234 ? welem[54] : _GEN_1975; // @[Execute.scala 117:10]
  assign _GEN_1977 = 6'h37 == _T_234 ? welem[55] : _GEN_1976; // @[Execute.scala 117:10]
  assign _GEN_1978 = 6'h38 == _T_234 ? welem[56] : _GEN_1977; // @[Execute.scala 117:10]
  assign _GEN_1979 = 6'h39 == _T_234 ? welem[57] : _GEN_1978; // @[Execute.scala 117:10]
  assign _GEN_1980 = 6'h3a == _T_234 ? welem[58] : _GEN_1979; // @[Execute.scala 117:10]
  assign _GEN_1981 = 6'h3b == _T_234 ? welem[59] : _GEN_1980; // @[Execute.scala 117:10]
  assign _GEN_1982 = 6'h3c == _T_234 ? welem[60] : _GEN_1981; // @[Execute.scala 117:10]
  assign _GEN_1983 = 6'h3d == _T_234 ? welem[61] : _GEN_1982; // @[Execute.scala 117:10]
  assign _GEN_1984 = 6'h3e == _T_234 ? welem[62] : _GEN_1983; // @[Execute.scala 117:10]
  assign _GEN_1985 = 6'h3f == _T_234 ? welem[63] : _GEN_1984; // @[Execute.scala 117:10]
  assign _GEN_1987 = 6'h1 == _T_238 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_1988 = 6'h2 == _T_238 ? welem[2] : _GEN_1987; // @[Execute.scala 117:10]
  assign _GEN_1989 = 6'h3 == _T_238 ? welem[3] : _GEN_1988; // @[Execute.scala 117:10]
  assign _GEN_1990 = 6'h4 == _T_238 ? welem[4] : _GEN_1989; // @[Execute.scala 117:10]
  assign _GEN_1991 = 6'h5 == _T_238 ? welem[5] : _GEN_1990; // @[Execute.scala 117:10]
  assign _GEN_1992 = 6'h6 == _T_238 ? welem[6] : _GEN_1991; // @[Execute.scala 117:10]
  assign _GEN_1993 = 6'h7 == _T_238 ? welem[7] : _GEN_1992; // @[Execute.scala 117:10]
  assign _GEN_1994 = 6'h8 == _T_238 ? welem[8] : _GEN_1993; // @[Execute.scala 117:10]
  assign _GEN_1995 = 6'h9 == _T_238 ? welem[9] : _GEN_1994; // @[Execute.scala 117:10]
  assign _GEN_1996 = 6'ha == _T_238 ? welem[10] : _GEN_1995; // @[Execute.scala 117:10]
  assign _GEN_1997 = 6'hb == _T_238 ? welem[11] : _GEN_1996; // @[Execute.scala 117:10]
  assign _GEN_1998 = 6'hc == _T_238 ? welem[12] : _GEN_1997; // @[Execute.scala 117:10]
  assign _GEN_1999 = 6'hd == _T_238 ? welem[13] : _GEN_1998; // @[Execute.scala 117:10]
  assign _GEN_2000 = 6'he == _T_238 ? welem[14] : _GEN_1999; // @[Execute.scala 117:10]
  assign _GEN_2001 = 6'hf == _T_238 ? welem[15] : _GEN_2000; // @[Execute.scala 117:10]
  assign _GEN_2002 = 6'h10 == _T_238 ? welem[16] : _GEN_2001; // @[Execute.scala 117:10]
  assign _GEN_2003 = 6'h11 == _T_238 ? welem[17] : _GEN_2002; // @[Execute.scala 117:10]
  assign _GEN_2004 = 6'h12 == _T_238 ? welem[18] : _GEN_2003; // @[Execute.scala 117:10]
  assign _GEN_2005 = 6'h13 == _T_238 ? welem[19] : _GEN_2004; // @[Execute.scala 117:10]
  assign _GEN_2006 = 6'h14 == _T_238 ? welem[20] : _GEN_2005; // @[Execute.scala 117:10]
  assign _GEN_2007 = 6'h15 == _T_238 ? welem[21] : _GEN_2006; // @[Execute.scala 117:10]
  assign _GEN_2008 = 6'h16 == _T_238 ? welem[22] : _GEN_2007; // @[Execute.scala 117:10]
  assign _GEN_2009 = 6'h17 == _T_238 ? welem[23] : _GEN_2008; // @[Execute.scala 117:10]
  assign _GEN_2010 = 6'h18 == _T_238 ? welem[24] : _GEN_2009; // @[Execute.scala 117:10]
  assign _GEN_2011 = 6'h19 == _T_238 ? welem[25] : _GEN_2010; // @[Execute.scala 117:10]
  assign _GEN_2012 = 6'h1a == _T_238 ? welem[26] : _GEN_2011; // @[Execute.scala 117:10]
  assign _GEN_2013 = 6'h1b == _T_238 ? welem[27] : _GEN_2012; // @[Execute.scala 117:10]
  assign _GEN_2014 = 6'h1c == _T_238 ? welem[28] : _GEN_2013; // @[Execute.scala 117:10]
  assign _GEN_2015 = 6'h1d == _T_238 ? welem[29] : _GEN_2014; // @[Execute.scala 117:10]
  assign _GEN_2016 = 6'h1e == _T_238 ? welem[30] : _GEN_2015; // @[Execute.scala 117:10]
  assign _GEN_2017 = 6'h1f == _T_238 ? welem[31] : _GEN_2016; // @[Execute.scala 117:10]
  assign _GEN_2018 = 6'h20 == _T_238 ? welem[32] : _GEN_2017; // @[Execute.scala 117:10]
  assign _GEN_2019 = 6'h21 == _T_238 ? welem[33] : _GEN_2018; // @[Execute.scala 117:10]
  assign _GEN_2020 = 6'h22 == _T_238 ? welem[34] : _GEN_2019; // @[Execute.scala 117:10]
  assign _GEN_2021 = 6'h23 == _T_238 ? welem[35] : _GEN_2020; // @[Execute.scala 117:10]
  assign _GEN_2022 = 6'h24 == _T_238 ? welem[36] : _GEN_2021; // @[Execute.scala 117:10]
  assign _GEN_2023 = 6'h25 == _T_238 ? welem[37] : _GEN_2022; // @[Execute.scala 117:10]
  assign _GEN_2024 = 6'h26 == _T_238 ? welem[38] : _GEN_2023; // @[Execute.scala 117:10]
  assign _GEN_2025 = 6'h27 == _T_238 ? welem[39] : _GEN_2024; // @[Execute.scala 117:10]
  assign _GEN_2026 = 6'h28 == _T_238 ? welem[40] : _GEN_2025; // @[Execute.scala 117:10]
  assign _GEN_2027 = 6'h29 == _T_238 ? welem[41] : _GEN_2026; // @[Execute.scala 117:10]
  assign _GEN_2028 = 6'h2a == _T_238 ? welem[42] : _GEN_2027; // @[Execute.scala 117:10]
  assign _GEN_2029 = 6'h2b == _T_238 ? welem[43] : _GEN_2028; // @[Execute.scala 117:10]
  assign _GEN_2030 = 6'h2c == _T_238 ? welem[44] : _GEN_2029; // @[Execute.scala 117:10]
  assign _GEN_2031 = 6'h2d == _T_238 ? welem[45] : _GEN_2030; // @[Execute.scala 117:10]
  assign _GEN_2032 = 6'h2e == _T_238 ? welem[46] : _GEN_2031; // @[Execute.scala 117:10]
  assign _GEN_2033 = 6'h2f == _T_238 ? welem[47] : _GEN_2032; // @[Execute.scala 117:10]
  assign _GEN_2034 = 6'h30 == _T_238 ? welem[48] : _GEN_2033; // @[Execute.scala 117:10]
  assign _GEN_2035 = 6'h31 == _T_238 ? welem[49] : _GEN_2034; // @[Execute.scala 117:10]
  assign _GEN_2036 = 6'h32 == _T_238 ? welem[50] : _GEN_2035; // @[Execute.scala 117:10]
  assign _GEN_2037 = 6'h33 == _T_238 ? welem[51] : _GEN_2036; // @[Execute.scala 117:10]
  assign _GEN_2038 = 6'h34 == _T_238 ? welem[52] : _GEN_2037; // @[Execute.scala 117:10]
  assign _GEN_2039 = 6'h35 == _T_238 ? welem[53] : _GEN_2038; // @[Execute.scala 117:10]
  assign _GEN_2040 = 6'h36 == _T_238 ? welem[54] : _GEN_2039; // @[Execute.scala 117:10]
  assign _GEN_2041 = 6'h37 == _T_238 ? welem[55] : _GEN_2040; // @[Execute.scala 117:10]
  assign _GEN_2042 = 6'h38 == _T_238 ? welem[56] : _GEN_2041; // @[Execute.scala 117:10]
  assign _GEN_2043 = 6'h39 == _T_238 ? welem[57] : _GEN_2042; // @[Execute.scala 117:10]
  assign _GEN_2044 = 6'h3a == _T_238 ? welem[58] : _GEN_2043; // @[Execute.scala 117:10]
  assign _GEN_2045 = 6'h3b == _T_238 ? welem[59] : _GEN_2044; // @[Execute.scala 117:10]
  assign _GEN_2046 = 6'h3c == _T_238 ? welem[60] : _GEN_2045; // @[Execute.scala 117:10]
  assign _GEN_2047 = 6'h3d == _T_238 ? welem[61] : _GEN_2046; // @[Execute.scala 117:10]
  assign _GEN_2048 = 6'h3e == _T_238 ? welem[62] : _GEN_2047; // @[Execute.scala 117:10]
  assign _GEN_2049 = 6'h3f == _T_238 ? welem[63] : _GEN_2048; // @[Execute.scala 117:10]
  assign _T_241 = _T_232 ? _GEN_1985 : _GEN_2049; // @[Execute.scala 117:10]
  assign _T_242 = r < 6'h31; // @[Execute.scala 117:15]
  assign _T_244 = r - 6'h31; // @[Execute.scala 117:37]
  assign _T_248 = 6'hf + r; // @[Execute.scala 117:60]
  assign _GEN_2051 = 6'h1 == _T_244 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2052 = 6'h2 == _T_244 ? welem[2] : _GEN_2051; // @[Execute.scala 117:10]
  assign _GEN_2053 = 6'h3 == _T_244 ? welem[3] : _GEN_2052; // @[Execute.scala 117:10]
  assign _GEN_2054 = 6'h4 == _T_244 ? welem[4] : _GEN_2053; // @[Execute.scala 117:10]
  assign _GEN_2055 = 6'h5 == _T_244 ? welem[5] : _GEN_2054; // @[Execute.scala 117:10]
  assign _GEN_2056 = 6'h6 == _T_244 ? welem[6] : _GEN_2055; // @[Execute.scala 117:10]
  assign _GEN_2057 = 6'h7 == _T_244 ? welem[7] : _GEN_2056; // @[Execute.scala 117:10]
  assign _GEN_2058 = 6'h8 == _T_244 ? welem[8] : _GEN_2057; // @[Execute.scala 117:10]
  assign _GEN_2059 = 6'h9 == _T_244 ? welem[9] : _GEN_2058; // @[Execute.scala 117:10]
  assign _GEN_2060 = 6'ha == _T_244 ? welem[10] : _GEN_2059; // @[Execute.scala 117:10]
  assign _GEN_2061 = 6'hb == _T_244 ? welem[11] : _GEN_2060; // @[Execute.scala 117:10]
  assign _GEN_2062 = 6'hc == _T_244 ? welem[12] : _GEN_2061; // @[Execute.scala 117:10]
  assign _GEN_2063 = 6'hd == _T_244 ? welem[13] : _GEN_2062; // @[Execute.scala 117:10]
  assign _GEN_2064 = 6'he == _T_244 ? welem[14] : _GEN_2063; // @[Execute.scala 117:10]
  assign _GEN_2065 = 6'hf == _T_244 ? welem[15] : _GEN_2064; // @[Execute.scala 117:10]
  assign _GEN_2066 = 6'h10 == _T_244 ? welem[16] : _GEN_2065; // @[Execute.scala 117:10]
  assign _GEN_2067 = 6'h11 == _T_244 ? welem[17] : _GEN_2066; // @[Execute.scala 117:10]
  assign _GEN_2068 = 6'h12 == _T_244 ? welem[18] : _GEN_2067; // @[Execute.scala 117:10]
  assign _GEN_2069 = 6'h13 == _T_244 ? welem[19] : _GEN_2068; // @[Execute.scala 117:10]
  assign _GEN_2070 = 6'h14 == _T_244 ? welem[20] : _GEN_2069; // @[Execute.scala 117:10]
  assign _GEN_2071 = 6'h15 == _T_244 ? welem[21] : _GEN_2070; // @[Execute.scala 117:10]
  assign _GEN_2072 = 6'h16 == _T_244 ? welem[22] : _GEN_2071; // @[Execute.scala 117:10]
  assign _GEN_2073 = 6'h17 == _T_244 ? welem[23] : _GEN_2072; // @[Execute.scala 117:10]
  assign _GEN_2074 = 6'h18 == _T_244 ? welem[24] : _GEN_2073; // @[Execute.scala 117:10]
  assign _GEN_2075 = 6'h19 == _T_244 ? welem[25] : _GEN_2074; // @[Execute.scala 117:10]
  assign _GEN_2076 = 6'h1a == _T_244 ? welem[26] : _GEN_2075; // @[Execute.scala 117:10]
  assign _GEN_2077 = 6'h1b == _T_244 ? welem[27] : _GEN_2076; // @[Execute.scala 117:10]
  assign _GEN_2078 = 6'h1c == _T_244 ? welem[28] : _GEN_2077; // @[Execute.scala 117:10]
  assign _GEN_2079 = 6'h1d == _T_244 ? welem[29] : _GEN_2078; // @[Execute.scala 117:10]
  assign _GEN_2080 = 6'h1e == _T_244 ? welem[30] : _GEN_2079; // @[Execute.scala 117:10]
  assign _GEN_2081 = 6'h1f == _T_244 ? welem[31] : _GEN_2080; // @[Execute.scala 117:10]
  assign _GEN_2082 = 6'h20 == _T_244 ? welem[32] : _GEN_2081; // @[Execute.scala 117:10]
  assign _GEN_2083 = 6'h21 == _T_244 ? welem[33] : _GEN_2082; // @[Execute.scala 117:10]
  assign _GEN_2084 = 6'h22 == _T_244 ? welem[34] : _GEN_2083; // @[Execute.scala 117:10]
  assign _GEN_2085 = 6'h23 == _T_244 ? welem[35] : _GEN_2084; // @[Execute.scala 117:10]
  assign _GEN_2086 = 6'h24 == _T_244 ? welem[36] : _GEN_2085; // @[Execute.scala 117:10]
  assign _GEN_2087 = 6'h25 == _T_244 ? welem[37] : _GEN_2086; // @[Execute.scala 117:10]
  assign _GEN_2088 = 6'h26 == _T_244 ? welem[38] : _GEN_2087; // @[Execute.scala 117:10]
  assign _GEN_2089 = 6'h27 == _T_244 ? welem[39] : _GEN_2088; // @[Execute.scala 117:10]
  assign _GEN_2090 = 6'h28 == _T_244 ? welem[40] : _GEN_2089; // @[Execute.scala 117:10]
  assign _GEN_2091 = 6'h29 == _T_244 ? welem[41] : _GEN_2090; // @[Execute.scala 117:10]
  assign _GEN_2092 = 6'h2a == _T_244 ? welem[42] : _GEN_2091; // @[Execute.scala 117:10]
  assign _GEN_2093 = 6'h2b == _T_244 ? welem[43] : _GEN_2092; // @[Execute.scala 117:10]
  assign _GEN_2094 = 6'h2c == _T_244 ? welem[44] : _GEN_2093; // @[Execute.scala 117:10]
  assign _GEN_2095 = 6'h2d == _T_244 ? welem[45] : _GEN_2094; // @[Execute.scala 117:10]
  assign _GEN_2096 = 6'h2e == _T_244 ? welem[46] : _GEN_2095; // @[Execute.scala 117:10]
  assign _GEN_2097 = 6'h2f == _T_244 ? welem[47] : _GEN_2096; // @[Execute.scala 117:10]
  assign _GEN_2098 = 6'h30 == _T_244 ? welem[48] : _GEN_2097; // @[Execute.scala 117:10]
  assign _GEN_2099 = 6'h31 == _T_244 ? welem[49] : _GEN_2098; // @[Execute.scala 117:10]
  assign _GEN_2100 = 6'h32 == _T_244 ? welem[50] : _GEN_2099; // @[Execute.scala 117:10]
  assign _GEN_2101 = 6'h33 == _T_244 ? welem[51] : _GEN_2100; // @[Execute.scala 117:10]
  assign _GEN_2102 = 6'h34 == _T_244 ? welem[52] : _GEN_2101; // @[Execute.scala 117:10]
  assign _GEN_2103 = 6'h35 == _T_244 ? welem[53] : _GEN_2102; // @[Execute.scala 117:10]
  assign _GEN_2104 = 6'h36 == _T_244 ? welem[54] : _GEN_2103; // @[Execute.scala 117:10]
  assign _GEN_2105 = 6'h37 == _T_244 ? welem[55] : _GEN_2104; // @[Execute.scala 117:10]
  assign _GEN_2106 = 6'h38 == _T_244 ? welem[56] : _GEN_2105; // @[Execute.scala 117:10]
  assign _GEN_2107 = 6'h39 == _T_244 ? welem[57] : _GEN_2106; // @[Execute.scala 117:10]
  assign _GEN_2108 = 6'h3a == _T_244 ? welem[58] : _GEN_2107; // @[Execute.scala 117:10]
  assign _GEN_2109 = 6'h3b == _T_244 ? welem[59] : _GEN_2108; // @[Execute.scala 117:10]
  assign _GEN_2110 = 6'h3c == _T_244 ? welem[60] : _GEN_2109; // @[Execute.scala 117:10]
  assign _GEN_2111 = 6'h3d == _T_244 ? welem[61] : _GEN_2110; // @[Execute.scala 117:10]
  assign _GEN_2112 = 6'h3e == _T_244 ? welem[62] : _GEN_2111; // @[Execute.scala 117:10]
  assign _GEN_2113 = 6'h3f == _T_244 ? welem[63] : _GEN_2112; // @[Execute.scala 117:10]
  assign _GEN_2115 = 6'h1 == _T_248 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2116 = 6'h2 == _T_248 ? welem[2] : _GEN_2115; // @[Execute.scala 117:10]
  assign _GEN_2117 = 6'h3 == _T_248 ? welem[3] : _GEN_2116; // @[Execute.scala 117:10]
  assign _GEN_2118 = 6'h4 == _T_248 ? welem[4] : _GEN_2117; // @[Execute.scala 117:10]
  assign _GEN_2119 = 6'h5 == _T_248 ? welem[5] : _GEN_2118; // @[Execute.scala 117:10]
  assign _GEN_2120 = 6'h6 == _T_248 ? welem[6] : _GEN_2119; // @[Execute.scala 117:10]
  assign _GEN_2121 = 6'h7 == _T_248 ? welem[7] : _GEN_2120; // @[Execute.scala 117:10]
  assign _GEN_2122 = 6'h8 == _T_248 ? welem[8] : _GEN_2121; // @[Execute.scala 117:10]
  assign _GEN_2123 = 6'h9 == _T_248 ? welem[9] : _GEN_2122; // @[Execute.scala 117:10]
  assign _GEN_2124 = 6'ha == _T_248 ? welem[10] : _GEN_2123; // @[Execute.scala 117:10]
  assign _GEN_2125 = 6'hb == _T_248 ? welem[11] : _GEN_2124; // @[Execute.scala 117:10]
  assign _GEN_2126 = 6'hc == _T_248 ? welem[12] : _GEN_2125; // @[Execute.scala 117:10]
  assign _GEN_2127 = 6'hd == _T_248 ? welem[13] : _GEN_2126; // @[Execute.scala 117:10]
  assign _GEN_2128 = 6'he == _T_248 ? welem[14] : _GEN_2127; // @[Execute.scala 117:10]
  assign _GEN_2129 = 6'hf == _T_248 ? welem[15] : _GEN_2128; // @[Execute.scala 117:10]
  assign _GEN_2130 = 6'h10 == _T_248 ? welem[16] : _GEN_2129; // @[Execute.scala 117:10]
  assign _GEN_2131 = 6'h11 == _T_248 ? welem[17] : _GEN_2130; // @[Execute.scala 117:10]
  assign _GEN_2132 = 6'h12 == _T_248 ? welem[18] : _GEN_2131; // @[Execute.scala 117:10]
  assign _GEN_2133 = 6'h13 == _T_248 ? welem[19] : _GEN_2132; // @[Execute.scala 117:10]
  assign _GEN_2134 = 6'h14 == _T_248 ? welem[20] : _GEN_2133; // @[Execute.scala 117:10]
  assign _GEN_2135 = 6'h15 == _T_248 ? welem[21] : _GEN_2134; // @[Execute.scala 117:10]
  assign _GEN_2136 = 6'h16 == _T_248 ? welem[22] : _GEN_2135; // @[Execute.scala 117:10]
  assign _GEN_2137 = 6'h17 == _T_248 ? welem[23] : _GEN_2136; // @[Execute.scala 117:10]
  assign _GEN_2138 = 6'h18 == _T_248 ? welem[24] : _GEN_2137; // @[Execute.scala 117:10]
  assign _GEN_2139 = 6'h19 == _T_248 ? welem[25] : _GEN_2138; // @[Execute.scala 117:10]
  assign _GEN_2140 = 6'h1a == _T_248 ? welem[26] : _GEN_2139; // @[Execute.scala 117:10]
  assign _GEN_2141 = 6'h1b == _T_248 ? welem[27] : _GEN_2140; // @[Execute.scala 117:10]
  assign _GEN_2142 = 6'h1c == _T_248 ? welem[28] : _GEN_2141; // @[Execute.scala 117:10]
  assign _GEN_2143 = 6'h1d == _T_248 ? welem[29] : _GEN_2142; // @[Execute.scala 117:10]
  assign _GEN_2144 = 6'h1e == _T_248 ? welem[30] : _GEN_2143; // @[Execute.scala 117:10]
  assign _GEN_2145 = 6'h1f == _T_248 ? welem[31] : _GEN_2144; // @[Execute.scala 117:10]
  assign _GEN_2146 = 6'h20 == _T_248 ? welem[32] : _GEN_2145; // @[Execute.scala 117:10]
  assign _GEN_2147 = 6'h21 == _T_248 ? welem[33] : _GEN_2146; // @[Execute.scala 117:10]
  assign _GEN_2148 = 6'h22 == _T_248 ? welem[34] : _GEN_2147; // @[Execute.scala 117:10]
  assign _GEN_2149 = 6'h23 == _T_248 ? welem[35] : _GEN_2148; // @[Execute.scala 117:10]
  assign _GEN_2150 = 6'h24 == _T_248 ? welem[36] : _GEN_2149; // @[Execute.scala 117:10]
  assign _GEN_2151 = 6'h25 == _T_248 ? welem[37] : _GEN_2150; // @[Execute.scala 117:10]
  assign _GEN_2152 = 6'h26 == _T_248 ? welem[38] : _GEN_2151; // @[Execute.scala 117:10]
  assign _GEN_2153 = 6'h27 == _T_248 ? welem[39] : _GEN_2152; // @[Execute.scala 117:10]
  assign _GEN_2154 = 6'h28 == _T_248 ? welem[40] : _GEN_2153; // @[Execute.scala 117:10]
  assign _GEN_2155 = 6'h29 == _T_248 ? welem[41] : _GEN_2154; // @[Execute.scala 117:10]
  assign _GEN_2156 = 6'h2a == _T_248 ? welem[42] : _GEN_2155; // @[Execute.scala 117:10]
  assign _GEN_2157 = 6'h2b == _T_248 ? welem[43] : _GEN_2156; // @[Execute.scala 117:10]
  assign _GEN_2158 = 6'h2c == _T_248 ? welem[44] : _GEN_2157; // @[Execute.scala 117:10]
  assign _GEN_2159 = 6'h2d == _T_248 ? welem[45] : _GEN_2158; // @[Execute.scala 117:10]
  assign _GEN_2160 = 6'h2e == _T_248 ? welem[46] : _GEN_2159; // @[Execute.scala 117:10]
  assign _GEN_2161 = 6'h2f == _T_248 ? welem[47] : _GEN_2160; // @[Execute.scala 117:10]
  assign _GEN_2162 = 6'h30 == _T_248 ? welem[48] : _GEN_2161; // @[Execute.scala 117:10]
  assign _GEN_2163 = 6'h31 == _T_248 ? welem[49] : _GEN_2162; // @[Execute.scala 117:10]
  assign _GEN_2164 = 6'h32 == _T_248 ? welem[50] : _GEN_2163; // @[Execute.scala 117:10]
  assign _GEN_2165 = 6'h33 == _T_248 ? welem[51] : _GEN_2164; // @[Execute.scala 117:10]
  assign _GEN_2166 = 6'h34 == _T_248 ? welem[52] : _GEN_2165; // @[Execute.scala 117:10]
  assign _GEN_2167 = 6'h35 == _T_248 ? welem[53] : _GEN_2166; // @[Execute.scala 117:10]
  assign _GEN_2168 = 6'h36 == _T_248 ? welem[54] : _GEN_2167; // @[Execute.scala 117:10]
  assign _GEN_2169 = 6'h37 == _T_248 ? welem[55] : _GEN_2168; // @[Execute.scala 117:10]
  assign _GEN_2170 = 6'h38 == _T_248 ? welem[56] : _GEN_2169; // @[Execute.scala 117:10]
  assign _GEN_2171 = 6'h39 == _T_248 ? welem[57] : _GEN_2170; // @[Execute.scala 117:10]
  assign _GEN_2172 = 6'h3a == _T_248 ? welem[58] : _GEN_2171; // @[Execute.scala 117:10]
  assign _GEN_2173 = 6'h3b == _T_248 ? welem[59] : _GEN_2172; // @[Execute.scala 117:10]
  assign _GEN_2174 = 6'h3c == _T_248 ? welem[60] : _GEN_2173; // @[Execute.scala 117:10]
  assign _GEN_2175 = 6'h3d == _T_248 ? welem[61] : _GEN_2174; // @[Execute.scala 117:10]
  assign _GEN_2176 = 6'h3e == _T_248 ? welem[62] : _GEN_2175; // @[Execute.scala 117:10]
  assign _GEN_2177 = 6'h3f == _T_248 ? welem[63] : _GEN_2176; // @[Execute.scala 117:10]
  assign _T_251 = _T_242 ? _GEN_2113 : _GEN_2177; // @[Execute.scala 117:10]
  assign _T_252 = r < 6'h30; // @[Execute.scala 117:15]
  assign _T_254 = r - 6'h30; // @[Execute.scala 117:37]
  assign _T_258 = 6'h10 + r; // @[Execute.scala 117:60]
  assign _GEN_2179 = 6'h1 == _T_254 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2180 = 6'h2 == _T_254 ? welem[2] : _GEN_2179; // @[Execute.scala 117:10]
  assign _GEN_2181 = 6'h3 == _T_254 ? welem[3] : _GEN_2180; // @[Execute.scala 117:10]
  assign _GEN_2182 = 6'h4 == _T_254 ? welem[4] : _GEN_2181; // @[Execute.scala 117:10]
  assign _GEN_2183 = 6'h5 == _T_254 ? welem[5] : _GEN_2182; // @[Execute.scala 117:10]
  assign _GEN_2184 = 6'h6 == _T_254 ? welem[6] : _GEN_2183; // @[Execute.scala 117:10]
  assign _GEN_2185 = 6'h7 == _T_254 ? welem[7] : _GEN_2184; // @[Execute.scala 117:10]
  assign _GEN_2186 = 6'h8 == _T_254 ? welem[8] : _GEN_2185; // @[Execute.scala 117:10]
  assign _GEN_2187 = 6'h9 == _T_254 ? welem[9] : _GEN_2186; // @[Execute.scala 117:10]
  assign _GEN_2188 = 6'ha == _T_254 ? welem[10] : _GEN_2187; // @[Execute.scala 117:10]
  assign _GEN_2189 = 6'hb == _T_254 ? welem[11] : _GEN_2188; // @[Execute.scala 117:10]
  assign _GEN_2190 = 6'hc == _T_254 ? welem[12] : _GEN_2189; // @[Execute.scala 117:10]
  assign _GEN_2191 = 6'hd == _T_254 ? welem[13] : _GEN_2190; // @[Execute.scala 117:10]
  assign _GEN_2192 = 6'he == _T_254 ? welem[14] : _GEN_2191; // @[Execute.scala 117:10]
  assign _GEN_2193 = 6'hf == _T_254 ? welem[15] : _GEN_2192; // @[Execute.scala 117:10]
  assign _GEN_2194 = 6'h10 == _T_254 ? welem[16] : _GEN_2193; // @[Execute.scala 117:10]
  assign _GEN_2195 = 6'h11 == _T_254 ? welem[17] : _GEN_2194; // @[Execute.scala 117:10]
  assign _GEN_2196 = 6'h12 == _T_254 ? welem[18] : _GEN_2195; // @[Execute.scala 117:10]
  assign _GEN_2197 = 6'h13 == _T_254 ? welem[19] : _GEN_2196; // @[Execute.scala 117:10]
  assign _GEN_2198 = 6'h14 == _T_254 ? welem[20] : _GEN_2197; // @[Execute.scala 117:10]
  assign _GEN_2199 = 6'h15 == _T_254 ? welem[21] : _GEN_2198; // @[Execute.scala 117:10]
  assign _GEN_2200 = 6'h16 == _T_254 ? welem[22] : _GEN_2199; // @[Execute.scala 117:10]
  assign _GEN_2201 = 6'h17 == _T_254 ? welem[23] : _GEN_2200; // @[Execute.scala 117:10]
  assign _GEN_2202 = 6'h18 == _T_254 ? welem[24] : _GEN_2201; // @[Execute.scala 117:10]
  assign _GEN_2203 = 6'h19 == _T_254 ? welem[25] : _GEN_2202; // @[Execute.scala 117:10]
  assign _GEN_2204 = 6'h1a == _T_254 ? welem[26] : _GEN_2203; // @[Execute.scala 117:10]
  assign _GEN_2205 = 6'h1b == _T_254 ? welem[27] : _GEN_2204; // @[Execute.scala 117:10]
  assign _GEN_2206 = 6'h1c == _T_254 ? welem[28] : _GEN_2205; // @[Execute.scala 117:10]
  assign _GEN_2207 = 6'h1d == _T_254 ? welem[29] : _GEN_2206; // @[Execute.scala 117:10]
  assign _GEN_2208 = 6'h1e == _T_254 ? welem[30] : _GEN_2207; // @[Execute.scala 117:10]
  assign _GEN_2209 = 6'h1f == _T_254 ? welem[31] : _GEN_2208; // @[Execute.scala 117:10]
  assign _GEN_2210 = 6'h20 == _T_254 ? welem[32] : _GEN_2209; // @[Execute.scala 117:10]
  assign _GEN_2211 = 6'h21 == _T_254 ? welem[33] : _GEN_2210; // @[Execute.scala 117:10]
  assign _GEN_2212 = 6'h22 == _T_254 ? welem[34] : _GEN_2211; // @[Execute.scala 117:10]
  assign _GEN_2213 = 6'h23 == _T_254 ? welem[35] : _GEN_2212; // @[Execute.scala 117:10]
  assign _GEN_2214 = 6'h24 == _T_254 ? welem[36] : _GEN_2213; // @[Execute.scala 117:10]
  assign _GEN_2215 = 6'h25 == _T_254 ? welem[37] : _GEN_2214; // @[Execute.scala 117:10]
  assign _GEN_2216 = 6'h26 == _T_254 ? welem[38] : _GEN_2215; // @[Execute.scala 117:10]
  assign _GEN_2217 = 6'h27 == _T_254 ? welem[39] : _GEN_2216; // @[Execute.scala 117:10]
  assign _GEN_2218 = 6'h28 == _T_254 ? welem[40] : _GEN_2217; // @[Execute.scala 117:10]
  assign _GEN_2219 = 6'h29 == _T_254 ? welem[41] : _GEN_2218; // @[Execute.scala 117:10]
  assign _GEN_2220 = 6'h2a == _T_254 ? welem[42] : _GEN_2219; // @[Execute.scala 117:10]
  assign _GEN_2221 = 6'h2b == _T_254 ? welem[43] : _GEN_2220; // @[Execute.scala 117:10]
  assign _GEN_2222 = 6'h2c == _T_254 ? welem[44] : _GEN_2221; // @[Execute.scala 117:10]
  assign _GEN_2223 = 6'h2d == _T_254 ? welem[45] : _GEN_2222; // @[Execute.scala 117:10]
  assign _GEN_2224 = 6'h2e == _T_254 ? welem[46] : _GEN_2223; // @[Execute.scala 117:10]
  assign _GEN_2225 = 6'h2f == _T_254 ? welem[47] : _GEN_2224; // @[Execute.scala 117:10]
  assign _GEN_2226 = 6'h30 == _T_254 ? welem[48] : _GEN_2225; // @[Execute.scala 117:10]
  assign _GEN_2227 = 6'h31 == _T_254 ? welem[49] : _GEN_2226; // @[Execute.scala 117:10]
  assign _GEN_2228 = 6'h32 == _T_254 ? welem[50] : _GEN_2227; // @[Execute.scala 117:10]
  assign _GEN_2229 = 6'h33 == _T_254 ? welem[51] : _GEN_2228; // @[Execute.scala 117:10]
  assign _GEN_2230 = 6'h34 == _T_254 ? welem[52] : _GEN_2229; // @[Execute.scala 117:10]
  assign _GEN_2231 = 6'h35 == _T_254 ? welem[53] : _GEN_2230; // @[Execute.scala 117:10]
  assign _GEN_2232 = 6'h36 == _T_254 ? welem[54] : _GEN_2231; // @[Execute.scala 117:10]
  assign _GEN_2233 = 6'h37 == _T_254 ? welem[55] : _GEN_2232; // @[Execute.scala 117:10]
  assign _GEN_2234 = 6'h38 == _T_254 ? welem[56] : _GEN_2233; // @[Execute.scala 117:10]
  assign _GEN_2235 = 6'h39 == _T_254 ? welem[57] : _GEN_2234; // @[Execute.scala 117:10]
  assign _GEN_2236 = 6'h3a == _T_254 ? welem[58] : _GEN_2235; // @[Execute.scala 117:10]
  assign _GEN_2237 = 6'h3b == _T_254 ? welem[59] : _GEN_2236; // @[Execute.scala 117:10]
  assign _GEN_2238 = 6'h3c == _T_254 ? welem[60] : _GEN_2237; // @[Execute.scala 117:10]
  assign _GEN_2239 = 6'h3d == _T_254 ? welem[61] : _GEN_2238; // @[Execute.scala 117:10]
  assign _GEN_2240 = 6'h3e == _T_254 ? welem[62] : _GEN_2239; // @[Execute.scala 117:10]
  assign _GEN_2241 = 6'h3f == _T_254 ? welem[63] : _GEN_2240; // @[Execute.scala 117:10]
  assign _GEN_2243 = 6'h1 == _T_258 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2244 = 6'h2 == _T_258 ? welem[2] : _GEN_2243; // @[Execute.scala 117:10]
  assign _GEN_2245 = 6'h3 == _T_258 ? welem[3] : _GEN_2244; // @[Execute.scala 117:10]
  assign _GEN_2246 = 6'h4 == _T_258 ? welem[4] : _GEN_2245; // @[Execute.scala 117:10]
  assign _GEN_2247 = 6'h5 == _T_258 ? welem[5] : _GEN_2246; // @[Execute.scala 117:10]
  assign _GEN_2248 = 6'h6 == _T_258 ? welem[6] : _GEN_2247; // @[Execute.scala 117:10]
  assign _GEN_2249 = 6'h7 == _T_258 ? welem[7] : _GEN_2248; // @[Execute.scala 117:10]
  assign _GEN_2250 = 6'h8 == _T_258 ? welem[8] : _GEN_2249; // @[Execute.scala 117:10]
  assign _GEN_2251 = 6'h9 == _T_258 ? welem[9] : _GEN_2250; // @[Execute.scala 117:10]
  assign _GEN_2252 = 6'ha == _T_258 ? welem[10] : _GEN_2251; // @[Execute.scala 117:10]
  assign _GEN_2253 = 6'hb == _T_258 ? welem[11] : _GEN_2252; // @[Execute.scala 117:10]
  assign _GEN_2254 = 6'hc == _T_258 ? welem[12] : _GEN_2253; // @[Execute.scala 117:10]
  assign _GEN_2255 = 6'hd == _T_258 ? welem[13] : _GEN_2254; // @[Execute.scala 117:10]
  assign _GEN_2256 = 6'he == _T_258 ? welem[14] : _GEN_2255; // @[Execute.scala 117:10]
  assign _GEN_2257 = 6'hf == _T_258 ? welem[15] : _GEN_2256; // @[Execute.scala 117:10]
  assign _GEN_2258 = 6'h10 == _T_258 ? welem[16] : _GEN_2257; // @[Execute.scala 117:10]
  assign _GEN_2259 = 6'h11 == _T_258 ? welem[17] : _GEN_2258; // @[Execute.scala 117:10]
  assign _GEN_2260 = 6'h12 == _T_258 ? welem[18] : _GEN_2259; // @[Execute.scala 117:10]
  assign _GEN_2261 = 6'h13 == _T_258 ? welem[19] : _GEN_2260; // @[Execute.scala 117:10]
  assign _GEN_2262 = 6'h14 == _T_258 ? welem[20] : _GEN_2261; // @[Execute.scala 117:10]
  assign _GEN_2263 = 6'h15 == _T_258 ? welem[21] : _GEN_2262; // @[Execute.scala 117:10]
  assign _GEN_2264 = 6'h16 == _T_258 ? welem[22] : _GEN_2263; // @[Execute.scala 117:10]
  assign _GEN_2265 = 6'h17 == _T_258 ? welem[23] : _GEN_2264; // @[Execute.scala 117:10]
  assign _GEN_2266 = 6'h18 == _T_258 ? welem[24] : _GEN_2265; // @[Execute.scala 117:10]
  assign _GEN_2267 = 6'h19 == _T_258 ? welem[25] : _GEN_2266; // @[Execute.scala 117:10]
  assign _GEN_2268 = 6'h1a == _T_258 ? welem[26] : _GEN_2267; // @[Execute.scala 117:10]
  assign _GEN_2269 = 6'h1b == _T_258 ? welem[27] : _GEN_2268; // @[Execute.scala 117:10]
  assign _GEN_2270 = 6'h1c == _T_258 ? welem[28] : _GEN_2269; // @[Execute.scala 117:10]
  assign _GEN_2271 = 6'h1d == _T_258 ? welem[29] : _GEN_2270; // @[Execute.scala 117:10]
  assign _GEN_2272 = 6'h1e == _T_258 ? welem[30] : _GEN_2271; // @[Execute.scala 117:10]
  assign _GEN_2273 = 6'h1f == _T_258 ? welem[31] : _GEN_2272; // @[Execute.scala 117:10]
  assign _GEN_2274 = 6'h20 == _T_258 ? welem[32] : _GEN_2273; // @[Execute.scala 117:10]
  assign _GEN_2275 = 6'h21 == _T_258 ? welem[33] : _GEN_2274; // @[Execute.scala 117:10]
  assign _GEN_2276 = 6'h22 == _T_258 ? welem[34] : _GEN_2275; // @[Execute.scala 117:10]
  assign _GEN_2277 = 6'h23 == _T_258 ? welem[35] : _GEN_2276; // @[Execute.scala 117:10]
  assign _GEN_2278 = 6'h24 == _T_258 ? welem[36] : _GEN_2277; // @[Execute.scala 117:10]
  assign _GEN_2279 = 6'h25 == _T_258 ? welem[37] : _GEN_2278; // @[Execute.scala 117:10]
  assign _GEN_2280 = 6'h26 == _T_258 ? welem[38] : _GEN_2279; // @[Execute.scala 117:10]
  assign _GEN_2281 = 6'h27 == _T_258 ? welem[39] : _GEN_2280; // @[Execute.scala 117:10]
  assign _GEN_2282 = 6'h28 == _T_258 ? welem[40] : _GEN_2281; // @[Execute.scala 117:10]
  assign _GEN_2283 = 6'h29 == _T_258 ? welem[41] : _GEN_2282; // @[Execute.scala 117:10]
  assign _GEN_2284 = 6'h2a == _T_258 ? welem[42] : _GEN_2283; // @[Execute.scala 117:10]
  assign _GEN_2285 = 6'h2b == _T_258 ? welem[43] : _GEN_2284; // @[Execute.scala 117:10]
  assign _GEN_2286 = 6'h2c == _T_258 ? welem[44] : _GEN_2285; // @[Execute.scala 117:10]
  assign _GEN_2287 = 6'h2d == _T_258 ? welem[45] : _GEN_2286; // @[Execute.scala 117:10]
  assign _GEN_2288 = 6'h2e == _T_258 ? welem[46] : _GEN_2287; // @[Execute.scala 117:10]
  assign _GEN_2289 = 6'h2f == _T_258 ? welem[47] : _GEN_2288; // @[Execute.scala 117:10]
  assign _GEN_2290 = 6'h30 == _T_258 ? welem[48] : _GEN_2289; // @[Execute.scala 117:10]
  assign _GEN_2291 = 6'h31 == _T_258 ? welem[49] : _GEN_2290; // @[Execute.scala 117:10]
  assign _GEN_2292 = 6'h32 == _T_258 ? welem[50] : _GEN_2291; // @[Execute.scala 117:10]
  assign _GEN_2293 = 6'h33 == _T_258 ? welem[51] : _GEN_2292; // @[Execute.scala 117:10]
  assign _GEN_2294 = 6'h34 == _T_258 ? welem[52] : _GEN_2293; // @[Execute.scala 117:10]
  assign _GEN_2295 = 6'h35 == _T_258 ? welem[53] : _GEN_2294; // @[Execute.scala 117:10]
  assign _GEN_2296 = 6'h36 == _T_258 ? welem[54] : _GEN_2295; // @[Execute.scala 117:10]
  assign _GEN_2297 = 6'h37 == _T_258 ? welem[55] : _GEN_2296; // @[Execute.scala 117:10]
  assign _GEN_2298 = 6'h38 == _T_258 ? welem[56] : _GEN_2297; // @[Execute.scala 117:10]
  assign _GEN_2299 = 6'h39 == _T_258 ? welem[57] : _GEN_2298; // @[Execute.scala 117:10]
  assign _GEN_2300 = 6'h3a == _T_258 ? welem[58] : _GEN_2299; // @[Execute.scala 117:10]
  assign _GEN_2301 = 6'h3b == _T_258 ? welem[59] : _GEN_2300; // @[Execute.scala 117:10]
  assign _GEN_2302 = 6'h3c == _T_258 ? welem[60] : _GEN_2301; // @[Execute.scala 117:10]
  assign _GEN_2303 = 6'h3d == _T_258 ? welem[61] : _GEN_2302; // @[Execute.scala 117:10]
  assign _GEN_2304 = 6'h3e == _T_258 ? welem[62] : _GEN_2303; // @[Execute.scala 117:10]
  assign _GEN_2305 = 6'h3f == _T_258 ? welem[63] : _GEN_2304; // @[Execute.scala 117:10]
  assign _T_261 = _T_252 ? _GEN_2241 : _GEN_2305; // @[Execute.scala 117:10]
  assign _T_262 = r < 6'h2f; // @[Execute.scala 117:15]
  assign _T_264 = r - 6'h2f; // @[Execute.scala 117:37]
  assign _T_268 = 6'h11 + r; // @[Execute.scala 117:60]
  assign _GEN_2307 = 6'h1 == _T_264 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2308 = 6'h2 == _T_264 ? welem[2] : _GEN_2307; // @[Execute.scala 117:10]
  assign _GEN_2309 = 6'h3 == _T_264 ? welem[3] : _GEN_2308; // @[Execute.scala 117:10]
  assign _GEN_2310 = 6'h4 == _T_264 ? welem[4] : _GEN_2309; // @[Execute.scala 117:10]
  assign _GEN_2311 = 6'h5 == _T_264 ? welem[5] : _GEN_2310; // @[Execute.scala 117:10]
  assign _GEN_2312 = 6'h6 == _T_264 ? welem[6] : _GEN_2311; // @[Execute.scala 117:10]
  assign _GEN_2313 = 6'h7 == _T_264 ? welem[7] : _GEN_2312; // @[Execute.scala 117:10]
  assign _GEN_2314 = 6'h8 == _T_264 ? welem[8] : _GEN_2313; // @[Execute.scala 117:10]
  assign _GEN_2315 = 6'h9 == _T_264 ? welem[9] : _GEN_2314; // @[Execute.scala 117:10]
  assign _GEN_2316 = 6'ha == _T_264 ? welem[10] : _GEN_2315; // @[Execute.scala 117:10]
  assign _GEN_2317 = 6'hb == _T_264 ? welem[11] : _GEN_2316; // @[Execute.scala 117:10]
  assign _GEN_2318 = 6'hc == _T_264 ? welem[12] : _GEN_2317; // @[Execute.scala 117:10]
  assign _GEN_2319 = 6'hd == _T_264 ? welem[13] : _GEN_2318; // @[Execute.scala 117:10]
  assign _GEN_2320 = 6'he == _T_264 ? welem[14] : _GEN_2319; // @[Execute.scala 117:10]
  assign _GEN_2321 = 6'hf == _T_264 ? welem[15] : _GEN_2320; // @[Execute.scala 117:10]
  assign _GEN_2322 = 6'h10 == _T_264 ? welem[16] : _GEN_2321; // @[Execute.scala 117:10]
  assign _GEN_2323 = 6'h11 == _T_264 ? welem[17] : _GEN_2322; // @[Execute.scala 117:10]
  assign _GEN_2324 = 6'h12 == _T_264 ? welem[18] : _GEN_2323; // @[Execute.scala 117:10]
  assign _GEN_2325 = 6'h13 == _T_264 ? welem[19] : _GEN_2324; // @[Execute.scala 117:10]
  assign _GEN_2326 = 6'h14 == _T_264 ? welem[20] : _GEN_2325; // @[Execute.scala 117:10]
  assign _GEN_2327 = 6'h15 == _T_264 ? welem[21] : _GEN_2326; // @[Execute.scala 117:10]
  assign _GEN_2328 = 6'h16 == _T_264 ? welem[22] : _GEN_2327; // @[Execute.scala 117:10]
  assign _GEN_2329 = 6'h17 == _T_264 ? welem[23] : _GEN_2328; // @[Execute.scala 117:10]
  assign _GEN_2330 = 6'h18 == _T_264 ? welem[24] : _GEN_2329; // @[Execute.scala 117:10]
  assign _GEN_2331 = 6'h19 == _T_264 ? welem[25] : _GEN_2330; // @[Execute.scala 117:10]
  assign _GEN_2332 = 6'h1a == _T_264 ? welem[26] : _GEN_2331; // @[Execute.scala 117:10]
  assign _GEN_2333 = 6'h1b == _T_264 ? welem[27] : _GEN_2332; // @[Execute.scala 117:10]
  assign _GEN_2334 = 6'h1c == _T_264 ? welem[28] : _GEN_2333; // @[Execute.scala 117:10]
  assign _GEN_2335 = 6'h1d == _T_264 ? welem[29] : _GEN_2334; // @[Execute.scala 117:10]
  assign _GEN_2336 = 6'h1e == _T_264 ? welem[30] : _GEN_2335; // @[Execute.scala 117:10]
  assign _GEN_2337 = 6'h1f == _T_264 ? welem[31] : _GEN_2336; // @[Execute.scala 117:10]
  assign _GEN_2338 = 6'h20 == _T_264 ? welem[32] : _GEN_2337; // @[Execute.scala 117:10]
  assign _GEN_2339 = 6'h21 == _T_264 ? welem[33] : _GEN_2338; // @[Execute.scala 117:10]
  assign _GEN_2340 = 6'h22 == _T_264 ? welem[34] : _GEN_2339; // @[Execute.scala 117:10]
  assign _GEN_2341 = 6'h23 == _T_264 ? welem[35] : _GEN_2340; // @[Execute.scala 117:10]
  assign _GEN_2342 = 6'h24 == _T_264 ? welem[36] : _GEN_2341; // @[Execute.scala 117:10]
  assign _GEN_2343 = 6'h25 == _T_264 ? welem[37] : _GEN_2342; // @[Execute.scala 117:10]
  assign _GEN_2344 = 6'h26 == _T_264 ? welem[38] : _GEN_2343; // @[Execute.scala 117:10]
  assign _GEN_2345 = 6'h27 == _T_264 ? welem[39] : _GEN_2344; // @[Execute.scala 117:10]
  assign _GEN_2346 = 6'h28 == _T_264 ? welem[40] : _GEN_2345; // @[Execute.scala 117:10]
  assign _GEN_2347 = 6'h29 == _T_264 ? welem[41] : _GEN_2346; // @[Execute.scala 117:10]
  assign _GEN_2348 = 6'h2a == _T_264 ? welem[42] : _GEN_2347; // @[Execute.scala 117:10]
  assign _GEN_2349 = 6'h2b == _T_264 ? welem[43] : _GEN_2348; // @[Execute.scala 117:10]
  assign _GEN_2350 = 6'h2c == _T_264 ? welem[44] : _GEN_2349; // @[Execute.scala 117:10]
  assign _GEN_2351 = 6'h2d == _T_264 ? welem[45] : _GEN_2350; // @[Execute.scala 117:10]
  assign _GEN_2352 = 6'h2e == _T_264 ? welem[46] : _GEN_2351; // @[Execute.scala 117:10]
  assign _GEN_2353 = 6'h2f == _T_264 ? welem[47] : _GEN_2352; // @[Execute.scala 117:10]
  assign _GEN_2354 = 6'h30 == _T_264 ? welem[48] : _GEN_2353; // @[Execute.scala 117:10]
  assign _GEN_2355 = 6'h31 == _T_264 ? welem[49] : _GEN_2354; // @[Execute.scala 117:10]
  assign _GEN_2356 = 6'h32 == _T_264 ? welem[50] : _GEN_2355; // @[Execute.scala 117:10]
  assign _GEN_2357 = 6'h33 == _T_264 ? welem[51] : _GEN_2356; // @[Execute.scala 117:10]
  assign _GEN_2358 = 6'h34 == _T_264 ? welem[52] : _GEN_2357; // @[Execute.scala 117:10]
  assign _GEN_2359 = 6'h35 == _T_264 ? welem[53] : _GEN_2358; // @[Execute.scala 117:10]
  assign _GEN_2360 = 6'h36 == _T_264 ? welem[54] : _GEN_2359; // @[Execute.scala 117:10]
  assign _GEN_2361 = 6'h37 == _T_264 ? welem[55] : _GEN_2360; // @[Execute.scala 117:10]
  assign _GEN_2362 = 6'h38 == _T_264 ? welem[56] : _GEN_2361; // @[Execute.scala 117:10]
  assign _GEN_2363 = 6'h39 == _T_264 ? welem[57] : _GEN_2362; // @[Execute.scala 117:10]
  assign _GEN_2364 = 6'h3a == _T_264 ? welem[58] : _GEN_2363; // @[Execute.scala 117:10]
  assign _GEN_2365 = 6'h3b == _T_264 ? welem[59] : _GEN_2364; // @[Execute.scala 117:10]
  assign _GEN_2366 = 6'h3c == _T_264 ? welem[60] : _GEN_2365; // @[Execute.scala 117:10]
  assign _GEN_2367 = 6'h3d == _T_264 ? welem[61] : _GEN_2366; // @[Execute.scala 117:10]
  assign _GEN_2368 = 6'h3e == _T_264 ? welem[62] : _GEN_2367; // @[Execute.scala 117:10]
  assign _GEN_2369 = 6'h3f == _T_264 ? welem[63] : _GEN_2368; // @[Execute.scala 117:10]
  assign _GEN_2371 = 6'h1 == _T_268 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2372 = 6'h2 == _T_268 ? welem[2] : _GEN_2371; // @[Execute.scala 117:10]
  assign _GEN_2373 = 6'h3 == _T_268 ? welem[3] : _GEN_2372; // @[Execute.scala 117:10]
  assign _GEN_2374 = 6'h4 == _T_268 ? welem[4] : _GEN_2373; // @[Execute.scala 117:10]
  assign _GEN_2375 = 6'h5 == _T_268 ? welem[5] : _GEN_2374; // @[Execute.scala 117:10]
  assign _GEN_2376 = 6'h6 == _T_268 ? welem[6] : _GEN_2375; // @[Execute.scala 117:10]
  assign _GEN_2377 = 6'h7 == _T_268 ? welem[7] : _GEN_2376; // @[Execute.scala 117:10]
  assign _GEN_2378 = 6'h8 == _T_268 ? welem[8] : _GEN_2377; // @[Execute.scala 117:10]
  assign _GEN_2379 = 6'h9 == _T_268 ? welem[9] : _GEN_2378; // @[Execute.scala 117:10]
  assign _GEN_2380 = 6'ha == _T_268 ? welem[10] : _GEN_2379; // @[Execute.scala 117:10]
  assign _GEN_2381 = 6'hb == _T_268 ? welem[11] : _GEN_2380; // @[Execute.scala 117:10]
  assign _GEN_2382 = 6'hc == _T_268 ? welem[12] : _GEN_2381; // @[Execute.scala 117:10]
  assign _GEN_2383 = 6'hd == _T_268 ? welem[13] : _GEN_2382; // @[Execute.scala 117:10]
  assign _GEN_2384 = 6'he == _T_268 ? welem[14] : _GEN_2383; // @[Execute.scala 117:10]
  assign _GEN_2385 = 6'hf == _T_268 ? welem[15] : _GEN_2384; // @[Execute.scala 117:10]
  assign _GEN_2386 = 6'h10 == _T_268 ? welem[16] : _GEN_2385; // @[Execute.scala 117:10]
  assign _GEN_2387 = 6'h11 == _T_268 ? welem[17] : _GEN_2386; // @[Execute.scala 117:10]
  assign _GEN_2388 = 6'h12 == _T_268 ? welem[18] : _GEN_2387; // @[Execute.scala 117:10]
  assign _GEN_2389 = 6'h13 == _T_268 ? welem[19] : _GEN_2388; // @[Execute.scala 117:10]
  assign _GEN_2390 = 6'h14 == _T_268 ? welem[20] : _GEN_2389; // @[Execute.scala 117:10]
  assign _GEN_2391 = 6'h15 == _T_268 ? welem[21] : _GEN_2390; // @[Execute.scala 117:10]
  assign _GEN_2392 = 6'h16 == _T_268 ? welem[22] : _GEN_2391; // @[Execute.scala 117:10]
  assign _GEN_2393 = 6'h17 == _T_268 ? welem[23] : _GEN_2392; // @[Execute.scala 117:10]
  assign _GEN_2394 = 6'h18 == _T_268 ? welem[24] : _GEN_2393; // @[Execute.scala 117:10]
  assign _GEN_2395 = 6'h19 == _T_268 ? welem[25] : _GEN_2394; // @[Execute.scala 117:10]
  assign _GEN_2396 = 6'h1a == _T_268 ? welem[26] : _GEN_2395; // @[Execute.scala 117:10]
  assign _GEN_2397 = 6'h1b == _T_268 ? welem[27] : _GEN_2396; // @[Execute.scala 117:10]
  assign _GEN_2398 = 6'h1c == _T_268 ? welem[28] : _GEN_2397; // @[Execute.scala 117:10]
  assign _GEN_2399 = 6'h1d == _T_268 ? welem[29] : _GEN_2398; // @[Execute.scala 117:10]
  assign _GEN_2400 = 6'h1e == _T_268 ? welem[30] : _GEN_2399; // @[Execute.scala 117:10]
  assign _GEN_2401 = 6'h1f == _T_268 ? welem[31] : _GEN_2400; // @[Execute.scala 117:10]
  assign _GEN_2402 = 6'h20 == _T_268 ? welem[32] : _GEN_2401; // @[Execute.scala 117:10]
  assign _GEN_2403 = 6'h21 == _T_268 ? welem[33] : _GEN_2402; // @[Execute.scala 117:10]
  assign _GEN_2404 = 6'h22 == _T_268 ? welem[34] : _GEN_2403; // @[Execute.scala 117:10]
  assign _GEN_2405 = 6'h23 == _T_268 ? welem[35] : _GEN_2404; // @[Execute.scala 117:10]
  assign _GEN_2406 = 6'h24 == _T_268 ? welem[36] : _GEN_2405; // @[Execute.scala 117:10]
  assign _GEN_2407 = 6'h25 == _T_268 ? welem[37] : _GEN_2406; // @[Execute.scala 117:10]
  assign _GEN_2408 = 6'h26 == _T_268 ? welem[38] : _GEN_2407; // @[Execute.scala 117:10]
  assign _GEN_2409 = 6'h27 == _T_268 ? welem[39] : _GEN_2408; // @[Execute.scala 117:10]
  assign _GEN_2410 = 6'h28 == _T_268 ? welem[40] : _GEN_2409; // @[Execute.scala 117:10]
  assign _GEN_2411 = 6'h29 == _T_268 ? welem[41] : _GEN_2410; // @[Execute.scala 117:10]
  assign _GEN_2412 = 6'h2a == _T_268 ? welem[42] : _GEN_2411; // @[Execute.scala 117:10]
  assign _GEN_2413 = 6'h2b == _T_268 ? welem[43] : _GEN_2412; // @[Execute.scala 117:10]
  assign _GEN_2414 = 6'h2c == _T_268 ? welem[44] : _GEN_2413; // @[Execute.scala 117:10]
  assign _GEN_2415 = 6'h2d == _T_268 ? welem[45] : _GEN_2414; // @[Execute.scala 117:10]
  assign _GEN_2416 = 6'h2e == _T_268 ? welem[46] : _GEN_2415; // @[Execute.scala 117:10]
  assign _GEN_2417 = 6'h2f == _T_268 ? welem[47] : _GEN_2416; // @[Execute.scala 117:10]
  assign _GEN_2418 = 6'h30 == _T_268 ? welem[48] : _GEN_2417; // @[Execute.scala 117:10]
  assign _GEN_2419 = 6'h31 == _T_268 ? welem[49] : _GEN_2418; // @[Execute.scala 117:10]
  assign _GEN_2420 = 6'h32 == _T_268 ? welem[50] : _GEN_2419; // @[Execute.scala 117:10]
  assign _GEN_2421 = 6'h33 == _T_268 ? welem[51] : _GEN_2420; // @[Execute.scala 117:10]
  assign _GEN_2422 = 6'h34 == _T_268 ? welem[52] : _GEN_2421; // @[Execute.scala 117:10]
  assign _GEN_2423 = 6'h35 == _T_268 ? welem[53] : _GEN_2422; // @[Execute.scala 117:10]
  assign _GEN_2424 = 6'h36 == _T_268 ? welem[54] : _GEN_2423; // @[Execute.scala 117:10]
  assign _GEN_2425 = 6'h37 == _T_268 ? welem[55] : _GEN_2424; // @[Execute.scala 117:10]
  assign _GEN_2426 = 6'h38 == _T_268 ? welem[56] : _GEN_2425; // @[Execute.scala 117:10]
  assign _GEN_2427 = 6'h39 == _T_268 ? welem[57] : _GEN_2426; // @[Execute.scala 117:10]
  assign _GEN_2428 = 6'h3a == _T_268 ? welem[58] : _GEN_2427; // @[Execute.scala 117:10]
  assign _GEN_2429 = 6'h3b == _T_268 ? welem[59] : _GEN_2428; // @[Execute.scala 117:10]
  assign _GEN_2430 = 6'h3c == _T_268 ? welem[60] : _GEN_2429; // @[Execute.scala 117:10]
  assign _GEN_2431 = 6'h3d == _T_268 ? welem[61] : _GEN_2430; // @[Execute.scala 117:10]
  assign _GEN_2432 = 6'h3e == _T_268 ? welem[62] : _GEN_2431; // @[Execute.scala 117:10]
  assign _GEN_2433 = 6'h3f == _T_268 ? welem[63] : _GEN_2432; // @[Execute.scala 117:10]
  assign _T_271 = _T_262 ? _GEN_2369 : _GEN_2433; // @[Execute.scala 117:10]
  assign _T_272 = r < 6'h2e; // @[Execute.scala 117:15]
  assign _T_274 = r - 6'h2e; // @[Execute.scala 117:37]
  assign _T_278 = 6'h12 + r; // @[Execute.scala 117:60]
  assign _GEN_2435 = 6'h1 == _T_274 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2436 = 6'h2 == _T_274 ? welem[2] : _GEN_2435; // @[Execute.scala 117:10]
  assign _GEN_2437 = 6'h3 == _T_274 ? welem[3] : _GEN_2436; // @[Execute.scala 117:10]
  assign _GEN_2438 = 6'h4 == _T_274 ? welem[4] : _GEN_2437; // @[Execute.scala 117:10]
  assign _GEN_2439 = 6'h5 == _T_274 ? welem[5] : _GEN_2438; // @[Execute.scala 117:10]
  assign _GEN_2440 = 6'h6 == _T_274 ? welem[6] : _GEN_2439; // @[Execute.scala 117:10]
  assign _GEN_2441 = 6'h7 == _T_274 ? welem[7] : _GEN_2440; // @[Execute.scala 117:10]
  assign _GEN_2442 = 6'h8 == _T_274 ? welem[8] : _GEN_2441; // @[Execute.scala 117:10]
  assign _GEN_2443 = 6'h9 == _T_274 ? welem[9] : _GEN_2442; // @[Execute.scala 117:10]
  assign _GEN_2444 = 6'ha == _T_274 ? welem[10] : _GEN_2443; // @[Execute.scala 117:10]
  assign _GEN_2445 = 6'hb == _T_274 ? welem[11] : _GEN_2444; // @[Execute.scala 117:10]
  assign _GEN_2446 = 6'hc == _T_274 ? welem[12] : _GEN_2445; // @[Execute.scala 117:10]
  assign _GEN_2447 = 6'hd == _T_274 ? welem[13] : _GEN_2446; // @[Execute.scala 117:10]
  assign _GEN_2448 = 6'he == _T_274 ? welem[14] : _GEN_2447; // @[Execute.scala 117:10]
  assign _GEN_2449 = 6'hf == _T_274 ? welem[15] : _GEN_2448; // @[Execute.scala 117:10]
  assign _GEN_2450 = 6'h10 == _T_274 ? welem[16] : _GEN_2449; // @[Execute.scala 117:10]
  assign _GEN_2451 = 6'h11 == _T_274 ? welem[17] : _GEN_2450; // @[Execute.scala 117:10]
  assign _GEN_2452 = 6'h12 == _T_274 ? welem[18] : _GEN_2451; // @[Execute.scala 117:10]
  assign _GEN_2453 = 6'h13 == _T_274 ? welem[19] : _GEN_2452; // @[Execute.scala 117:10]
  assign _GEN_2454 = 6'h14 == _T_274 ? welem[20] : _GEN_2453; // @[Execute.scala 117:10]
  assign _GEN_2455 = 6'h15 == _T_274 ? welem[21] : _GEN_2454; // @[Execute.scala 117:10]
  assign _GEN_2456 = 6'h16 == _T_274 ? welem[22] : _GEN_2455; // @[Execute.scala 117:10]
  assign _GEN_2457 = 6'h17 == _T_274 ? welem[23] : _GEN_2456; // @[Execute.scala 117:10]
  assign _GEN_2458 = 6'h18 == _T_274 ? welem[24] : _GEN_2457; // @[Execute.scala 117:10]
  assign _GEN_2459 = 6'h19 == _T_274 ? welem[25] : _GEN_2458; // @[Execute.scala 117:10]
  assign _GEN_2460 = 6'h1a == _T_274 ? welem[26] : _GEN_2459; // @[Execute.scala 117:10]
  assign _GEN_2461 = 6'h1b == _T_274 ? welem[27] : _GEN_2460; // @[Execute.scala 117:10]
  assign _GEN_2462 = 6'h1c == _T_274 ? welem[28] : _GEN_2461; // @[Execute.scala 117:10]
  assign _GEN_2463 = 6'h1d == _T_274 ? welem[29] : _GEN_2462; // @[Execute.scala 117:10]
  assign _GEN_2464 = 6'h1e == _T_274 ? welem[30] : _GEN_2463; // @[Execute.scala 117:10]
  assign _GEN_2465 = 6'h1f == _T_274 ? welem[31] : _GEN_2464; // @[Execute.scala 117:10]
  assign _GEN_2466 = 6'h20 == _T_274 ? welem[32] : _GEN_2465; // @[Execute.scala 117:10]
  assign _GEN_2467 = 6'h21 == _T_274 ? welem[33] : _GEN_2466; // @[Execute.scala 117:10]
  assign _GEN_2468 = 6'h22 == _T_274 ? welem[34] : _GEN_2467; // @[Execute.scala 117:10]
  assign _GEN_2469 = 6'h23 == _T_274 ? welem[35] : _GEN_2468; // @[Execute.scala 117:10]
  assign _GEN_2470 = 6'h24 == _T_274 ? welem[36] : _GEN_2469; // @[Execute.scala 117:10]
  assign _GEN_2471 = 6'h25 == _T_274 ? welem[37] : _GEN_2470; // @[Execute.scala 117:10]
  assign _GEN_2472 = 6'h26 == _T_274 ? welem[38] : _GEN_2471; // @[Execute.scala 117:10]
  assign _GEN_2473 = 6'h27 == _T_274 ? welem[39] : _GEN_2472; // @[Execute.scala 117:10]
  assign _GEN_2474 = 6'h28 == _T_274 ? welem[40] : _GEN_2473; // @[Execute.scala 117:10]
  assign _GEN_2475 = 6'h29 == _T_274 ? welem[41] : _GEN_2474; // @[Execute.scala 117:10]
  assign _GEN_2476 = 6'h2a == _T_274 ? welem[42] : _GEN_2475; // @[Execute.scala 117:10]
  assign _GEN_2477 = 6'h2b == _T_274 ? welem[43] : _GEN_2476; // @[Execute.scala 117:10]
  assign _GEN_2478 = 6'h2c == _T_274 ? welem[44] : _GEN_2477; // @[Execute.scala 117:10]
  assign _GEN_2479 = 6'h2d == _T_274 ? welem[45] : _GEN_2478; // @[Execute.scala 117:10]
  assign _GEN_2480 = 6'h2e == _T_274 ? welem[46] : _GEN_2479; // @[Execute.scala 117:10]
  assign _GEN_2481 = 6'h2f == _T_274 ? welem[47] : _GEN_2480; // @[Execute.scala 117:10]
  assign _GEN_2482 = 6'h30 == _T_274 ? welem[48] : _GEN_2481; // @[Execute.scala 117:10]
  assign _GEN_2483 = 6'h31 == _T_274 ? welem[49] : _GEN_2482; // @[Execute.scala 117:10]
  assign _GEN_2484 = 6'h32 == _T_274 ? welem[50] : _GEN_2483; // @[Execute.scala 117:10]
  assign _GEN_2485 = 6'h33 == _T_274 ? welem[51] : _GEN_2484; // @[Execute.scala 117:10]
  assign _GEN_2486 = 6'h34 == _T_274 ? welem[52] : _GEN_2485; // @[Execute.scala 117:10]
  assign _GEN_2487 = 6'h35 == _T_274 ? welem[53] : _GEN_2486; // @[Execute.scala 117:10]
  assign _GEN_2488 = 6'h36 == _T_274 ? welem[54] : _GEN_2487; // @[Execute.scala 117:10]
  assign _GEN_2489 = 6'h37 == _T_274 ? welem[55] : _GEN_2488; // @[Execute.scala 117:10]
  assign _GEN_2490 = 6'h38 == _T_274 ? welem[56] : _GEN_2489; // @[Execute.scala 117:10]
  assign _GEN_2491 = 6'h39 == _T_274 ? welem[57] : _GEN_2490; // @[Execute.scala 117:10]
  assign _GEN_2492 = 6'h3a == _T_274 ? welem[58] : _GEN_2491; // @[Execute.scala 117:10]
  assign _GEN_2493 = 6'h3b == _T_274 ? welem[59] : _GEN_2492; // @[Execute.scala 117:10]
  assign _GEN_2494 = 6'h3c == _T_274 ? welem[60] : _GEN_2493; // @[Execute.scala 117:10]
  assign _GEN_2495 = 6'h3d == _T_274 ? welem[61] : _GEN_2494; // @[Execute.scala 117:10]
  assign _GEN_2496 = 6'h3e == _T_274 ? welem[62] : _GEN_2495; // @[Execute.scala 117:10]
  assign _GEN_2497 = 6'h3f == _T_274 ? welem[63] : _GEN_2496; // @[Execute.scala 117:10]
  assign _GEN_2499 = 6'h1 == _T_278 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2500 = 6'h2 == _T_278 ? welem[2] : _GEN_2499; // @[Execute.scala 117:10]
  assign _GEN_2501 = 6'h3 == _T_278 ? welem[3] : _GEN_2500; // @[Execute.scala 117:10]
  assign _GEN_2502 = 6'h4 == _T_278 ? welem[4] : _GEN_2501; // @[Execute.scala 117:10]
  assign _GEN_2503 = 6'h5 == _T_278 ? welem[5] : _GEN_2502; // @[Execute.scala 117:10]
  assign _GEN_2504 = 6'h6 == _T_278 ? welem[6] : _GEN_2503; // @[Execute.scala 117:10]
  assign _GEN_2505 = 6'h7 == _T_278 ? welem[7] : _GEN_2504; // @[Execute.scala 117:10]
  assign _GEN_2506 = 6'h8 == _T_278 ? welem[8] : _GEN_2505; // @[Execute.scala 117:10]
  assign _GEN_2507 = 6'h9 == _T_278 ? welem[9] : _GEN_2506; // @[Execute.scala 117:10]
  assign _GEN_2508 = 6'ha == _T_278 ? welem[10] : _GEN_2507; // @[Execute.scala 117:10]
  assign _GEN_2509 = 6'hb == _T_278 ? welem[11] : _GEN_2508; // @[Execute.scala 117:10]
  assign _GEN_2510 = 6'hc == _T_278 ? welem[12] : _GEN_2509; // @[Execute.scala 117:10]
  assign _GEN_2511 = 6'hd == _T_278 ? welem[13] : _GEN_2510; // @[Execute.scala 117:10]
  assign _GEN_2512 = 6'he == _T_278 ? welem[14] : _GEN_2511; // @[Execute.scala 117:10]
  assign _GEN_2513 = 6'hf == _T_278 ? welem[15] : _GEN_2512; // @[Execute.scala 117:10]
  assign _GEN_2514 = 6'h10 == _T_278 ? welem[16] : _GEN_2513; // @[Execute.scala 117:10]
  assign _GEN_2515 = 6'h11 == _T_278 ? welem[17] : _GEN_2514; // @[Execute.scala 117:10]
  assign _GEN_2516 = 6'h12 == _T_278 ? welem[18] : _GEN_2515; // @[Execute.scala 117:10]
  assign _GEN_2517 = 6'h13 == _T_278 ? welem[19] : _GEN_2516; // @[Execute.scala 117:10]
  assign _GEN_2518 = 6'h14 == _T_278 ? welem[20] : _GEN_2517; // @[Execute.scala 117:10]
  assign _GEN_2519 = 6'h15 == _T_278 ? welem[21] : _GEN_2518; // @[Execute.scala 117:10]
  assign _GEN_2520 = 6'h16 == _T_278 ? welem[22] : _GEN_2519; // @[Execute.scala 117:10]
  assign _GEN_2521 = 6'h17 == _T_278 ? welem[23] : _GEN_2520; // @[Execute.scala 117:10]
  assign _GEN_2522 = 6'h18 == _T_278 ? welem[24] : _GEN_2521; // @[Execute.scala 117:10]
  assign _GEN_2523 = 6'h19 == _T_278 ? welem[25] : _GEN_2522; // @[Execute.scala 117:10]
  assign _GEN_2524 = 6'h1a == _T_278 ? welem[26] : _GEN_2523; // @[Execute.scala 117:10]
  assign _GEN_2525 = 6'h1b == _T_278 ? welem[27] : _GEN_2524; // @[Execute.scala 117:10]
  assign _GEN_2526 = 6'h1c == _T_278 ? welem[28] : _GEN_2525; // @[Execute.scala 117:10]
  assign _GEN_2527 = 6'h1d == _T_278 ? welem[29] : _GEN_2526; // @[Execute.scala 117:10]
  assign _GEN_2528 = 6'h1e == _T_278 ? welem[30] : _GEN_2527; // @[Execute.scala 117:10]
  assign _GEN_2529 = 6'h1f == _T_278 ? welem[31] : _GEN_2528; // @[Execute.scala 117:10]
  assign _GEN_2530 = 6'h20 == _T_278 ? welem[32] : _GEN_2529; // @[Execute.scala 117:10]
  assign _GEN_2531 = 6'h21 == _T_278 ? welem[33] : _GEN_2530; // @[Execute.scala 117:10]
  assign _GEN_2532 = 6'h22 == _T_278 ? welem[34] : _GEN_2531; // @[Execute.scala 117:10]
  assign _GEN_2533 = 6'h23 == _T_278 ? welem[35] : _GEN_2532; // @[Execute.scala 117:10]
  assign _GEN_2534 = 6'h24 == _T_278 ? welem[36] : _GEN_2533; // @[Execute.scala 117:10]
  assign _GEN_2535 = 6'h25 == _T_278 ? welem[37] : _GEN_2534; // @[Execute.scala 117:10]
  assign _GEN_2536 = 6'h26 == _T_278 ? welem[38] : _GEN_2535; // @[Execute.scala 117:10]
  assign _GEN_2537 = 6'h27 == _T_278 ? welem[39] : _GEN_2536; // @[Execute.scala 117:10]
  assign _GEN_2538 = 6'h28 == _T_278 ? welem[40] : _GEN_2537; // @[Execute.scala 117:10]
  assign _GEN_2539 = 6'h29 == _T_278 ? welem[41] : _GEN_2538; // @[Execute.scala 117:10]
  assign _GEN_2540 = 6'h2a == _T_278 ? welem[42] : _GEN_2539; // @[Execute.scala 117:10]
  assign _GEN_2541 = 6'h2b == _T_278 ? welem[43] : _GEN_2540; // @[Execute.scala 117:10]
  assign _GEN_2542 = 6'h2c == _T_278 ? welem[44] : _GEN_2541; // @[Execute.scala 117:10]
  assign _GEN_2543 = 6'h2d == _T_278 ? welem[45] : _GEN_2542; // @[Execute.scala 117:10]
  assign _GEN_2544 = 6'h2e == _T_278 ? welem[46] : _GEN_2543; // @[Execute.scala 117:10]
  assign _GEN_2545 = 6'h2f == _T_278 ? welem[47] : _GEN_2544; // @[Execute.scala 117:10]
  assign _GEN_2546 = 6'h30 == _T_278 ? welem[48] : _GEN_2545; // @[Execute.scala 117:10]
  assign _GEN_2547 = 6'h31 == _T_278 ? welem[49] : _GEN_2546; // @[Execute.scala 117:10]
  assign _GEN_2548 = 6'h32 == _T_278 ? welem[50] : _GEN_2547; // @[Execute.scala 117:10]
  assign _GEN_2549 = 6'h33 == _T_278 ? welem[51] : _GEN_2548; // @[Execute.scala 117:10]
  assign _GEN_2550 = 6'h34 == _T_278 ? welem[52] : _GEN_2549; // @[Execute.scala 117:10]
  assign _GEN_2551 = 6'h35 == _T_278 ? welem[53] : _GEN_2550; // @[Execute.scala 117:10]
  assign _GEN_2552 = 6'h36 == _T_278 ? welem[54] : _GEN_2551; // @[Execute.scala 117:10]
  assign _GEN_2553 = 6'h37 == _T_278 ? welem[55] : _GEN_2552; // @[Execute.scala 117:10]
  assign _GEN_2554 = 6'h38 == _T_278 ? welem[56] : _GEN_2553; // @[Execute.scala 117:10]
  assign _GEN_2555 = 6'h39 == _T_278 ? welem[57] : _GEN_2554; // @[Execute.scala 117:10]
  assign _GEN_2556 = 6'h3a == _T_278 ? welem[58] : _GEN_2555; // @[Execute.scala 117:10]
  assign _GEN_2557 = 6'h3b == _T_278 ? welem[59] : _GEN_2556; // @[Execute.scala 117:10]
  assign _GEN_2558 = 6'h3c == _T_278 ? welem[60] : _GEN_2557; // @[Execute.scala 117:10]
  assign _GEN_2559 = 6'h3d == _T_278 ? welem[61] : _GEN_2558; // @[Execute.scala 117:10]
  assign _GEN_2560 = 6'h3e == _T_278 ? welem[62] : _GEN_2559; // @[Execute.scala 117:10]
  assign _GEN_2561 = 6'h3f == _T_278 ? welem[63] : _GEN_2560; // @[Execute.scala 117:10]
  assign _T_281 = _T_272 ? _GEN_2497 : _GEN_2561; // @[Execute.scala 117:10]
  assign _T_282 = r < 6'h2d; // @[Execute.scala 117:15]
  assign _T_284 = r - 6'h2d; // @[Execute.scala 117:37]
  assign _T_288 = 6'h13 + r; // @[Execute.scala 117:60]
  assign _GEN_2563 = 6'h1 == _T_284 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2564 = 6'h2 == _T_284 ? welem[2] : _GEN_2563; // @[Execute.scala 117:10]
  assign _GEN_2565 = 6'h3 == _T_284 ? welem[3] : _GEN_2564; // @[Execute.scala 117:10]
  assign _GEN_2566 = 6'h4 == _T_284 ? welem[4] : _GEN_2565; // @[Execute.scala 117:10]
  assign _GEN_2567 = 6'h5 == _T_284 ? welem[5] : _GEN_2566; // @[Execute.scala 117:10]
  assign _GEN_2568 = 6'h6 == _T_284 ? welem[6] : _GEN_2567; // @[Execute.scala 117:10]
  assign _GEN_2569 = 6'h7 == _T_284 ? welem[7] : _GEN_2568; // @[Execute.scala 117:10]
  assign _GEN_2570 = 6'h8 == _T_284 ? welem[8] : _GEN_2569; // @[Execute.scala 117:10]
  assign _GEN_2571 = 6'h9 == _T_284 ? welem[9] : _GEN_2570; // @[Execute.scala 117:10]
  assign _GEN_2572 = 6'ha == _T_284 ? welem[10] : _GEN_2571; // @[Execute.scala 117:10]
  assign _GEN_2573 = 6'hb == _T_284 ? welem[11] : _GEN_2572; // @[Execute.scala 117:10]
  assign _GEN_2574 = 6'hc == _T_284 ? welem[12] : _GEN_2573; // @[Execute.scala 117:10]
  assign _GEN_2575 = 6'hd == _T_284 ? welem[13] : _GEN_2574; // @[Execute.scala 117:10]
  assign _GEN_2576 = 6'he == _T_284 ? welem[14] : _GEN_2575; // @[Execute.scala 117:10]
  assign _GEN_2577 = 6'hf == _T_284 ? welem[15] : _GEN_2576; // @[Execute.scala 117:10]
  assign _GEN_2578 = 6'h10 == _T_284 ? welem[16] : _GEN_2577; // @[Execute.scala 117:10]
  assign _GEN_2579 = 6'h11 == _T_284 ? welem[17] : _GEN_2578; // @[Execute.scala 117:10]
  assign _GEN_2580 = 6'h12 == _T_284 ? welem[18] : _GEN_2579; // @[Execute.scala 117:10]
  assign _GEN_2581 = 6'h13 == _T_284 ? welem[19] : _GEN_2580; // @[Execute.scala 117:10]
  assign _GEN_2582 = 6'h14 == _T_284 ? welem[20] : _GEN_2581; // @[Execute.scala 117:10]
  assign _GEN_2583 = 6'h15 == _T_284 ? welem[21] : _GEN_2582; // @[Execute.scala 117:10]
  assign _GEN_2584 = 6'h16 == _T_284 ? welem[22] : _GEN_2583; // @[Execute.scala 117:10]
  assign _GEN_2585 = 6'h17 == _T_284 ? welem[23] : _GEN_2584; // @[Execute.scala 117:10]
  assign _GEN_2586 = 6'h18 == _T_284 ? welem[24] : _GEN_2585; // @[Execute.scala 117:10]
  assign _GEN_2587 = 6'h19 == _T_284 ? welem[25] : _GEN_2586; // @[Execute.scala 117:10]
  assign _GEN_2588 = 6'h1a == _T_284 ? welem[26] : _GEN_2587; // @[Execute.scala 117:10]
  assign _GEN_2589 = 6'h1b == _T_284 ? welem[27] : _GEN_2588; // @[Execute.scala 117:10]
  assign _GEN_2590 = 6'h1c == _T_284 ? welem[28] : _GEN_2589; // @[Execute.scala 117:10]
  assign _GEN_2591 = 6'h1d == _T_284 ? welem[29] : _GEN_2590; // @[Execute.scala 117:10]
  assign _GEN_2592 = 6'h1e == _T_284 ? welem[30] : _GEN_2591; // @[Execute.scala 117:10]
  assign _GEN_2593 = 6'h1f == _T_284 ? welem[31] : _GEN_2592; // @[Execute.scala 117:10]
  assign _GEN_2594 = 6'h20 == _T_284 ? welem[32] : _GEN_2593; // @[Execute.scala 117:10]
  assign _GEN_2595 = 6'h21 == _T_284 ? welem[33] : _GEN_2594; // @[Execute.scala 117:10]
  assign _GEN_2596 = 6'h22 == _T_284 ? welem[34] : _GEN_2595; // @[Execute.scala 117:10]
  assign _GEN_2597 = 6'h23 == _T_284 ? welem[35] : _GEN_2596; // @[Execute.scala 117:10]
  assign _GEN_2598 = 6'h24 == _T_284 ? welem[36] : _GEN_2597; // @[Execute.scala 117:10]
  assign _GEN_2599 = 6'h25 == _T_284 ? welem[37] : _GEN_2598; // @[Execute.scala 117:10]
  assign _GEN_2600 = 6'h26 == _T_284 ? welem[38] : _GEN_2599; // @[Execute.scala 117:10]
  assign _GEN_2601 = 6'h27 == _T_284 ? welem[39] : _GEN_2600; // @[Execute.scala 117:10]
  assign _GEN_2602 = 6'h28 == _T_284 ? welem[40] : _GEN_2601; // @[Execute.scala 117:10]
  assign _GEN_2603 = 6'h29 == _T_284 ? welem[41] : _GEN_2602; // @[Execute.scala 117:10]
  assign _GEN_2604 = 6'h2a == _T_284 ? welem[42] : _GEN_2603; // @[Execute.scala 117:10]
  assign _GEN_2605 = 6'h2b == _T_284 ? welem[43] : _GEN_2604; // @[Execute.scala 117:10]
  assign _GEN_2606 = 6'h2c == _T_284 ? welem[44] : _GEN_2605; // @[Execute.scala 117:10]
  assign _GEN_2607 = 6'h2d == _T_284 ? welem[45] : _GEN_2606; // @[Execute.scala 117:10]
  assign _GEN_2608 = 6'h2e == _T_284 ? welem[46] : _GEN_2607; // @[Execute.scala 117:10]
  assign _GEN_2609 = 6'h2f == _T_284 ? welem[47] : _GEN_2608; // @[Execute.scala 117:10]
  assign _GEN_2610 = 6'h30 == _T_284 ? welem[48] : _GEN_2609; // @[Execute.scala 117:10]
  assign _GEN_2611 = 6'h31 == _T_284 ? welem[49] : _GEN_2610; // @[Execute.scala 117:10]
  assign _GEN_2612 = 6'h32 == _T_284 ? welem[50] : _GEN_2611; // @[Execute.scala 117:10]
  assign _GEN_2613 = 6'h33 == _T_284 ? welem[51] : _GEN_2612; // @[Execute.scala 117:10]
  assign _GEN_2614 = 6'h34 == _T_284 ? welem[52] : _GEN_2613; // @[Execute.scala 117:10]
  assign _GEN_2615 = 6'h35 == _T_284 ? welem[53] : _GEN_2614; // @[Execute.scala 117:10]
  assign _GEN_2616 = 6'h36 == _T_284 ? welem[54] : _GEN_2615; // @[Execute.scala 117:10]
  assign _GEN_2617 = 6'h37 == _T_284 ? welem[55] : _GEN_2616; // @[Execute.scala 117:10]
  assign _GEN_2618 = 6'h38 == _T_284 ? welem[56] : _GEN_2617; // @[Execute.scala 117:10]
  assign _GEN_2619 = 6'h39 == _T_284 ? welem[57] : _GEN_2618; // @[Execute.scala 117:10]
  assign _GEN_2620 = 6'h3a == _T_284 ? welem[58] : _GEN_2619; // @[Execute.scala 117:10]
  assign _GEN_2621 = 6'h3b == _T_284 ? welem[59] : _GEN_2620; // @[Execute.scala 117:10]
  assign _GEN_2622 = 6'h3c == _T_284 ? welem[60] : _GEN_2621; // @[Execute.scala 117:10]
  assign _GEN_2623 = 6'h3d == _T_284 ? welem[61] : _GEN_2622; // @[Execute.scala 117:10]
  assign _GEN_2624 = 6'h3e == _T_284 ? welem[62] : _GEN_2623; // @[Execute.scala 117:10]
  assign _GEN_2625 = 6'h3f == _T_284 ? welem[63] : _GEN_2624; // @[Execute.scala 117:10]
  assign _GEN_2627 = 6'h1 == _T_288 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2628 = 6'h2 == _T_288 ? welem[2] : _GEN_2627; // @[Execute.scala 117:10]
  assign _GEN_2629 = 6'h3 == _T_288 ? welem[3] : _GEN_2628; // @[Execute.scala 117:10]
  assign _GEN_2630 = 6'h4 == _T_288 ? welem[4] : _GEN_2629; // @[Execute.scala 117:10]
  assign _GEN_2631 = 6'h5 == _T_288 ? welem[5] : _GEN_2630; // @[Execute.scala 117:10]
  assign _GEN_2632 = 6'h6 == _T_288 ? welem[6] : _GEN_2631; // @[Execute.scala 117:10]
  assign _GEN_2633 = 6'h7 == _T_288 ? welem[7] : _GEN_2632; // @[Execute.scala 117:10]
  assign _GEN_2634 = 6'h8 == _T_288 ? welem[8] : _GEN_2633; // @[Execute.scala 117:10]
  assign _GEN_2635 = 6'h9 == _T_288 ? welem[9] : _GEN_2634; // @[Execute.scala 117:10]
  assign _GEN_2636 = 6'ha == _T_288 ? welem[10] : _GEN_2635; // @[Execute.scala 117:10]
  assign _GEN_2637 = 6'hb == _T_288 ? welem[11] : _GEN_2636; // @[Execute.scala 117:10]
  assign _GEN_2638 = 6'hc == _T_288 ? welem[12] : _GEN_2637; // @[Execute.scala 117:10]
  assign _GEN_2639 = 6'hd == _T_288 ? welem[13] : _GEN_2638; // @[Execute.scala 117:10]
  assign _GEN_2640 = 6'he == _T_288 ? welem[14] : _GEN_2639; // @[Execute.scala 117:10]
  assign _GEN_2641 = 6'hf == _T_288 ? welem[15] : _GEN_2640; // @[Execute.scala 117:10]
  assign _GEN_2642 = 6'h10 == _T_288 ? welem[16] : _GEN_2641; // @[Execute.scala 117:10]
  assign _GEN_2643 = 6'h11 == _T_288 ? welem[17] : _GEN_2642; // @[Execute.scala 117:10]
  assign _GEN_2644 = 6'h12 == _T_288 ? welem[18] : _GEN_2643; // @[Execute.scala 117:10]
  assign _GEN_2645 = 6'h13 == _T_288 ? welem[19] : _GEN_2644; // @[Execute.scala 117:10]
  assign _GEN_2646 = 6'h14 == _T_288 ? welem[20] : _GEN_2645; // @[Execute.scala 117:10]
  assign _GEN_2647 = 6'h15 == _T_288 ? welem[21] : _GEN_2646; // @[Execute.scala 117:10]
  assign _GEN_2648 = 6'h16 == _T_288 ? welem[22] : _GEN_2647; // @[Execute.scala 117:10]
  assign _GEN_2649 = 6'h17 == _T_288 ? welem[23] : _GEN_2648; // @[Execute.scala 117:10]
  assign _GEN_2650 = 6'h18 == _T_288 ? welem[24] : _GEN_2649; // @[Execute.scala 117:10]
  assign _GEN_2651 = 6'h19 == _T_288 ? welem[25] : _GEN_2650; // @[Execute.scala 117:10]
  assign _GEN_2652 = 6'h1a == _T_288 ? welem[26] : _GEN_2651; // @[Execute.scala 117:10]
  assign _GEN_2653 = 6'h1b == _T_288 ? welem[27] : _GEN_2652; // @[Execute.scala 117:10]
  assign _GEN_2654 = 6'h1c == _T_288 ? welem[28] : _GEN_2653; // @[Execute.scala 117:10]
  assign _GEN_2655 = 6'h1d == _T_288 ? welem[29] : _GEN_2654; // @[Execute.scala 117:10]
  assign _GEN_2656 = 6'h1e == _T_288 ? welem[30] : _GEN_2655; // @[Execute.scala 117:10]
  assign _GEN_2657 = 6'h1f == _T_288 ? welem[31] : _GEN_2656; // @[Execute.scala 117:10]
  assign _GEN_2658 = 6'h20 == _T_288 ? welem[32] : _GEN_2657; // @[Execute.scala 117:10]
  assign _GEN_2659 = 6'h21 == _T_288 ? welem[33] : _GEN_2658; // @[Execute.scala 117:10]
  assign _GEN_2660 = 6'h22 == _T_288 ? welem[34] : _GEN_2659; // @[Execute.scala 117:10]
  assign _GEN_2661 = 6'h23 == _T_288 ? welem[35] : _GEN_2660; // @[Execute.scala 117:10]
  assign _GEN_2662 = 6'h24 == _T_288 ? welem[36] : _GEN_2661; // @[Execute.scala 117:10]
  assign _GEN_2663 = 6'h25 == _T_288 ? welem[37] : _GEN_2662; // @[Execute.scala 117:10]
  assign _GEN_2664 = 6'h26 == _T_288 ? welem[38] : _GEN_2663; // @[Execute.scala 117:10]
  assign _GEN_2665 = 6'h27 == _T_288 ? welem[39] : _GEN_2664; // @[Execute.scala 117:10]
  assign _GEN_2666 = 6'h28 == _T_288 ? welem[40] : _GEN_2665; // @[Execute.scala 117:10]
  assign _GEN_2667 = 6'h29 == _T_288 ? welem[41] : _GEN_2666; // @[Execute.scala 117:10]
  assign _GEN_2668 = 6'h2a == _T_288 ? welem[42] : _GEN_2667; // @[Execute.scala 117:10]
  assign _GEN_2669 = 6'h2b == _T_288 ? welem[43] : _GEN_2668; // @[Execute.scala 117:10]
  assign _GEN_2670 = 6'h2c == _T_288 ? welem[44] : _GEN_2669; // @[Execute.scala 117:10]
  assign _GEN_2671 = 6'h2d == _T_288 ? welem[45] : _GEN_2670; // @[Execute.scala 117:10]
  assign _GEN_2672 = 6'h2e == _T_288 ? welem[46] : _GEN_2671; // @[Execute.scala 117:10]
  assign _GEN_2673 = 6'h2f == _T_288 ? welem[47] : _GEN_2672; // @[Execute.scala 117:10]
  assign _GEN_2674 = 6'h30 == _T_288 ? welem[48] : _GEN_2673; // @[Execute.scala 117:10]
  assign _GEN_2675 = 6'h31 == _T_288 ? welem[49] : _GEN_2674; // @[Execute.scala 117:10]
  assign _GEN_2676 = 6'h32 == _T_288 ? welem[50] : _GEN_2675; // @[Execute.scala 117:10]
  assign _GEN_2677 = 6'h33 == _T_288 ? welem[51] : _GEN_2676; // @[Execute.scala 117:10]
  assign _GEN_2678 = 6'h34 == _T_288 ? welem[52] : _GEN_2677; // @[Execute.scala 117:10]
  assign _GEN_2679 = 6'h35 == _T_288 ? welem[53] : _GEN_2678; // @[Execute.scala 117:10]
  assign _GEN_2680 = 6'h36 == _T_288 ? welem[54] : _GEN_2679; // @[Execute.scala 117:10]
  assign _GEN_2681 = 6'h37 == _T_288 ? welem[55] : _GEN_2680; // @[Execute.scala 117:10]
  assign _GEN_2682 = 6'h38 == _T_288 ? welem[56] : _GEN_2681; // @[Execute.scala 117:10]
  assign _GEN_2683 = 6'h39 == _T_288 ? welem[57] : _GEN_2682; // @[Execute.scala 117:10]
  assign _GEN_2684 = 6'h3a == _T_288 ? welem[58] : _GEN_2683; // @[Execute.scala 117:10]
  assign _GEN_2685 = 6'h3b == _T_288 ? welem[59] : _GEN_2684; // @[Execute.scala 117:10]
  assign _GEN_2686 = 6'h3c == _T_288 ? welem[60] : _GEN_2685; // @[Execute.scala 117:10]
  assign _GEN_2687 = 6'h3d == _T_288 ? welem[61] : _GEN_2686; // @[Execute.scala 117:10]
  assign _GEN_2688 = 6'h3e == _T_288 ? welem[62] : _GEN_2687; // @[Execute.scala 117:10]
  assign _GEN_2689 = 6'h3f == _T_288 ? welem[63] : _GEN_2688; // @[Execute.scala 117:10]
  assign _T_291 = _T_282 ? _GEN_2625 : _GEN_2689; // @[Execute.scala 117:10]
  assign _T_292 = r < 6'h2c; // @[Execute.scala 117:15]
  assign _T_294 = r - 6'h2c; // @[Execute.scala 117:37]
  assign _T_298 = 6'h14 + r; // @[Execute.scala 117:60]
  assign _GEN_2691 = 6'h1 == _T_294 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2692 = 6'h2 == _T_294 ? welem[2] : _GEN_2691; // @[Execute.scala 117:10]
  assign _GEN_2693 = 6'h3 == _T_294 ? welem[3] : _GEN_2692; // @[Execute.scala 117:10]
  assign _GEN_2694 = 6'h4 == _T_294 ? welem[4] : _GEN_2693; // @[Execute.scala 117:10]
  assign _GEN_2695 = 6'h5 == _T_294 ? welem[5] : _GEN_2694; // @[Execute.scala 117:10]
  assign _GEN_2696 = 6'h6 == _T_294 ? welem[6] : _GEN_2695; // @[Execute.scala 117:10]
  assign _GEN_2697 = 6'h7 == _T_294 ? welem[7] : _GEN_2696; // @[Execute.scala 117:10]
  assign _GEN_2698 = 6'h8 == _T_294 ? welem[8] : _GEN_2697; // @[Execute.scala 117:10]
  assign _GEN_2699 = 6'h9 == _T_294 ? welem[9] : _GEN_2698; // @[Execute.scala 117:10]
  assign _GEN_2700 = 6'ha == _T_294 ? welem[10] : _GEN_2699; // @[Execute.scala 117:10]
  assign _GEN_2701 = 6'hb == _T_294 ? welem[11] : _GEN_2700; // @[Execute.scala 117:10]
  assign _GEN_2702 = 6'hc == _T_294 ? welem[12] : _GEN_2701; // @[Execute.scala 117:10]
  assign _GEN_2703 = 6'hd == _T_294 ? welem[13] : _GEN_2702; // @[Execute.scala 117:10]
  assign _GEN_2704 = 6'he == _T_294 ? welem[14] : _GEN_2703; // @[Execute.scala 117:10]
  assign _GEN_2705 = 6'hf == _T_294 ? welem[15] : _GEN_2704; // @[Execute.scala 117:10]
  assign _GEN_2706 = 6'h10 == _T_294 ? welem[16] : _GEN_2705; // @[Execute.scala 117:10]
  assign _GEN_2707 = 6'h11 == _T_294 ? welem[17] : _GEN_2706; // @[Execute.scala 117:10]
  assign _GEN_2708 = 6'h12 == _T_294 ? welem[18] : _GEN_2707; // @[Execute.scala 117:10]
  assign _GEN_2709 = 6'h13 == _T_294 ? welem[19] : _GEN_2708; // @[Execute.scala 117:10]
  assign _GEN_2710 = 6'h14 == _T_294 ? welem[20] : _GEN_2709; // @[Execute.scala 117:10]
  assign _GEN_2711 = 6'h15 == _T_294 ? welem[21] : _GEN_2710; // @[Execute.scala 117:10]
  assign _GEN_2712 = 6'h16 == _T_294 ? welem[22] : _GEN_2711; // @[Execute.scala 117:10]
  assign _GEN_2713 = 6'h17 == _T_294 ? welem[23] : _GEN_2712; // @[Execute.scala 117:10]
  assign _GEN_2714 = 6'h18 == _T_294 ? welem[24] : _GEN_2713; // @[Execute.scala 117:10]
  assign _GEN_2715 = 6'h19 == _T_294 ? welem[25] : _GEN_2714; // @[Execute.scala 117:10]
  assign _GEN_2716 = 6'h1a == _T_294 ? welem[26] : _GEN_2715; // @[Execute.scala 117:10]
  assign _GEN_2717 = 6'h1b == _T_294 ? welem[27] : _GEN_2716; // @[Execute.scala 117:10]
  assign _GEN_2718 = 6'h1c == _T_294 ? welem[28] : _GEN_2717; // @[Execute.scala 117:10]
  assign _GEN_2719 = 6'h1d == _T_294 ? welem[29] : _GEN_2718; // @[Execute.scala 117:10]
  assign _GEN_2720 = 6'h1e == _T_294 ? welem[30] : _GEN_2719; // @[Execute.scala 117:10]
  assign _GEN_2721 = 6'h1f == _T_294 ? welem[31] : _GEN_2720; // @[Execute.scala 117:10]
  assign _GEN_2722 = 6'h20 == _T_294 ? welem[32] : _GEN_2721; // @[Execute.scala 117:10]
  assign _GEN_2723 = 6'h21 == _T_294 ? welem[33] : _GEN_2722; // @[Execute.scala 117:10]
  assign _GEN_2724 = 6'h22 == _T_294 ? welem[34] : _GEN_2723; // @[Execute.scala 117:10]
  assign _GEN_2725 = 6'h23 == _T_294 ? welem[35] : _GEN_2724; // @[Execute.scala 117:10]
  assign _GEN_2726 = 6'h24 == _T_294 ? welem[36] : _GEN_2725; // @[Execute.scala 117:10]
  assign _GEN_2727 = 6'h25 == _T_294 ? welem[37] : _GEN_2726; // @[Execute.scala 117:10]
  assign _GEN_2728 = 6'h26 == _T_294 ? welem[38] : _GEN_2727; // @[Execute.scala 117:10]
  assign _GEN_2729 = 6'h27 == _T_294 ? welem[39] : _GEN_2728; // @[Execute.scala 117:10]
  assign _GEN_2730 = 6'h28 == _T_294 ? welem[40] : _GEN_2729; // @[Execute.scala 117:10]
  assign _GEN_2731 = 6'h29 == _T_294 ? welem[41] : _GEN_2730; // @[Execute.scala 117:10]
  assign _GEN_2732 = 6'h2a == _T_294 ? welem[42] : _GEN_2731; // @[Execute.scala 117:10]
  assign _GEN_2733 = 6'h2b == _T_294 ? welem[43] : _GEN_2732; // @[Execute.scala 117:10]
  assign _GEN_2734 = 6'h2c == _T_294 ? welem[44] : _GEN_2733; // @[Execute.scala 117:10]
  assign _GEN_2735 = 6'h2d == _T_294 ? welem[45] : _GEN_2734; // @[Execute.scala 117:10]
  assign _GEN_2736 = 6'h2e == _T_294 ? welem[46] : _GEN_2735; // @[Execute.scala 117:10]
  assign _GEN_2737 = 6'h2f == _T_294 ? welem[47] : _GEN_2736; // @[Execute.scala 117:10]
  assign _GEN_2738 = 6'h30 == _T_294 ? welem[48] : _GEN_2737; // @[Execute.scala 117:10]
  assign _GEN_2739 = 6'h31 == _T_294 ? welem[49] : _GEN_2738; // @[Execute.scala 117:10]
  assign _GEN_2740 = 6'h32 == _T_294 ? welem[50] : _GEN_2739; // @[Execute.scala 117:10]
  assign _GEN_2741 = 6'h33 == _T_294 ? welem[51] : _GEN_2740; // @[Execute.scala 117:10]
  assign _GEN_2742 = 6'h34 == _T_294 ? welem[52] : _GEN_2741; // @[Execute.scala 117:10]
  assign _GEN_2743 = 6'h35 == _T_294 ? welem[53] : _GEN_2742; // @[Execute.scala 117:10]
  assign _GEN_2744 = 6'h36 == _T_294 ? welem[54] : _GEN_2743; // @[Execute.scala 117:10]
  assign _GEN_2745 = 6'h37 == _T_294 ? welem[55] : _GEN_2744; // @[Execute.scala 117:10]
  assign _GEN_2746 = 6'h38 == _T_294 ? welem[56] : _GEN_2745; // @[Execute.scala 117:10]
  assign _GEN_2747 = 6'h39 == _T_294 ? welem[57] : _GEN_2746; // @[Execute.scala 117:10]
  assign _GEN_2748 = 6'h3a == _T_294 ? welem[58] : _GEN_2747; // @[Execute.scala 117:10]
  assign _GEN_2749 = 6'h3b == _T_294 ? welem[59] : _GEN_2748; // @[Execute.scala 117:10]
  assign _GEN_2750 = 6'h3c == _T_294 ? welem[60] : _GEN_2749; // @[Execute.scala 117:10]
  assign _GEN_2751 = 6'h3d == _T_294 ? welem[61] : _GEN_2750; // @[Execute.scala 117:10]
  assign _GEN_2752 = 6'h3e == _T_294 ? welem[62] : _GEN_2751; // @[Execute.scala 117:10]
  assign _GEN_2753 = 6'h3f == _T_294 ? welem[63] : _GEN_2752; // @[Execute.scala 117:10]
  assign _GEN_2755 = 6'h1 == _T_298 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2756 = 6'h2 == _T_298 ? welem[2] : _GEN_2755; // @[Execute.scala 117:10]
  assign _GEN_2757 = 6'h3 == _T_298 ? welem[3] : _GEN_2756; // @[Execute.scala 117:10]
  assign _GEN_2758 = 6'h4 == _T_298 ? welem[4] : _GEN_2757; // @[Execute.scala 117:10]
  assign _GEN_2759 = 6'h5 == _T_298 ? welem[5] : _GEN_2758; // @[Execute.scala 117:10]
  assign _GEN_2760 = 6'h6 == _T_298 ? welem[6] : _GEN_2759; // @[Execute.scala 117:10]
  assign _GEN_2761 = 6'h7 == _T_298 ? welem[7] : _GEN_2760; // @[Execute.scala 117:10]
  assign _GEN_2762 = 6'h8 == _T_298 ? welem[8] : _GEN_2761; // @[Execute.scala 117:10]
  assign _GEN_2763 = 6'h9 == _T_298 ? welem[9] : _GEN_2762; // @[Execute.scala 117:10]
  assign _GEN_2764 = 6'ha == _T_298 ? welem[10] : _GEN_2763; // @[Execute.scala 117:10]
  assign _GEN_2765 = 6'hb == _T_298 ? welem[11] : _GEN_2764; // @[Execute.scala 117:10]
  assign _GEN_2766 = 6'hc == _T_298 ? welem[12] : _GEN_2765; // @[Execute.scala 117:10]
  assign _GEN_2767 = 6'hd == _T_298 ? welem[13] : _GEN_2766; // @[Execute.scala 117:10]
  assign _GEN_2768 = 6'he == _T_298 ? welem[14] : _GEN_2767; // @[Execute.scala 117:10]
  assign _GEN_2769 = 6'hf == _T_298 ? welem[15] : _GEN_2768; // @[Execute.scala 117:10]
  assign _GEN_2770 = 6'h10 == _T_298 ? welem[16] : _GEN_2769; // @[Execute.scala 117:10]
  assign _GEN_2771 = 6'h11 == _T_298 ? welem[17] : _GEN_2770; // @[Execute.scala 117:10]
  assign _GEN_2772 = 6'h12 == _T_298 ? welem[18] : _GEN_2771; // @[Execute.scala 117:10]
  assign _GEN_2773 = 6'h13 == _T_298 ? welem[19] : _GEN_2772; // @[Execute.scala 117:10]
  assign _GEN_2774 = 6'h14 == _T_298 ? welem[20] : _GEN_2773; // @[Execute.scala 117:10]
  assign _GEN_2775 = 6'h15 == _T_298 ? welem[21] : _GEN_2774; // @[Execute.scala 117:10]
  assign _GEN_2776 = 6'h16 == _T_298 ? welem[22] : _GEN_2775; // @[Execute.scala 117:10]
  assign _GEN_2777 = 6'h17 == _T_298 ? welem[23] : _GEN_2776; // @[Execute.scala 117:10]
  assign _GEN_2778 = 6'h18 == _T_298 ? welem[24] : _GEN_2777; // @[Execute.scala 117:10]
  assign _GEN_2779 = 6'h19 == _T_298 ? welem[25] : _GEN_2778; // @[Execute.scala 117:10]
  assign _GEN_2780 = 6'h1a == _T_298 ? welem[26] : _GEN_2779; // @[Execute.scala 117:10]
  assign _GEN_2781 = 6'h1b == _T_298 ? welem[27] : _GEN_2780; // @[Execute.scala 117:10]
  assign _GEN_2782 = 6'h1c == _T_298 ? welem[28] : _GEN_2781; // @[Execute.scala 117:10]
  assign _GEN_2783 = 6'h1d == _T_298 ? welem[29] : _GEN_2782; // @[Execute.scala 117:10]
  assign _GEN_2784 = 6'h1e == _T_298 ? welem[30] : _GEN_2783; // @[Execute.scala 117:10]
  assign _GEN_2785 = 6'h1f == _T_298 ? welem[31] : _GEN_2784; // @[Execute.scala 117:10]
  assign _GEN_2786 = 6'h20 == _T_298 ? welem[32] : _GEN_2785; // @[Execute.scala 117:10]
  assign _GEN_2787 = 6'h21 == _T_298 ? welem[33] : _GEN_2786; // @[Execute.scala 117:10]
  assign _GEN_2788 = 6'h22 == _T_298 ? welem[34] : _GEN_2787; // @[Execute.scala 117:10]
  assign _GEN_2789 = 6'h23 == _T_298 ? welem[35] : _GEN_2788; // @[Execute.scala 117:10]
  assign _GEN_2790 = 6'h24 == _T_298 ? welem[36] : _GEN_2789; // @[Execute.scala 117:10]
  assign _GEN_2791 = 6'h25 == _T_298 ? welem[37] : _GEN_2790; // @[Execute.scala 117:10]
  assign _GEN_2792 = 6'h26 == _T_298 ? welem[38] : _GEN_2791; // @[Execute.scala 117:10]
  assign _GEN_2793 = 6'h27 == _T_298 ? welem[39] : _GEN_2792; // @[Execute.scala 117:10]
  assign _GEN_2794 = 6'h28 == _T_298 ? welem[40] : _GEN_2793; // @[Execute.scala 117:10]
  assign _GEN_2795 = 6'h29 == _T_298 ? welem[41] : _GEN_2794; // @[Execute.scala 117:10]
  assign _GEN_2796 = 6'h2a == _T_298 ? welem[42] : _GEN_2795; // @[Execute.scala 117:10]
  assign _GEN_2797 = 6'h2b == _T_298 ? welem[43] : _GEN_2796; // @[Execute.scala 117:10]
  assign _GEN_2798 = 6'h2c == _T_298 ? welem[44] : _GEN_2797; // @[Execute.scala 117:10]
  assign _GEN_2799 = 6'h2d == _T_298 ? welem[45] : _GEN_2798; // @[Execute.scala 117:10]
  assign _GEN_2800 = 6'h2e == _T_298 ? welem[46] : _GEN_2799; // @[Execute.scala 117:10]
  assign _GEN_2801 = 6'h2f == _T_298 ? welem[47] : _GEN_2800; // @[Execute.scala 117:10]
  assign _GEN_2802 = 6'h30 == _T_298 ? welem[48] : _GEN_2801; // @[Execute.scala 117:10]
  assign _GEN_2803 = 6'h31 == _T_298 ? welem[49] : _GEN_2802; // @[Execute.scala 117:10]
  assign _GEN_2804 = 6'h32 == _T_298 ? welem[50] : _GEN_2803; // @[Execute.scala 117:10]
  assign _GEN_2805 = 6'h33 == _T_298 ? welem[51] : _GEN_2804; // @[Execute.scala 117:10]
  assign _GEN_2806 = 6'h34 == _T_298 ? welem[52] : _GEN_2805; // @[Execute.scala 117:10]
  assign _GEN_2807 = 6'h35 == _T_298 ? welem[53] : _GEN_2806; // @[Execute.scala 117:10]
  assign _GEN_2808 = 6'h36 == _T_298 ? welem[54] : _GEN_2807; // @[Execute.scala 117:10]
  assign _GEN_2809 = 6'h37 == _T_298 ? welem[55] : _GEN_2808; // @[Execute.scala 117:10]
  assign _GEN_2810 = 6'h38 == _T_298 ? welem[56] : _GEN_2809; // @[Execute.scala 117:10]
  assign _GEN_2811 = 6'h39 == _T_298 ? welem[57] : _GEN_2810; // @[Execute.scala 117:10]
  assign _GEN_2812 = 6'h3a == _T_298 ? welem[58] : _GEN_2811; // @[Execute.scala 117:10]
  assign _GEN_2813 = 6'h3b == _T_298 ? welem[59] : _GEN_2812; // @[Execute.scala 117:10]
  assign _GEN_2814 = 6'h3c == _T_298 ? welem[60] : _GEN_2813; // @[Execute.scala 117:10]
  assign _GEN_2815 = 6'h3d == _T_298 ? welem[61] : _GEN_2814; // @[Execute.scala 117:10]
  assign _GEN_2816 = 6'h3e == _T_298 ? welem[62] : _GEN_2815; // @[Execute.scala 117:10]
  assign _GEN_2817 = 6'h3f == _T_298 ? welem[63] : _GEN_2816; // @[Execute.scala 117:10]
  assign _T_301 = _T_292 ? _GEN_2753 : _GEN_2817; // @[Execute.scala 117:10]
  assign _T_302 = r < 6'h2b; // @[Execute.scala 117:15]
  assign _T_304 = r - 6'h2b; // @[Execute.scala 117:37]
  assign _T_308 = 6'h15 + r; // @[Execute.scala 117:60]
  assign _GEN_2819 = 6'h1 == _T_304 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2820 = 6'h2 == _T_304 ? welem[2] : _GEN_2819; // @[Execute.scala 117:10]
  assign _GEN_2821 = 6'h3 == _T_304 ? welem[3] : _GEN_2820; // @[Execute.scala 117:10]
  assign _GEN_2822 = 6'h4 == _T_304 ? welem[4] : _GEN_2821; // @[Execute.scala 117:10]
  assign _GEN_2823 = 6'h5 == _T_304 ? welem[5] : _GEN_2822; // @[Execute.scala 117:10]
  assign _GEN_2824 = 6'h6 == _T_304 ? welem[6] : _GEN_2823; // @[Execute.scala 117:10]
  assign _GEN_2825 = 6'h7 == _T_304 ? welem[7] : _GEN_2824; // @[Execute.scala 117:10]
  assign _GEN_2826 = 6'h8 == _T_304 ? welem[8] : _GEN_2825; // @[Execute.scala 117:10]
  assign _GEN_2827 = 6'h9 == _T_304 ? welem[9] : _GEN_2826; // @[Execute.scala 117:10]
  assign _GEN_2828 = 6'ha == _T_304 ? welem[10] : _GEN_2827; // @[Execute.scala 117:10]
  assign _GEN_2829 = 6'hb == _T_304 ? welem[11] : _GEN_2828; // @[Execute.scala 117:10]
  assign _GEN_2830 = 6'hc == _T_304 ? welem[12] : _GEN_2829; // @[Execute.scala 117:10]
  assign _GEN_2831 = 6'hd == _T_304 ? welem[13] : _GEN_2830; // @[Execute.scala 117:10]
  assign _GEN_2832 = 6'he == _T_304 ? welem[14] : _GEN_2831; // @[Execute.scala 117:10]
  assign _GEN_2833 = 6'hf == _T_304 ? welem[15] : _GEN_2832; // @[Execute.scala 117:10]
  assign _GEN_2834 = 6'h10 == _T_304 ? welem[16] : _GEN_2833; // @[Execute.scala 117:10]
  assign _GEN_2835 = 6'h11 == _T_304 ? welem[17] : _GEN_2834; // @[Execute.scala 117:10]
  assign _GEN_2836 = 6'h12 == _T_304 ? welem[18] : _GEN_2835; // @[Execute.scala 117:10]
  assign _GEN_2837 = 6'h13 == _T_304 ? welem[19] : _GEN_2836; // @[Execute.scala 117:10]
  assign _GEN_2838 = 6'h14 == _T_304 ? welem[20] : _GEN_2837; // @[Execute.scala 117:10]
  assign _GEN_2839 = 6'h15 == _T_304 ? welem[21] : _GEN_2838; // @[Execute.scala 117:10]
  assign _GEN_2840 = 6'h16 == _T_304 ? welem[22] : _GEN_2839; // @[Execute.scala 117:10]
  assign _GEN_2841 = 6'h17 == _T_304 ? welem[23] : _GEN_2840; // @[Execute.scala 117:10]
  assign _GEN_2842 = 6'h18 == _T_304 ? welem[24] : _GEN_2841; // @[Execute.scala 117:10]
  assign _GEN_2843 = 6'h19 == _T_304 ? welem[25] : _GEN_2842; // @[Execute.scala 117:10]
  assign _GEN_2844 = 6'h1a == _T_304 ? welem[26] : _GEN_2843; // @[Execute.scala 117:10]
  assign _GEN_2845 = 6'h1b == _T_304 ? welem[27] : _GEN_2844; // @[Execute.scala 117:10]
  assign _GEN_2846 = 6'h1c == _T_304 ? welem[28] : _GEN_2845; // @[Execute.scala 117:10]
  assign _GEN_2847 = 6'h1d == _T_304 ? welem[29] : _GEN_2846; // @[Execute.scala 117:10]
  assign _GEN_2848 = 6'h1e == _T_304 ? welem[30] : _GEN_2847; // @[Execute.scala 117:10]
  assign _GEN_2849 = 6'h1f == _T_304 ? welem[31] : _GEN_2848; // @[Execute.scala 117:10]
  assign _GEN_2850 = 6'h20 == _T_304 ? welem[32] : _GEN_2849; // @[Execute.scala 117:10]
  assign _GEN_2851 = 6'h21 == _T_304 ? welem[33] : _GEN_2850; // @[Execute.scala 117:10]
  assign _GEN_2852 = 6'h22 == _T_304 ? welem[34] : _GEN_2851; // @[Execute.scala 117:10]
  assign _GEN_2853 = 6'h23 == _T_304 ? welem[35] : _GEN_2852; // @[Execute.scala 117:10]
  assign _GEN_2854 = 6'h24 == _T_304 ? welem[36] : _GEN_2853; // @[Execute.scala 117:10]
  assign _GEN_2855 = 6'h25 == _T_304 ? welem[37] : _GEN_2854; // @[Execute.scala 117:10]
  assign _GEN_2856 = 6'h26 == _T_304 ? welem[38] : _GEN_2855; // @[Execute.scala 117:10]
  assign _GEN_2857 = 6'h27 == _T_304 ? welem[39] : _GEN_2856; // @[Execute.scala 117:10]
  assign _GEN_2858 = 6'h28 == _T_304 ? welem[40] : _GEN_2857; // @[Execute.scala 117:10]
  assign _GEN_2859 = 6'h29 == _T_304 ? welem[41] : _GEN_2858; // @[Execute.scala 117:10]
  assign _GEN_2860 = 6'h2a == _T_304 ? welem[42] : _GEN_2859; // @[Execute.scala 117:10]
  assign _GEN_2861 = 6'h2b == _T_304 ? welem[43] : _GEN_2860; // @[Execute.scala 117:10]
  assign _GEN_2862 = 6'h2c == _T_304 ? welem[44] : _GEN_2861; // @[Execute.scala 117:10]
  assign _GEN_2863 = 6'h2d == _T_304 ? welem[45] : _GEN_2862; // @[Execute.scala 117:10]
  assign _GEN_2864 = 6'h2e == _T_304 ? welem[46] : _GEN_2863; // @[Execute.scala 117:10]
  assign _GEN_2865 = 6'h2f == _T_304 ? welem[47] : _GEN_2864; // @[Execute.scala 117:10]
  assign _GEN_2866 = 6'h30 == _T_304 ? welem[48] : _GEN_2865; // @[Execute.scala 117:10]
  assign _GEN_2867 = 6'h31 == _T_304 ? welem[49] : _GEN_2866; // @[Execute.scala 117:10]
  assign _GEN_2868 = 6'h32 == _T_304 ? welem[50] : _GEN_2867; // @[Execute.scala 117:10]
  assign _GEN_2869 = 6'h33 == _T_304 ? welem[51] : _GEN_2868; // @[Execute.scala 117:10]
  assign _GEN_2870 = 6'h34 == _T_304 ? welem[52] : _GEN_2869; // @[Execute.scala 117:10]
  assign _GEN_2871 = 6'h35 == _T_304 ? welem[53] : _GEN_2870; // @[Execute.scala 117:10]
  assign _GEN_2872 = 6'h36 == _T_304 ? welem[54] : _GEN_2871; // @[Execute.scala 117:10]
  assign _GEN_2873 = 6'h37 == _T_304 ? welem[55] : _GEN_2872; // @[Execute.scala 117:10]
  assign _GEN_2874 = 6'h38 == _T_304 ? welem[56] : _GEN_2873; // @[Execute.scala 117:10]
  assign _GEN_2875 = 6'h39 == _T_304 ? welem[57] : _GEN_2874; // @[Execute.scala 117:10]
  assign _GEN_2876 = 6'h3a == _T_304 ? welem[58] : _GEN_2875; // @[Execute.scala 117:10]
  assign _GEN_2877 = 6'h3b == _T_304 ? welem[59] : _GEN_2876; // @[Execute.scala 117:10]
  assign _GEN_2878 = 6'h3c == _T_304 ? welem[60] : _GEN_2877; // @[Execute.scala 117:10]
  assign _GEN_2879 = 6'h3d == _T_304 ? welem[61] : _GEN_2878; // @[Execute.scala 117:10]
  assign _GEN_2880 = 6'h3e == _T_304 ? welem[62] : _GEN_2879; // @[Execute.scala 117:10]
  assign _GEN_2881 = 6'h3f == _T_304 ? welem[63] : _GEN_2880; // @[Execute.scala 117:10]
  assign _GEN_2883 = 6'h1 == _T_308 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2884 = 6'h2 == _T_308 ? welem[2] : _GEN_2883; // @[Execute.scala 117:10]
  assign _GEN_2885 = 6'h3 == _T_308 ? welem[3] : _GEN_2884; // @[Execute.scala 117:10]
  assign _GEN_2886 = 6'h4 == _T_308 ? welem[4] : _GEN_2885; // @[Execute.scala 117:10]
  assign _GEN_2887 = 6'h5 == _T_308 ? welem[5] : _GEN_2886; // @[Execute.scala 117:10]
  assign _GEN_2888 = 6'h6 == _T_308 ? welem[6] : _GEN_2887; // @[Execute.scala 117:10]
  assign _GEN_2889 = 6'h7 == _T_308 ? welem[7] : _GEN_2888; // @[Execute.scala 117:10]
  assign _GEN_2890 = 6'h8 == _T_308 ? welem[8] : _GEN_2889; // @[Execute.scala 117:10]
  assign _GEN_2891 = 6'h9 == _T_308 ? welem[9] : _GEN_2890; // @[Execute.scala 117:10]
  assign _GEN_2892 = 6'ha == _T_308 ? welem[10] : _GEN_2891; // @[Execute.scala 117:10]
  assign _GEN_2893 = 6'hb == _T_308 ? welem[11] : _GEN_2892; // @[Execute.scala 117:10]
  assign _GEN_2894 = 6'hc == _T_308 ? welem[12] : _GEN_2893; // @[Execute.scala 117:10]
  assign _GEN_2895 = 6'hd == _T_308 ? welem[13] : _GEN_2894; // @[Execute.scala 117:10]
  assign _GEN_2896 = 6'he == _T_308 ? welem[14] : _GEN_2895; // @[Execute.scala 117:10]
  assign _GEN_2897 = 6'hf == _T_308 ? welem[15] : _GEN_2896; // @[Execute.scala 117:10]
  assign _GEN_2898 = 6'h10 == _T_308 ? welem[16] : _GEN_2897; // @[Execute.scala 117:10]
  assign _GEN_2899 = 6'h11 == _T_308 ? welem[17] : _GEN_2898; // @[Execute.scala 117:10]
  assign _GEN_2900 = 6'h12 == _T_308 ? welem[18] : _GEN_2899; // @[Execute.scala 117:10]
  assign _GEN_2901 = 6'h13 == _T_308 ? welem[19] : _GEN_2900; // @[Execute.scala 117:10]
  assign _GEN_2902 = 6'h14 == _T_308 ? welem[20] : _GEN_2901; // @[Execute.scala 117:10]
  assign _GEN_2903 = 6'h15 == _T_308 ? welem[21] : _GEN_2902; // @[Execute.scala 117:10]
  assign _GEN_2904 = 6'h16 == _T_308 ? welem[22] : _GEN_2903; // @[Execute.scala 117:10]
  assign _GEN_2905 = 6'h17 == _T_308 ? welem[23] : _GEN_2904; // @[Execute.scala 117:10]
  assign _GEN_2906 = 6'h18 == _T_308 ? welem[24] : _GEN_2905; // @[Execute.scala 117:10]
  assign _GEN_2907 = 6'h19 == _T_308 ? welem[25] : _GEN_2906; // @[Execute.scala 117:10]
  assign _GEN_2908 = 6'h1a == _T_308 ? welem[26] : _GEN_2907; // @[Execute.scala 117:10]
  assign _GEN_2909 = 6'h1b == _T_308 ? welem[27] : _GEN_2908; // @[Execute.scala 117:10]
  assign _GEN_2910 = 6'h1c == _T_308 ? welem[28] : _GEN_2909; // @[Execute.scala 117:10]
  assign _GEN_2911 = 6'h1d == _T_308 ? welem[29] : _GEN_2910; // @[Execute.scala 117:10]
  assign _GEN_2912 = 6'h1e == _T_308 ? welem[30] : _GEN_2911; // @[Execute.scala 117:10]
  assign _GEN_2913 = 6'h1f == _T_308 ? welem[31] : _GEN_2912; // @[Execute.scala 117:10]
  assign _GEN_2914 = 6'h20 == _T_308 ? welem[32] : _GEN_2913; // @[Execute.scala 117:10]
  assign _GEN_2915 = 6'h21 == _T_308 ? welem[33] : _GEN_2914; // @[Execute.scala 117:10]
  assign _GEN_2916 = 6'h22 == _T_308 ? welem[34] : _GEN_2915; // @[Execute.scala 117:10]
  assign _GEN_2917 = 6'h23 == _T_308 ? welem[35] : _GEN_2916; // @[Execute.scala 117:10]
  assign _GEN_2918 = 6'h24 == _T_308 ? welem[36] : _GEN_2917; // @[Execute.scala 117:10]
  assign _GEN_2919 = 6'h25 == _T_308 ? welem[37] : _GEN_2918; // @[Execute.scala 117:10]
  assign _GEN_2920 = 6'h26 == _T_308 ? welem[38] : _GEN_2919; // @[Execute.scala 117:10]
  assign _GEN_2921 = 6'h27 == _T_308 ? welem[39] : _GEN_2920; // @[Execute.scala 117:10]
  assign _GEN_2922 = 6'h28 == _T_308 ? welem[40] : _GEN_2921; // @[Execute.scala 117:10]
  assign _GEN_2923 = 6'h29 == _T_308 ? welem[41] : _GEN_2922; // @[Execute.scala 117:10]
  assign _GEN_2924 = 6'h2a == _T_308 ? welem[42] : _GEN_2923; // @[Execute.scala 117:10]
  assign _GEN_2925 = 6'h2b == _T_308 ? welem[43] : _GEN_2924; // @[Execute.scala 117:10]
  assign _GEN_2926 = 6'h2c == _T_308 ? welem[44] : _GEN_2925; // @[Execute.scala 117:10]
  assign _GEN_2927 = 6'h2d == _T_308 ? welem[45] : _GEN_2926; // @[Execute.scala 117:10]
  assign _GEN_2928 = 6'h2e == _T_308 ? welem[46] : _GEN_2927; // @[Execute.scala 117:10]
  assign _GEN_2929 = 6'h2f == _T_308 ? welem[47] : _GEN_2928; // @[Execute.scala 117:10]
  assign _GEN_2930 = 6'h30 == _T_308 ? welem[48] : _GEN_2929; // @[Execute.scala 117:10]
  assign _GEN_2931 = 6'h31 == _T_308 ? welem[49] : _GEN_2930; // @[Execute.scala 117:10]
  assign _GEN_2932 = 6'h32 == _T_308 ? welem[50] : _GEN_2931; // @[Execute.scala 117:10]
  assign _GEN_2933 = 6'h33 == _T_308 ? welem[51] : _GEN_2932; // @[Execute.scala 117:10]
  assign _GEN_2934 = 6'h34 == _T_308 ? welem[52] : _GEN_2933; // @[Execute.scala 117:10]
  assign _GEN_2935 = 6'h35 == _T_308 ? welem[53] : _GEN_2934; // @[Execute.scala 117:10]
  assign _GEN_2936 = 6'h36 == _T_308 ? welem[54] : _GEN_2935; // @[Execute.scala 117:10]
  assign _GEN_2937 = 6'h37 == _T_308 ? welem[55] : _GEN_2936; // @[Execute.scala 117:10]
  assign _GEN_2938 = 6'h38 == _T_308 ? welem[56] : _GEN_2937; // @[Execute.scala 117:10]
  assign _GEN_2939 = 6'h39 == _T_308 ? welem[57] : _GEN_2938; // @[Execute.scala 117:10]
  assign _GEN_2940 = 6'h3a == _T_308 ? welem[58] : _GEN_2939; // @[Execute.scala 117:10]
  assign _GEN_2941 = 6'h3b == _T_308 ? welem[59] : _GEN_2940; // @[Execute.scala 117:10]
  assign _GEN_2942 = 6'h3c == _T_308 ? welem[60] : _GEN_2941; // @[Execute.scala 117:10]
  assign _GEN_2943 = 6'h3d == _T_308 ? welem[61] : _GEN_2942; // @[Execute.scala 117:10]
  assign _GEN_2944 = 6'h3e == _T_308 ? welem[62] : _GEN_2943; // @[Execute.scala 117:10]
  assign _GEN_2945 = 6'h3f == _T_308 ? welem[63] : _GEN_2944; // @[Execute.scala 117:10]
  assign _T_311 = _T_302 ? _GEN_2881 : _GEN_2945; // @[Execute.scala 117:10]
  assign _T_312 = r < 6'h2a; // @[Execute.scala 117:15]
  assign _T_314 = r - 6'h2a; // @[Execute.scala 117:37]
  assign _T_318 = 6'h16 + r; // @[Execute.scala 117:60]
  assign _GEN_2947 = 6'h1 == _T_314 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_2948 = 6'h2 == _T_314 ? welem[2] : _GEN_2947; // @[Execute.scala 117:10]
  assign _GEN_2949 = 6'h3 == _T_314 ? welem[3] : _GEN_2948; // @[Execute.scala 117:10]
  assign _GEN_2950 = 6'h4 == _T_314 ? welem[4] : _GEN_2949; // @[Execute.scala 117:10]
  assign _GEN_2951 = 6'h5 == _T_314 ? welem[5] : _GEN_2950; // @[Execute.scala 117:10]
  assign _GEN_2952 = 6'h6 == _T_314 ? welem[6] : _GEN_2951; // @[Execute.scala 117:10]
  assign _GEN_2953 = 6'h7 == _T_314 ? welem[7] : _GEN_2952; // @[Execute.scala 117:10]
  assign _GEN_2954 = 6'h8 == _T_314 ? welem[8] : _GEN_2953; // @[Execute.scala 117:10]
  assign _GEN_2955 = 6'h9 == _T_314 ? welem[9] : _GEN_2954; // @[Execute.scala 117:10]
  assign _GEN_2956 = 6'ha == _T_314 ? welem[10] : _GEN_2955; // @[Execute.scala 117:10]
  assign _GEN_2957 = 6'hb == _T_314 ? welem[11] : _GEN_2956; // @[Execute.scala 117:10]
  assign _GEN_2958 = 6'hc == _T_314 ? welem[12] : _GEN_2957; // @[Execute.scala 117:10]
  assign _GEN_2959 = 6'hd == _T_314 ? welem[13] : _GEN_2958; // @[Execute.scala 117:10]
  assign _GEN_2960 = 6'he == _T_314 ? welem[14] : _GEN_2959; // @[Execute.scala 117:10]
  assign _GEN_2961 = 6'hf == _T_314 ? welem[15] : _GEN_2960; // @[Execute.scala 117:10]
  assign _GEN_2962 = 6'h10 == _T_314 ? welem[16] : _GEN_2961; // @[Execute.scala 117:10]
  assign _GEN_2963 = 6'h11 == _T_314 ? welem[17] : _GEN_2962; // @[Execute.scala 117:10]
  assign _GEN_2964 = 6'h12 == _T_314 ? welem[18] : _GEN_2963; // @[Execute.scala 117:10]
  assign _GEN_2965 = 6'h13 == _T_314 ? welem[19] : _GEN_2964; // @[Execute.scala 117:10]
  assign _GEN_2966 = 6'h14 == _T_314 ? welem[20] : _GEN_2965; // @[Execute.scala 117:10]
  assign _GEN_2967 = 6'h15 == _T_314 ? welem[21] : _GEN_2966; // @[Execute.scala 117:10]
  assign _GEN_2968 = 6'h16 == _T_314 ? welem[22] : _GEN_2967; // @[Execute.scala 117:10]
  assign _GEN_2969 = 6'h17 == _T_314 ? welem[23] : _GEN_2968; // @[Execute.scala 117:10]
  assign _GEN_2970 = 6'h18 == _T_314 ? welem[24] : _GEN_2969; // @[Execute.scala 117:10]
  assign _GEN_2971 = 6'h19 == _T_314 ? welem[25] : _GEN_2970; // @[Execute.scala 117:10]
  assign _GEN_2972 = 6'h1a == _T_314 ? welem[26] : _GEN_2971; // @[Execute.scala 117:10]
  assign _GEN_2973 = 6'h1b == _T_314 ? welem[27] : _GEN_2972; // @[Execute.scala 117:10]
  assign _GEN_2974 = 6'h1c == _T_314 ? welem[28] : _GEN_2973; // @[Execute.scala 117:10]
  assign _GEN_2975 = 6'h1d == _T_314 ? welem[29] : _GEN_2974; // @[Execute.scala 117:10]
  assign _GEN_2976 = 6'h1e == _T_314 ? welem[30] : _GEN_2975; // @[Execute.scala 117:10]
  assign _GEN_2977 = 6'h1f == _T_314 ? welem[31] : _GEN_2976; // @[Execute.scala 117:10]
  assign _GEN_2978 = 6'h20 == _T_314 ? welem[32] : _GEN_2977; // @[Execute.scala 117:10]
  assign _GEN_2979 = 6'h21 == _T_314 ? welem[33] : _GEN_2978; // @[Execute.scala 117:10]
  assign _GEN_2980 = 6'h22 == _T_314 ? welem[34] : _GEN_2979; // @[Execute.scala 117:10]
  assign _GEN_2981 = 6'h23 == _T_314 ? welem[35] : _GEN_2980; // @[Execute.scala 117:10]
  assign _GEN_2982 = 6'h24 == _T_314 ? welem[36] : _GEN_2981; // @[Execute.scala 117:10]
  assign _GEN_2983 = 6'h25 == _T_314 ? welem[37] : _GEN_2982; // @[Execute.scala 117:10]
  assign _GEN_2984 = 6'h26 == _T_314 ? welem[38] : _GEN_2983; // @[Execute.scala 117:10]
  assign _GEN_2985 = 6'h27 == _T_314 ? welem[39] : _GEN_2984; // @[Execute.scala 117:10]
  assign _GEN_2986 = 6'h28 == _T_314 ? welem[40] : _GEN_2985; // @[Execute.scala 117:10]
  assign _GEN_2987 = 6'h29 == _T_314 ? welem[41] : _GEN_2986; // @[Execute.scala 117:10]
  assign _GEN_2988 = 6'h2a == _T_314 ? welem[42] : _GEN_2987; // @[Execute.scala 117:10]
  assign _GEN_2989 = 6'h2b == _T_314 ? welem[43] : _GEN_2988; // @[Execute.scala 117:10]
  assign _GEN_2990 = 6'h2c == _T_314 ? welem[44] : _GEN_2989; // @[Execute.scala 117:10]
  assign _GEN_2991 = 6'h2d == _T_314 ? welem[45] : _GEN_2990; // @[Execute.scala 117:10]
  assign _GEN_2992 = 6'h2e == _T_314 ? welem[46] : _GEN_2991; // @[Execute.scala 117:10]
  assign _GEN_2993 = 6'h2f == _T_314 ? welem[47] : _GEN_2992; // @[Execute.scala 117:10]
  assign _GEN_2994 = 6'h30 == _T_314 ? welem[48] : _GEN_2993; // @[Execute.scala 117:10]
  assign _GEN_2995 = 6'h31 == _T_314 ? welem[49] : _GEN_2994; // @[Execute.scala 117:10]
  assign _GEN_2996 = 6'h32 == _T_314 ? welem[50] : _GEN_2995; // @[Execute.scala 117:10]
  assign _GEN_2997 = 6'h33 == _T_314 ? welem[51] : _GEN_2996; // @[Execute.scala 117:10]
  assign _GEN_2998 = 6'h34 == _T_314 ? welem[52] : _GEN_2997; // @[Execute.scala 117:10]
  assign _GEN_2999 = 6'h35 == _T_314 ? welem[53] : _GEN_2998; // @[Execute.scala 117:10]
  assign _GEN_3000 = 6'h36 == _T_314 ? welem[54] : _GEN_2999; // @[Execute.scala 117:10]
  assign _GEN_3001 = 6'h37 == _T_314 ? welem[55] : _GEN_3000; // @[Execute.scala 117:10]
  assign _GEN_3002 = 6'h38 == _T_314 ? welem[56] : _GEN_3001; // @[Execute.scala 117:10]
  assign _GEN_3003 = 6'h39 == _T_314 ? welem[57] : _GEN_3002; // @[Execute.scala 117:10]
  assign _GEN_3004 = 6'h3a == _T_314 ? welem[58] : _GEN_3003; // @[Execute.scala 117:10]
  assign _GEN_3005 = 6'h3b == _T_314 ? welem[59] : _GEN_3004; // @[Execute.scala 117:10]
  assign _GEN_3006 = 6'h3c == _T_314 ? welem[60] : _GEN_3005; // @[Execute.scala 117:10]
  assign _GEN_3007 = 6'h3d == _T_314 ? welem[61] : _GEN_3006; // @[Execute.scala 117:10]
  assign _GEN_3008 = 6'h3e == _T_314 ? welem[62] : _GEN_3007; // @[Execute.scala 117:10]
  assign _GEN_3009 = 6'h3f == _T_314 ? welem[63] : _GEN_3008; // @[Execute.scala 117:10]
  assign _GEN_3011 = 6'h1 == _T_318 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3012 = 6'h2 == _T_318 ? welem[2] : _GEN_3011; // @[Execute.scala 117:10]
  assign _GEN_3013 = 6'h3 == _T_318 ? welem[3] : _GEN_3012; // @[Execute.scala 117:10]
  assign _GEN_3014 = 6'h4 == _T_318 ? welem[4] : _GEN_3013; // @[Execute.scala 117:10]
  assign _GEN_3015 = 6'h5 == _T_318 ? welem[5] : _GEN_3014; // @[Execute.scala 117:10]
  assign _GEN_3016 = 6'h6 == _T_318 ? welem[6] : _GEN_3015; // @[Execute.scala 117:10]
  assign _GEN_3017 = 6'h7 == _T_318 ? welem[7] : _GEN_3016; // @[Execute.scala 117:10]
  assign _GEN_3018 = 6'h8 == _T_318 ? welem[8] : _GEN_3017; // @[Execute.scala 117:10]
  assign _GEN_3019 = 6'h9 == _T_318 ? welem[9] : _GEN_3018; // @[Execute.scala 117:10]
  assign _GEN_3020 = 6'ha == _T_318 ? welem[10] : _GEN_3019; // @[Execute.scala 117:10]
  assign _GEN_3021 = 6'hb == _T_318 ? welem[11] : _GEN_3020; // @[Execute.scala 117:10]
  assign _GEN_3022 = 6'hc == _T_318 ? welem[12] : _GEN_3021; // @[Execute.scala 117:10]
  assign _GEN_3023 = 6'hd == _T_318 ? welem[13] : _GEN_3022; // @[Execute.scala 117:10]
  assign _GEN_3024 = 6'he == _T_318 ? welem[14] : _GEN_3023; // @[Execute.scala 117:10]
  assign _GEN_3025 = 6'hf == _T_318 ? welem[15] : _GEN_3024; // @[Execute.scala 117:10]
  assign _GEN_3026 = 6'h10 == _T_318 ? welem[16] : _GEN_3025; // @[Execute.scala 117:10]
  assign _GEN_3027 = 6'h11 == _T_318 ? welem[17] : _GEN_3026; // @[Execute.scala 117:10]
  assign _GEN_3028 = 6'h12 == _T_318 ? welem[18] : _GEN_3027; // @[Execute.scala 117:10]
  assign _GEN_3029 = 6'h13 == _T_318 ? welem[19] : _GEN_3028; // @[Execute.scala 117:10]
  assign _GEN_3030 = 6'h14 == _T_318 ? welem[20] : _GEN_3029; // @[Execute.scala 117:10]
  assign _GEN_3031 = 6'h15 == _T_318 ? welem[21] : _GEN_3030; // @[Execute.scala 117:10]
  assign _GEN_3032 = 6'h16 == _T_318 ? welem[22] : _GEN_3031; // @[Execute.scala 117:10]
  assign _GEN_3033 = 6'h17 == _T_318 ? welem[23] : _GEN_3032; // @[Execute.scala 117:10]
  assign _GEN_3034 = 6'h18 == _T_318 ? welem[24] : _GEN_3033; // @[Execute.scala 117:10]
  assign _GEN_3035 = 6'h19 == _T_318 ? welem[25] : _GEN_3034; // @[Execute.scala 117:10]
  assign _GEN_3036 = 6'h1a == _T_318 ? welem[26] : _GEN_3035; // @[Execute.scala 117:10]
  assign _GEN_3037 = 6'h1b == _T_318 ? welem[27] : _GEN_3036; // @[Execute.scala 117:10]
  assign _GEN_3038 = 6'h1c == _T_318 ? welem[28] : _GEN_3037; // @[Execute.scala 117:10]
  assign _GEN_3039 = 6'h1d == _T_318 ? welem[29] : _GEN_3038; // @[Execute.scala 117:10]
  assign _GEN_3040 = 6'h1e == _T_318 ? welem[30] : _GEN_3039; // @[Execute.scala 117:10]
  assign _GEN_3041 = 6'h1f == _T_318 ? welem[31] : _GEN_3040; // @[Execute.scala 117:10]
  assign _GEN_3042 = 6'h20 == _T_318 ? welem[32] : _GEN_3041; // @[Execute.scala 117:10]
  assign _GEN_3043 = 6'h21 == _T_318 ? welem[33] : _GEN_3042; // @[Execute.scala 117:10]
  assign _GEN_3044 = 6'h22 == _T_318 ? welem[34] : _GEN_3043; // @[Execute.scala 117:10]
  assign _GEN_3045 = 6'h23 == _T_318 ? welem[35] : _GEN_3044; // @[Execute.scala 117:10]
  assign _GEN_3046 = 6'h24 == _T_318 ? welem[36] : _GEN_3045; // @[Execute.scala 117:10]
  assign _GEN_3047 = 6'h25 == _T_318 ? welem[37] : _GEN_3046; // @[Execute.scala 117:10]
  assign _GEN_3048 = 6'h26 == _T_318 ? welem[38] : _GEN_3047; // @[Execute.scala 117:10]
  assign _GEN_3049 = 6'h27 == _T_318 ? welem[39] : _GEN_3048; // @[Execute.scala 117:10]
  assign _GEN_3050 = 6'h28 == _T_318 ? welem[40] : _GEN_3049; // @[Execute.scala 117:10]
  assign _GEN_3051 = 6'h29 == _T_318 ? welem[41] : _GEN_3050; // @[Execute.scala 117:10]
  assign _GEN_3052 = 6'h2a == _T_318 ? welem[42] : _GEN_3051; // @[Execute.scala 117:10]
  assign _GEN_3053 = 6'h2b == _T_318 ? welem[43] : _GEN_3052; // @[Execute.scala 117:10]
  assign _GEN_3054 = 6'h2c == _T_318 ? welem[44] : _GEN_3053; // @[Execute.scala 117:10]
  assign _GEN_3055 = 6'h2d == _T_318 ? welem[45] : _GEN_3054; // @[Execute.scala 117:10]
  assign _GEN_3056 = 6'h2e == _T_318 ? welem[46] : _GEN_3055; // @[Execute.scala 117:10]
  assign _GEN_3057 = 6'h2f == _T_318 ? welem[47] : _GEN_3056; // @[Execute.scala 117:10]
  assign _GEN_3058 = 6'h30 == _T_318 ? welem[48] : _GEN_3057; // @[Execute.scala 117:10]
  assign _GEN_3059 = 6'h31 == _T_318 ? welem[49] : _GEN_3058; // @[Execute.scala 117:10]
  assign _GEN_3060 = 6'h32 == _T_318 ? welem[50] : _GEN_3059; // @[Execute.scala 117:10]
  assign _GEN_3061 = 6'h33 == _T_318 ? welem[51] : _GEN_3060; // @[Execute.scala 117:10]
  assign _GEN_3062 = 6'h34 == _T_318 ? welem[52] : _GEN_3061; // @[Execute.scala 117:10]
  assign _GEN_3063 = 6'h35 == _T_318 ? welem[53] : _GEN_3062; // @[Execute.scala 117:10]
  assign _GEN_3064 = 6'h36 == _T_318 ? welem[54] : _GEN_3063; // @[Execute.scala 117:10]
  assign _GEN_3065 = 6'h37 == _T_318 ? welem[55] : _GEN_3064; // @[Execute.scala 117:10]
  assign _GEN_3066 = 6'h38 == _T_318 ? welem[56] : _GEN_3065; // @[Execute.scala 117:10]
  assign _GEN_3067 = 6'h39 == _T_318 ? welem[57] : _GEN_3066; // @[Execute.scala 117:10]
  assign _GEN_3068 = 6'h3a == _T_318 ? welem[58] : _GEN_3067; // @[Execute.scala 117:10]
  assign _GEN_3069 = 6'h3b == _T_318 ? welem[59] : _GEN_3068; // @[Execute.scala 117:10]
  assign _GEN_3070 = 6'h3c == _T_318 ? welem[60] : _GEN_3069; // @[Execute.scala 117:10]
  assign _GEN_3071 = 6'h3d == _T_318 ? welem[61] : _GEN_3070; // @[Execute.scala 117:10]
  assign _GEN_3072 = 6'h3e == _T_318 ? welem[62] : _GEN_3071; // @[Execute.scala 117:10]
  assign _GEN_3073 = 6'h3f == _T_318 ? welem[63] : _GEN_3072; // @[Execute.scala 117:10]
  assign _T_321 = _T_312 ? _GEN_3009 : _GEN_3073; // @[Execute.scala 117:10]
  assign _T_322 = r < 6'h29; // @[Execute.scala 117:15]
  assign _T_324 = r - 6'h29; // @[Execute.scala 117:37]
  assign _T_328 = 6'h17 + r; // @[Execute.scala 117:60]
  assign _GEN_3075 = 6'h1 == _T_324 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3076 = 6'h2 == _T_324 ? welem[2] : _GEN_3075; // @[Execute.scala 117:10]
  assign _GEN_3077 = 6'h3 == _T_324 ? welem[3] : _GEN_3076; // @[Execute.scala 117:10]
  assign _GEN_3078 = 6'h4 == _T_324 ? welem[4] : _GEN_3077; // @[Execute.scala 117:10]
  assign _GEN_3079 = 6'h5 == _T_324 ? welem[5] : _GEN_3078; // @[Execute.scala 117:10]
  assign _GEN_3080 = 6'h6 == _T_324 ? welem[6] : _GEN_3079; // @[Execute.scala 117:10]
  assign _GEN_3081 = 6'h7 == _T_324 ? welem[7] : _GEN_3080; // @[Execute.scala 117:10]
  assign _GEN_3082 = 6'h8 == _T_324 ? welem[8] : _GEN_3081; // @[Execute.scala 117:10]
  assign _GEN_3083 = 6'h9 == _T_324 ? welem[9] : _GEN_3082; // @[Execute.scala 117:10]
  assign _GEN_3084 = 6'ha == _T_324 ? welem[10] : _GEN_3083; // @[Execute.scala 117:10]
  assign _GEN_3085 = 6'hb == _T_324 ? welem[11] : _GEN_3084; // @[Execute.scala 117:10]
  assign _GEN_3086 = 6'hc == _T_324 ? welem[12] : _GEN_3085; // @[Execute.scala 117:10]
  assign _GEN_3087 = 6'hd == _T_324 ? welem[13] : _GEN_3086; // @[Execute.scala 117:10]
  assign _GEN_3088 = 6'he == _T_324 ? welem[14] : _GEN_3087; // @[Execute.scala 117:10]
  assign _GEN_3089 = 6'hf == _T_324 ? welem[15] : _GEN_3088; // @[Execute.scala 117:10]
  assign _GEN_3090 = 6'h10 == _T_324 ? welem[16] : _GEN_3089; // @[Execute.scala 117:10]
  assign _GEN_3091 = 6'h11 == _T_324 ? welem[17] : _GEN_3090; // @[Execute.scala 117:10]
  assign _GEN_3092 = 6'h12 == _T_324 ? welem[18] : _GEN_3091; // @[Execute.scala 117:10]
  assign _GEN_3093 = 6'h13 == _T_324 ? welem[19] : _GEN_3092; // @[Execute.scala 117:10]
  assign _GEN_3094 = 6'h14 == _T_324 ? welem[20] : _GEN_3093; // @[Execute.scala 117:10]
  assign _GEN_3095 = 6'h15 == _T_324 ? welem[21] : _GEN_3094; // @[Execute.scala 117:10]
  assign _GEN_3096 = 6'h16 == _T_324 ? welem[22] : _GEN_3095; // @[Execute.scala 117:10]
  assign _GEN_3097 = 6'h17 == _T_324 ? welem[23] : _GEN_3096; // @[Execute.scala 117:10]
  assign _GEN_3098 = 6'h18 == _T_324 ? welem[24] : _GEN_3097; // @[Execute.scala 117:10]
  assign _GEN_3099 = 6'h19 == _T_324 ? welem[25] : _GEN_3098; // @[Execute.scala 117:10]
  assign _GEN_3100 = 6'h1a == _T_324 ? welem[26] : _GEN_3099; // @[Execute.scala 117:10]
  assign _GEN_3101 = 6'h1b == _T_324 ? welem[27] : _GEN_3100; // @[Execute.scala 117:10]
  assign _GEN_3102 = 6'h1c == _T_324 ? welem[28] : _GEN_3101; // @[Execute.scala 117:10]
  assign _GEN_3103 = 6'h1d == _T_324 ? welem[29] : _GEN_3102; // @[Execute.scala 117:10]
  assign _GEN_3104 = 6'h1e == _T_324 ? welem[30] : _GEN_3103; // @[Execute.scala 117:10]
  assign _GEN_3105 = 6'h1f == _T_324 ? welem[31] : _GEN_3104; // @[Execute.scala 117:10]
  assign _GEN_3106 = 6'h20 == _T_324 ? welem[32] : _GEN_3105; // @[Execute.scala 117:10]
  assign _GEN_3107 = 6'h21 == _T_324 ? welem[33] : _GEN_3106; // @[Execute.scala 117:10]
  assign _GEN_3108 = 6'h22 == _T_324 ? welem[34] : _GEN_3107; // @[Execute.scala 117:10]
  assign _GEN_3109 = 6'h23 == _T_324 ? welem[35] : _GEN_3108; // @[Execute.scala 117:10]
  assign _GEN_3110 = 6'h24 == _T_324 ? welem[36] : _GEN_3109; // @[Execute.scala 117:10]
  assign _GEN_3111 = 6'h25 == _T_324 ? welem[37] : _GEN_3110; // @[Execute.scala 117:10]
  assign _GEN_3112 = 6'h26 == _T_324 ? welem[38] : _GEN_3111; // @[Execute.scala 117:10]
  assign _GEN_3113 = 6'h27 == _T_324 ? welem[39] : _GEN_3112; // @[Execute.scala 117:10]
  assign _GEN_3114 = 6'h28 == _T_324 ? welem[40] : _GEN_3113; // @[Execute.scala 117:10]
  assign _GEN_3115 = 6'h29 == _T_324 ? welem[41] : _GEN_3114; // @[Execute.scala 117:10]
  assign _GEN_3116 = 6'h2a == _T_324 ? welem[42] : _GEN_3115; // @[Execute.scala 117:10]
  assign _GEN_3117 = 6'h2b == _T_324 ? welem[43] : _GEN_3116; // @[Execute.scala 117:10]
  assign _GEN_3118 = 6'h2c == _T_324 ? welem[44] : _GEN_3117; // @[Execute.scala 117:10]
  assign _GEN_3119 = 6'h2d == _T_324 ? welem[45] : _GEN_3118; // @[Execute.scala 117:10]
  assign _GEN_3120 = 6'h2e == _T_324 ? welem[46] : _GEN_3119; // @[Execute.scala 117:10]
  assign _GEN_3121 = 6'h2f == _T_324 ? welem[47] : _GEN_3120; // @[Execute.scala 117:10]
  assign _GEN_3122 = 6'h30 == _T_324 ? welem[48] : _GEN_3121; // @[Execute.scala 117:10]
  assign _GEN_3123 = 6'h31 == _T_324 ? welem[49] : _GEN_3122; // @[Execute.scala 117:10]
  assign _GEN_3124 = 6'h32 == _T_324 ? welem[50] : _GEN_3123; // @[Execute.scala 117:10]
  assign _GEN_3125 = 6'h33 == _T_324 ? welem[51] : _GEN_3124; // @[Execute.scala 117:10]
  assign _GEN_3126 = 6'h34 == _T_324 ? welem[52] : _GEN_3125; // @[Execute.scala 117:10]
  assign _GEN_3127 = 6'h35 == _T_324 ? welem[53] : _GEN_3126; // @[Execute.scala 117:10]
  assign _GEN_3128 = 6'h36 == _T_324 ? welem[54] : _GEN_3127; // @[Execute.scala 117:10]
  assign _GEN_3129 = 6'h37 == _T_324 ? welem[55] : _GEN_3128; // @[Execute.scala 117:10]
  assign _GEN_3130 = 6'h38 == _T_324 ? welem[56] : _GEN_3129; // @[Execute.scala 117:10]
  assign _GEN_3131 = 6'h39 == _T_324 ? welem[57] : _GEN_3130; // @[Execute.scala 117:10]
  assign _GEN_3132 = 6'h3a == _T_324 ? welem[58] : _GEN_3131; // @[Execute.scala 117:10]
  assign _GEN_3133 = 6'h3b == _T_324 ? welem[59] : _GEN_3132; // @[Execute.scala 117:10]
  assign _GEN_3134 = 6'h3c == _T_324 ? welem[60] : _GEN_3133; // @[Execute.scala 117:10]
  assign _GEN_3135 = 6'h3d == _T_324 ? welem[61] : _GEN_3134; // @[Execute.scala 117:10]
  assign _GEN_3136 = 6'h3e == _T_324 ? welem[62] : _GEN_3135; // @[Execute.scala 117:10]
  assign _GEN_3137 = 6'h3f == _T_324 ? welem[63] : _GEN_3136; // @[Execute.scala 117:10]
  assign _GEN_3139 = 6'h1 == _T_328 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3140 = 6'h2 == _T_328 ? welem[2] : _GEN_3139; // @[Execute.scala 117:10]
  assign _GEN_3141 = 6'h3 == _T_328 ? welem[3] : _GEN_3140; // @[Execute.scala 117:10]
  assign _GEN_3142 = 6'h4 == _T_328 ? welem[4] : _GEN_3141; // @[Execute.scala 117:10]
  assign _GEN_3143 = 6'h5 == _T_328 ? welem[5] : _GEN_3142; // @[Execute.scala 117:10]
  assign _GEN_3144 = 6'h6 == _T_328 ? welem[6] : _GEN_3143; // @[Execute.scala 117:10]
  assign _GEN_3145 = 6'h7 == _T_328 ? welem[7] : _GEN_3144; // @[Execute.scala 117:10]
  assign _GEN_3146 = 6'h8 == _T_328 ? welem[8] : _GEN_3145; // @[Execute.scala 117:10]
  assign _GEN_3147 = 6'h9 == _T_328 ? welem[9] : _GEN_3146; // @[Execute.scala 117:10]
  assign _GEN_3148 = 6'ha == _T_328 ? welem[10] : _GEN_3147; // @[Execute.scala 117:10]
  assign _GEN_3149 = 6'hb == _T_328 ? welem[11] : _GEN_3148; // @[Execute.scala 117:10]
  assign _GEN_3150 = 6'hc == _T_328 ? welem[12] : _GEN_3149; // @[Execute.scala 117:10]
  assign _GEN_3151 = 6'hd == _T_328 ? welem[13] : _GEN_3150; // @[Execute.scala 117:10]
  assign _GEN_3152 = 6'he == _T_328 ? welem[14] : _GEN_3151; // @[Execute.scala 117:10]
  assign _GEN_3153 = 6'hf == _T_328 ? welem[15] : _GEN_3152; // @[Execute.scala 117:10]
  assign _GEN_3154 = 6'h10 == _T_328 ? welem[16] : _GEN_3153; // @[Execute.scala 117:10]
  assign _GEN_3155 = 6'h11 == _T_328 ? welem[17] : _GEN_3154; // @[Execute.scala 117:10]
  assign _GEN_3156 = 6'h12 == _T_328 ? welem[18] : _GEN_3155; // @[Execute.scala 117:10]
  assign _GEN_3157 = 6'h13 == _T_328 ? welem[19] : _GEN_3156; // @[Execute.scala 117:10]
  assign _GEN_3158 = 6'h14 == _T_328 ? welem[20] : _GEN_3157; // @[Execute.scala 117:10]
  assign _GEN_3159 = 6'h15 == _T_328 ? welem[21] : _GEN_3158; // @[Execute.scala 117:10]
  assign _GEN_3160 = 6'h16 == _T_328 ? welem[22] : _GEN_3159; // @[Execute.scala 117:10]
  assign _GEN_3161 = 6'h17 == _T_328 ? welem[23] : _GEN_3160; // @[Execute.scala 117:10]
  assign _GEN_3162 = 6'h18 == _T_328 ? welem[24] : _GEN_3161; // @[Execute.scala 117:10]
  assign _GEN_3163 = 6'h19 == _T_328 ? welem[25] : _GEN_3162; // @[Execute.scala 117:10]
  assign _GEN_3164 = 6'h1a == _T_328 ? welem[26] : _GEN_3163; // @[Execute.scala 117:10]
  assign _GEN_3165 = 6'h1b == _T_328 ? welem[27] : _GEN_3164; // @[Execute.scala 117:10]
  assign _GEN_3166 = 6'h1c == _T_328 ? welem[28] : _GEN_3165; // @[Execute.scala 117:10]
  assign _GEN_3167 = 6'h1d == _T_328 ? welem[29] : _GEN_3166; // @[Execute.scala 117:10]
  assign _GEN_3168 = 6'h1e == _T_328 ? welem[30] : _GEN_3167; // @[Execute.scala 117:10]
  assign _GEN_3169 = 6'h1f == _T_328 ? welem[31] : _GEN_3168; // @[Execute.scala 117:10]
  assign _GEN_3170 = 6'h20 == _T_328 ? welem[32] : _GEN_3169; // @[Execute.scala 117:10]
  assign _GEN_3171 = 6'h21 == _T_328 ? welem[33] : _GEN_3170; // @[Execute.scala 117:10]
  assign _GEN_3172 = 6'h22 == _T_328 ? welem[34] : _GEN_3171; // @[Execute.scala 117:10]
  assign _GEN_3173 = 6'h23 == _T_328 ? welem[35] : _GEN_3172; // @[Execute.scala 117:10]
  assign _GEN_3174 = 6'h24 == _T_328 ? welem[36] : _GEN_3173; // @[Execute.scala 117:10]
  assign _GEN_3175 = 6'h25 == _T_328 ? welem[37] : _GEN_3174; // @[Execute.scala 117:10]
  assign _GEN_3176 = 6'h26 == _T_328 ? welem[38] : _GEN_3175; // @[Execute.scala 117:10]
  assign _GEN_3177 = 6'h27 == _T_328 ? welem[39] : _GEN_3176; // @[Execute.scala 117:10]
  assign _GEN_3178 = 6'h28 == _T_328 ? welem[40] : _GEN_3177; // @[Execute.scala 117:10]
  assign _GEN_3179 = 6'h29 == _T_328 ? welem[41] : _GEN_3178; // @[Execute.scala 117:10]
  assign _GEN_3180 = 6'h2a == _T_328 ? welem[42] : _GEN_3179; // @[Execute.scala 117:10]
  assign _GEN_3181 = 6'h2b == _T_328 ? welem[43] : _GEN_3180; // @[Execute.scala 117:10]
  assign _GEN_3182 = 6'h2c == _T_328 ? welem[44] : _GEN_3181; // @[Execute.scala 117:10]
  assign _GEN_3183 = 6'h2d == _T_328 ? welem[45] : _GEN_3182; // @[Execute.scala 117:10]
  assign _GEN_3184 = 6'h2e == _T_328 ? welem[46] : _GEN_3183; // @[Execute.scala 117:10]
  assign _GEN_3185 = 6'h2f == _T_328 ? welem[47] : _GEN_3184; // @[Execute.scala 117:10]
  assign _GEN_3186 = 6'h30 == _T_328 ? welem[48] : _GEN_3185; // @[Execute.scala 117:10]
  assign _GEN_3187 = 6'h31 == _T_328 ? welem[49] : _GEN_3186; // @[Execute.scala 117:10]
  assign _GEN_3188 = 6'h32 == _T_328 ? welem[50] : _GEN_3187; // @[Execute.scala 117:10]
  assign _GEN_3189 = 6'h33 == _T_328 ? welem[51] : _GEN_3188; // @[Execute.scala 117:10]
  assign _GEN_3190 = 6'h34 == _T_328 ? welem[52] : _GEN_3189; // @[Execute.scala 117:10]
  assign _GEN_3191 = 6'h35 == _T_328 ? welem[53] : _GEN_3190; // @[Execute.scala 117:10]
  assign _GEN_3192 = 6'h36 == _T_328 ? welem[54] : _GEN_3191; // @[Execute.scala 117:10]
  assign _GEN_3193 = 6'h37 == _T_328 ? welem[55] : _GEN_3192; // @[Execute.scala 117:10]
  assign _GEN_3194 = 6'h38 == _T_328 ? welem[56] : _GEN_3193; // @[Execute.scala 117:10]
  assign _GEN_3195 = 6'h39 == _T_328 ? welem[57] : _GEN_3194; // @[Execute.scala 117:10]
  assign _GEN_3196 = 6'h3a == _T_328 ? welem[58] : _GEN_3195; // @[Execute.scala 117:10]
  assign _GEN_3197 = 6'h3b == _T_328 ? welem[59] : _GEN_3196; // @[Execute.scala 117:10]
  assign _GEN_3198 = 6'h3c == _T_328 ? welem[60] : _GEN_3197; // @[Execute.scala 117:10]
  assign _GEN_3199 = 6'h3d == _T_328 ? welem[61] : _GEN_3198; // @[Execute.scala 117:10]
  assign _GEN_3200 = 6'h3e == _T_328 ? welem[62] : _GEN_3199; // @[Execute.scala 117:10]
  assign _GEN_3201 = 6'h3f == _T_328 ? welem[63] : _GEN_3200; // @[Execute.scala 117:10]
  assign _T_331 = _T_322 ? _GEN_3137 : _GEN_3201; // @[Execute.scala 117:10]
  assign _T_332 = r < 6'h28; // @[Execute.scala 117:15]
  assign _T_334 = r - 6'h28; // @[Execute.scala 117:37]
  assign _T_338 = 6'h18 + r; // @[Execute.scala 117:60]
  assign _GEN_3203 = 6'h1 == _T_334 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3204 = 6'h2 == _T_334 ? welem[2] : _GEN_3203; // @[Execute.scala 117:10]
  assign _GEN_3205 = 6'h3 == _T_334 ? welem[3] : _GEN_3204; // @[Execute.scala 117:10]
  assign _GEN_3206 = 6'h4 == _T_334 ? welem[4] : _GEN_3205; // @[Execute.scala 117:10]
  assign _GEN_3207 = 6'h5 == _T_334 ? welem[5] : _GEN_3206; // @[Execute.scala 117:10]
  assign _GEN_3208 = 6'h6 == _T_334 ? welem[6] : _GEN_3207; // @[Execute.scala 117:10]
  assign _GEN_3209 = 6'h7 == _T_334 ? welem[7] : _GEN_3208; // @[Execute.scala 117:10]
  assign _GEN_3210 = 6'h8 == _T_334 ? welem[8] : _GEN_3209; // @[Execute.scala 117:10]
  assign _GEN_3211 = 6'h9 == _T_334 ? welem[9] : _GEN_3210; // @[Execute.scala 117:10]
  assign _GEN_3212 = 6'ha == _T_334 ? welem[10] : _GEN_3211; // @[Execute.scala 117:10]
  assign _GEN_3213 = 6'hb == _T_334 ? welem[11] : _GEN_3212; // @[Execute.scala 117:10]
  assign _GEN_3214 = 6'hc == _T_334 ? welem[12] : _GEN_3213; // @[Execute.scala 117:10]
  assign _GEN_3215 = 6'hd == _T_334 ? welem[13] : _GEN_3214; // @[Execute.scala 117:10]
  assign _GEN_3216 = 6'he == _T_334 ? welem[14] : _GEN_3215; // @[Execute.scala 117:10]
  assign _GEN_3217 = 6'hf == _T_334 ? welem[15] : _GEN_3216; // @[Execute.scala 117:10]
  assign _GEN_3218 = 6'h10 == _T_334 ? welem[16] : _GEN_3217; // @[Execute.scala 117:10]
  assign _GEN_3219 = 6'h11 == _T_334 ? welem[17] : _GEN_3218; // @[Execute.scala 117:10]
  assign _GEN_3220 = 6'h12 == _T_334 ? welem[18] : _GEN_3219; // @[Execute.scala 117:10]
  assign _GEN_3221 = 6'h13 == _T_334 ? welem[19] : _GEN_3220; // @[Execute.scala 117:10]
  assign _GEN_3222 = 6'h14 == _T_334 ? welem[20] : _GEN_3221; // @[Execute.scala 117:10]
  assign _GEN_3223 = 6'h15 == _T_334 ? welem[21] : _GEN_3222; // @[Execute.scala 117:10]
  assign _GEN_3224 = 6'h16 == _T_334 ? welem[22] : _GEN_3223; // @[Execute.scala 117:10]
  assign _GEN_3225 = 6'h17 == _T_334 ? welem[23] : _GEN_3224; // @[Execute.scala 117:10]
  assign _GEN_3226 = 6'h18 == _T_334 ? welem[24] : _GEN_3225; // @[Execute.scala 117:10]
  assign _GEN_3227 = 6'h19 == _T_334 ? welem[25] : _GEN_3226; // @[Execute.scala 117:10]
  assign _GEN_3228 = 6'h1a == _T_334 ? welem[26] : _GEN_3227; // @[Execute.scala 117:10]
  assign _GEN_3229 = 6'h1b == _T_334 ? welem[27] : _GEN_3228; // @[Execute.scala 117:10]
  assign _GEN_3230 = 6'h1c == _T_334 ? welem[28] : _GEN_3229; // @[Execute.scala 117:10]
  assign _GEN_3231 = 6'h1d == _T_334 ? welem[29] : _GEN_3230; // @[Execute.scala 117:10]
  assign _GEN_3232 = 6'h1e == _T_334 ? welem[30] : _GEN_3231; // @[Execute.scala 117:10]
  assign _GEN_3233 = 6'h1f == _T_334 ? welem[31] : _GEN_3232; // @[Execute.scala 117:10]
  assign _GEN_3234 = 6'h20 == _T_334 ? welem[32] : _GEN_3233; // @[Execute.scala 117:10]
  assign _GEN_3235 = 6'h21 == _T_334 ? welem[33] : _GEN_3234; // @[Execute.scala 117:10]
  assign _GEN_3236 = 6'h22 == _T_334 ? welem[34] : _GEN_3235; // @[Execute.scala 117:10]
  assign _GEN_3237 = 6'h23 == _T_334 ? welem[35] : _GEN_3236; // @[Execute.scala 117:10]
  assign _GEN_3238 = 6'h24 == _T_334 ? welem[36] : _GEN_3237; // @[Execute.scala 117:10]
  assign _GEN_3239 = 6'h25 == _T_334 ? welem[37] : _GEN_3238; // @[Execute.scala 117:10]
  assign _GEN_3240 = 6'h26 == _T_334 ? welem[38] : _GEN_3239; // @[Execute.scala 117:10]
  assign _GEN_3241 = 6'h27 == _T_334 ? welem[39] : _GEN_3240; // @[Execute.scala 117:10]
  assign _GEN_3242 = 6'h28 == _T_334 ? welem[40] : _GEN_3241; // @[Execute.scala 117:10]
  assign _GEN_3243 = 6'h29 == _T_334 ? welem[41] : _GEN_3242; // @[Execute.scala 117:10]
  assign _GEN_3244 = 6'h2a == _T_334 ? welem[42] : _GEN_3243; // @[Execute.scala 117:10]
  assign _GEN_3245 = 6'h2b == _T_334 ? welem[43] : _GEN_3244; // @[Execute.scala 117:10]
  assign _GEN_3246 = 6'h2c == _T_334 ? welem[44] : _GEN_3245; // @[Execute.scala 117:10]
  assign _GEN_3247 = 6'h2d == _T_334 ? welem[45] : _GEN_3246; // @[Execute.scala 117:10]
  assign _GEN_3248 = 6'h2e == _T_334 ? welem[46] : _GEN_3247; // @[Execute.scala 117:10]
  assign _GEN_3249 = 6'h2f == _T_334 ? welem[47] : _GEN_3248; // @[Execute.scala 117:10]
  assign _GEN_3250 = 6'h30 == _T_334 ? welem[48] : _GEN_3249; // @[Execute.scala 117:10]
  assign _GEN_3251 = 6'h31 == _T_334 ? welem[49] : _GEN_3250; // @[Execute.scala 117:10]
  assign _GEN_3252 = 6'h32 == _T_334 ? welem[50] : _GEN_3251; // @[Execute.scala 117:10]
  assign _GEN_3253 = 6'h33 == _T_334 ? welem[51] : _GEN_3252; // @[Execute.scala 117:10]
  assign _GEN_3254 = 6'h34 == _T_334 ? welem[52] : _GEN_3253; // @[Execute.scala 117:10]
  assign _GEN_3255 = 6'h35 == _T_334 ? welem[53] : _GEN_3254; // @[Execute.scala 117:10]
  assign _GEN_3256 = 6'h36 == _T_334 ? welem[54] : _GEN_3255; // @[Execute.scala 117:10]
  assign _GEN_3257 = 6'h37 == _T_334 ? welem[55] : _GEN_3256; // @[Execute.scala 117:10]
  assign _GEN_3258 = 6'h38 == _T_334 ? welem[56] : _GEN_3257; // @[Execute.scala 117:10]
  assign _GEN_3259 = 6'h39 == _T_334 ? welem[57] : _GEN_3258; // @[Execute.scala 117:10]
  assign _GEN_3260 = 6'h3a == _T_334 ? welem[58] : _GEN_3259; // @[Execute.scala 117:10]
  assign _GEN_3261 = 6'h3b == _T_334 ? welem[59] : _GEN_3260; // @[Execute.scala 117:10]
  assign _GEN_3262 = 6'h3c == _T_334 ? welem[60] : _GEN_3261; // @[Execute.scala 117:10]
  assign _GEN_3263 = 6'h3d == _T_334 ? welem[61] : _GEN_3262; // @[Execute.scala 117:10]
  assign _GEN_3264 = 6'h3e == _T_334 ? welem[62] : _GEN_3263; // @[Execute.scala 117:10]
  assign _GEN_3265 = 6'h3f == _T_334 ? welem[63] : _GEN_3264; // @[Execute.scala 117:10]
  assign _GEN_3267 = 6'h1 == _T_338 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3268 = 6'h2 == _T_338 ? welem[2] : _GEN_3267; // @[Execute.scala 117:10]
  assign _GEN_3269 = 6'h3 == _T_338 ? welem[3] : _GEN_3268; // @[Execute.scala 117:10]
  assign _GEN_3270 = 6'h4 == _T_338 ? welem[4] : _GEN_3269; // @[Execute.scala 117:10]
  assign _GEN_3271 = 6'h5 == _T_338 ? welem[5] : _GEN_3270; // @[Execute.scala 117:10]
  assign _GEN_3272 = 6'h6 == _T_338 ? welem[6] : _GEN_3271; // @[Execute.scala 117:10]
  assign _GEN_3273 = 6'h7 == _T_338 ? welem[7] : _GEN_3272; // @[Execute.scala 117:10]
  assign _GEN_3274 = 6'h8 == _T_338 ? welem[8] : _GEN_3273; // @[Execute.scala 117:10]
  assign _GEN_3275 = 6'h9 == _T_338 ? welem[9] : _GEN_3274; // @[Execute.scala 117:10]
  assign _GEN_3276 = 6'ha == _T_338 ? welem[10] : _GEN_3275; // @[Execute.scala 117:10]
  assign _GEN_3277 = 6'hb == _T_338 ? welem[11] : _GEN_3276; // @[Execute.scala 117:10]
  assign _GEN_3278 = 6'hc == _T_338 ? welem[12] : _GEN_3277; // @[Execute.scala 117:10]
  assign _GEN_3279 = 6'hd == _T_338 ? welem[13] : _GEN_3278; // @[Execute.scala 117:10]
  assign _GEN_3280 = 6'he == _T_338 ? welem[14] : _GEN_3279; // @[Execute.scala 117:10]
  assign _GEN_3281 = 6'hf == _T_338 ? welem[15] : _GEN_3280; // @[Execute.scala 117:10]
  assign _GEN_3282 = 6'h10 == _T_338 ? welem[16] : _GEN_3281; // @[Execute.scala 117:10]
  assign _GEN_3283 = 6'h11 == _T_338 ? welem[17] : _GEN_3282; // @[Execute.scala 117:10]
  assign _GEN_3284 = 6'h12 == _T_338 ? welem[18] : _GEN_3283; // @[Execute.scala 117:10]
  assign _GEN_3285 = 6'h13 == _T_338 ? welem[19] : _GEN_3284; // @[Execute.scala 117:10]
  assign _GEN_3286 = 6'h14 == _T_338 ? welem[20] : _GEN_3285; // @[Execute.scala 117:10]
  assign _GEN_3287 = 6'h15 == _T_338 ? welem[21] : _GEN_3286; // @[Execute.scala 117:10]
  assign _GEN_3288 = 6'h16 == _T_338 ? welem[22] : _GEN_3287; // @[Execute.scala 117:10]
  assign _GEN_3289 = 6'h17 == _T_338 ? welem[23] : _GEN_3288; // @[Execute.scala 117:10]
  assign _GEN_3290 = 6'h18 == _T_338 ? welem[24] : _GEN_3289; // @[Execute.scala 117:10]
  assign _GEN_3291 = 6'h19 == _T_338 ? welem[25] : _GEN_3290; // @[Execute.scala 117:10]
  assign _GEN_3292 = 6'h1a == _T_338 ? welem[26] : _GEN_3291; // @[Execute.scala 117:10]
  assign _GEN_3293 = 6'h1b == _T_338 ? welem[27] : _GEN_3292; // @[Execute.scala 117:10]
  assign _GEN_3294 = 6'h1c == _T_338 ? welem[28] : _GEN_3293; // @[Execute.scala 117:10]
  assign _GEN_3295 = 6'h1d == _T_338 ? welem[29] : _GEN_3294; // @[Execute.scala 117:10]
  assign _GEN_3296 = 6'h1e == _T_338 ? welem[30] : _GEN_3295; // @[Execute.scala 117:10]
  assign _GEN_3297 = 6'h1f == _T_338 ? welem[31] : _GEN_3296; // @[Execute.scala 117:10]
  assign _GEN_3298 = 6'h20 == _T_338 ? welem[32] : _GEN_3297; // @[Execute.scala 117:10]
  assign _GEN_3299 = 6'h21 == _T_338 ? welem[33] : _GEN_3298; // @[Execute.scala 117:10]
  assign _GEN_3300 = 6'h22 == _T_338 ? welem[34] : _GEN_3299; // @[Execute.scala 117:10]
  assign _GEN_3301 = 6'h23 == _T_338 ? welem[35] : _GEN_3300; // @[Execute.scala 117:10]
  assign _GEN_3302 = 6'h24 == _T_338 ? welem[36] : _GEN_3301; // @[Execute.scala 117:10]
  assign _GEN_3303 = 6'h25 == _T_338 ? welem[37] : _GEN_3302; // @[Execute.scala 117:10]
  assign _GEN_3304 = 6'h26 == _T_338 ? welem[38] : _GEN_3303; // @[Execute.scala 117:10]
  assign _GEN_3305 = 6'h27 == _T_338 ? welem[39] : _GEN_3304; // @[Execute.scala 117:10]
  assign _GEN_3306 = 6'h28 == _T_338 ? welem[40] : _GEN_3305; // @[Execute.scala 117:10]
  assign _GEN_3307 = 6'h29 == _T_338 ? welem[41] : _GEN_3306; // @[Execute.scala 117:10]
  assign _GEN_3308 = 6'h2a == _T_338 ? welem[42] : _GEN_3307; // @[Execute.scala 117:10]
  assign _GEN_3309 = 6'h2b == _T_338 ? welem[43] : _GEN_3308; // @[Execute.scala 117:10]
  assign _GEN_3310 = 6'h2c == _T_338 ? welem[44] : _GEN_3309; // @[Execute.scala 117:10]
  assign _GEN_3311 = 6'h2d == _T_338 ? welem[45] : _GEN_3310; // @[Execute.scala 117:10]
  assign _GEN_3312 = 6'h2e == _T_338 ? welem[46] : _GEN_3311; // @[Execute.scala 117:10]
  assign _GEN_3313 = 6'h2f == _T_338 ? welem[47] : _GEN_3312; // @[Execute.scala 117:10]
  assign _GEN_3314 = 6'h30 == _T_338 ? welem[48] : _GEN_3313; // @[Execute.scala 117:10]
  assign _GEN_3315 = 6'h31 == _T_338 ? welem[49] : _GEN_3314; // @[Execute.scala 117:10]
  assign _GEN_3316 = 6'h32 == _T_338 ? welem[50] : _GEN_3315; // @[Execute.scala 117:10]
  assign _GEN_3317 = 6'h33 == _T_338 ? welem[51] : _GEN_3316; // @[Execute.scala 117:10]
  assign _GEN_3318 = 6'h34 == _T_338 ? welem[52] : _GEN_3317; // @[Execute.scala 117:10]
  assign _GEN_3319 = 6'h35 == _T_338 ? welem[53] : _GEN_3318; // @[Execute.scala 117:10]
  assign _GEN_3320 = 6'h36 == _T_338 ? welem[54] : _GEN_3319; // @[Execute.scala 117:10]
  assign _GEN_3321 = 6'h37 == _T_338 ? welem[55] : _GEN_3320; // @[Execute.scala 117:10]
  assign _GEN_3322 = 6'h38 == _T_338 ? welem[56] : _GEN_3321; // @[Execute.scala 117:10]
  assign _GEN_3323 = 6'h39 == _T_338 ? welem[57] : _GEN_3322; // @[Execute.scala 117:10]
  assign _GEN_3324 = 6'h3a == _T_338 ? welem[58] : _GEN_3323; // @[Execute.scala 117:10]
  assign _GEN_3325 = 6'h3b == _T_338 ? welem[59] : _GEN_3324; // @[Execute.scala 117:10]
  assign _GEN_3326 = 6'h3c == _T_338 ? welem[60] : _GEN_3325; // @[Execute.scala 117:10]
  assign _GEN_3327 = 6'h3d == _T_338 ? welem[61] : _GEN_3326; // @[Execute.scala 117:10]
  assign _GEN_3328 = 6'h3e == _T_338 ? welem[62] : _GEN_3327; // @[Execute.scala 117:10]
  assign _GEN_3329 = 6'h3f == _T_338 ? welem[63] : _GEN_3328; // @[Execute.scala 117:10]
  assign _T_341 = _T_332 ? _GEN_3265 : _GEN_3329; // @[Execute.scala 117:10]
  assign _T_342 = r < 6'h27; // @[Execute.scala 117:15]
  assign _T_344 = r - 6'h27; // @[Execute.scala 117:37]
  assign _T_348 = 6'h19 + r; // @[Execute.scala 117:60]
  assign _GEN_3331 = 6'h1 == _T_344 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3332 = 6'h2 == _T_344 ? welem[2] : _GEN_3331; // @[Execute.scala 117:10]
  assign _GEN_3333 = 6'h3 == _T_344 ? welem[3] : _GEN_3332; // @[Execute.scala 117:10]
  assign _GEN_3334 = 6'h4 == _T_344 ? welem[4] : _GEN_3333; // @[Execute.scala 117:10]
  assign _GEN_3335 = 6'h5 == _T_344 ? welem[5] : _GEN_3334; // @[Execute.scala 117:10]
  assign _GEN_3336 = 6'h6 == _T_344 ? welem[6] : _GEN_3335; // @[Execute.scala 117:10]
  assign _GEN_3337 = 6'h7 == _T_344 ? welem[7] : _GEN_3336; // @[Execute.scala 117:10]
  assign _GEN_3338 = 6'h8 == _T_344 ? welem[8] : _GEN_3337; // @[Execute.scala 117:10]
  assign _GEN_3339 = 6'h9 == _T_344 ? welem[9] : _GEN_3338; // @[Execute.scala 117:10]
  assign _GEN_3340 = 6'ha == _T_344 ? welem[10] : _GEN_3339; // @[Execute.scala 117:10]
  assign _GEN_3341 = 6'hb == _T_344 ? welem[11] : _GEN_3340; // @[Execute.scala 117:10]
  assign _GEN_3342 = 6'hc == _T_344 ? welem[12] : _GEN_3341; // @[Execute.scala 117:10]
  assign _GEN_3343 = 6'hd == _T_344 ? welem[13] : _GEN_3342; // @[Execute.scala 117:10]
  assign _GEN_3344 = 6'he == _T_344 ? welem[14] : _GEN_3343; // @[Execute.scala 117:10]
  assign _GEN_3345 = 6'hf == _T_344 ? welem[15] : _GEN_3344; // @[Execute.scala 117:10]
  assign _GEN_3346 = 6'h10 == _T_344 ? welem[16] : _GEN_3345; // @[Execute.scala 117:10]
  assign _GEN_3347 = 6'h11 == _T_344 ? welem[17] : _GEN_3346; // @[Execute.scala 117:10]
  assign _GEN_3348 = 6'h12 == _T_344 ? welem[18] : _GEN_3347; // @[Execute.scala 117:10]
  assign _GEN_3349 = 6'h13 == _T_344 ? welem[19] : _GEN_3348; // @[Execute.scala 117:10]
  assign _GEN_3350 = 6'h14 == _T_344 ? welem[20] : _GEN_3349; // @[Execute.scala 117:10]
  assign _GEN_3351 = 6'h15 == _T_344 ? welem[21] : _GEN_3350; // @[Execute.scala 117:10]
  assign _GEN_3352 = 6'h16 == _T_344 ? welem[22] : _GEN_3351; // @[Execute.scala 117:10]
  assign _GEN_3353 = 6'h17 == _T_344 ? welem[23] : _GEN_3352; // @[Execute.scala 117:10]
  assign _GEN_3354 = 6'h18 == _T_344 ? welem[24] : _GEN_3353; // @[Execute.scala 117:10]
  assign _GEN_3355 = 6'h19 == _T_344 ? welem[25] : _GEN_3354; // @[Execute.scala 117:10]
  assign _GEN_3356 = 6'h1a == _T_344 ? welem[26] : _GEN_3355; // @[Execute.scala 117:10]
  assign _GEN_3357 = 6'h1b == _T_344 ? welem[27] : _GEN_3356; // @[Execute.scala 117:10]
  assign _GEN_3358 = 6'h1c == _T_344 ? welem[28] : _GEN_3357; // @[Execute.scala 117:10]
  assign _GEN_3359 = 6'h1d == _T_344 ? welem[29] : _GEN_3358; // @[Execute.scala 117:10]
  assign _GEN_3360 = 6'h1e == _T_344 ? welem[30] : _GEN_3359; // @[Execute.scala 117:10]
  assign _GEN_3361 = 6'h1f == _T_344 ? welem[31] : _GEN_3360; // @[Execute.scala 117:10]
  assign _GEN_3362 = 6'h20 == _T_344 ? welem[32] : _GEN_3361; // @[Execute.scala 117:10]
  assign _GEN_3363 = 6'h21 == _T_344 ? welem[33] : _GEN_3362; // @[Execute.scala 117:10]
  assign _GEN_3364 = 6'h22 == _T_344 ? welem[34] : _GEN_3363; // @[Execute.scala 117:10]
  assign _GEN_3365 = 6'h23 == _T_344 ? welem[35] : _GEN_3364; // @[Execute.scala 117:10]
  assign _GEN_3366 = 6'h24 == _T_344 ? welem[36] : _GEN_3365; // @[Execute.scala 117:10]
  assign _GEN_3367 = 6'h25 == _T_344 ? welem[37] : _GEN_3366; // @[Execute.scala 117:10]
  assign _GEN_3368 = 6'h26 == _T_344 ? welem[38] : _GEN_3367; // @[Execute.scala 117:10]
  assign _GEN_3369 = 6'h27 == _T_344 ? welem[39] : _GEN_3368; // @[Execute.scala 117:10]
  assign _GEN_3370 = 6'h28 == _T_344 ? welem[40] : _GEN_3369; // @[Execute.scala 117:10]
  assign _GEN_3371 = 6'h29 == _T_344 ? welem[41] : _GEN_3370; // @[Execute.scala 117:10]
  assign _GEN_3372 = 6'h2a == _T_344 ? welem[42] : _GEN_3371; // @[Execute.scala 117:10]
  assign _GEN_3373 = 6'h2b == _T_344 ? welem[43] : _GEN_3372; // @[Execute.scala 117:10]
  assign _GEN_3374 = 6'h2c == _T_344 ? welem[44] : _GEN_3373; // @[Execute.scala 117:10]
  assign _GEN_3375 = 6'h2d == _T_344 ? welem[45] : _GEN_3374; // @[Execute.scala 117:10]
  assign _GEN_3376 = 6'h2e == _T_344 ? welem[46] : _GEN_3375; // @[Execute.scala 117:10]
  assign _GEN_3377 = 6'h2f == _T_344 ? welem[47] : _GEN_3376; // @[Execute.scala 117:10]
  assign _GEN_3378 = 6'h30 == _T_344 ? welem[48] : _GEN_3377; // @[Execute.scala 117:10]
  assign _GEN_3379 = 6'h31 == _T_344 ? welem[49] : _GEN_3378; // @[Execute.scala 117:10]
  assign _GEN_3380 = 6'h32 == _T_344 ? welem[50] : _GEN_3379; // @[Execute.scala 117:10]
  assign _GEN_3381 = 6'h33 == _T_344 ? welem[51] : _GEN_3380; // @[Execute.scala 117:10]
  assign _GEN_3382 = 6'h34 == _T_344 ? welem[52] : _GEN_3381; // @[Execute.scala 117:10]
  assign _GEN_3383 = 6'h35 == _T_344 ? welem[53] : _GEN_3382; // @[Execute.scala 117:10]
  assign _GEN_3384 = 6'h36 == _T_344 ? welem[54] : _GEN_3383; // @[Execute.scala 117:10]
  assign _GEN_3385 = 6'h37 == _T_344 ? welem[55] : _GEN_3384; // @[Execute.scala 117:10]
  assign _GEN_3386 = 6'h38 == _T_344 ? welem[56] : _GEN_3385; // @[Execute.scala 117:10]
  assign _GEN_3387 = 6'h39 == _T_344 ? welem[57] : _GEN_3386; // @[Execute.scala 117:10]
  assign _GEN_3388 = 6'h3a == _T_344 ? welem[58] : _GEN_3387; // @[Execute.scala 117:10]
  assign _GEN_3389 = 6'h3b == _T_344 ? welem[59] : _GEN_3388; // @[Execute.scala 117:10]
  assign _GEN_3390 = 6'h3c == _T_344 ? welem[60] : _GEN_3389; // @[Execute.scala 117:10]
  assign _GEN_3391 = 6'h3d == _T_344 ? welem[61] : _GEN_3390; // @[Execute.scala 117:10]
  assign _GEN_3392 = 6'h3e == _T_344 ? welem[62] : _GEN_3391; // @[Execute.scala 117:10]
  assign _GEN_3393 = 6'h3f == _T_344 ? welem[63] : _GEN_3392; // @[Execute.scala 117:10]
  assign _GEN_3395 = 6'h1 == _T_348 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3396 = 6'h2 == _T_348 ? welem[2] : _GEN_3395; // @[Execute.scala 117:10]
  assign _GEN_3397 = 6'h3 == _T_348 ? welem[3] : _GEN_3396; // @[Execute.scala 117:10]
  assign _GEN_3398 = 6'h4 == _T_348 ? welem[4] : _GEN_3397; // @[Execute.scala 117:10]
  assign _GEN_3399 = 6'h5 == _T_348 ? welem[5] : _GEN_3398; // @[Execute.scala 117:10]
  assign _GEN_3400 = 6'h6 == _T_348 ? welem[6] : _GEN_3399; // @[Execute.scala 117:10]
  assign _GEN_3401 = 6'h7 == _T_348 ? welem[7] : _GEN_3400; // @[Execute.scala 117:10]
  assign _GEN_3402 = 6'h8 == _T_348 ? welem[8] : _GEN_3401; // @[Execute.scala 117:10]
  assign _GEN_3403 = 6'h9 == _T_348 ? welem[9] : _GEN_3402; // @[Execute.scala 117:10]
  assign _GEN_3404 = 6'ha == _T_348 ? welem[10] : _GEN_3403; // @[Execute.scala 117:10]
  assign _GEN_3405 = 6'hb == _T_348 ? welem[11] : _GEN_3404; // @[Execute.scala 117:10]
  assign _GEN_3406 = 6'hc == _T_348 ? welem[12] : _GEN_3405; // @[Execute.scala 117:10]
  assign _GEN_3407 = 6'hd == _T_348 ? welem[13] : _GEN_3406; // @[Execute.scala 117:10]
  assign _GEN_3408 = 6'he == _T_348 ? welem[14] : _GEN_3407; // @[Execute.scala 117:10]
  assign _GEN_3409 = 6'hf == _T_348 ? welem[15] : _GEN_3408; // @[Execute.scala 117:10]
  assign _GEN_3410 = 6'h10 == _T_348 ? welem[16] : _GEN_3409; // @[Execute.scala 117:10]
  assign _GEN_3411 = 6'h11 == _T_348 ? welem[17] : _GEN_3410; // @[Execute.scala 117:10]
  assign _GEN_3412 = 6'h12 == _T_348 ? welem[18] : _GEN_3411; // @[Execute.scala 117:10]
  assign _GEN_3413 = 6'h13 == _T_348 ? welem[19] : _GEN_3412; // @[Execute.scala 117:10]
  assign _GEN_3414 = 6'h14 == _T_348 ? welem[20] : _GEN_3413; // @[Execute.scala 117:10]
  assign _GEN_3415 = 6'h15 == _T_348 ? welem[21] : _GEN_3414; // @[Execute.scala 117:10]
  assign _GEN_3416 = 6'h16 == _T_348 ? welem[22] : _GEN_3415; // @[Execute.scala 117:10]
  assign _GEN_3417 = 6'h17 == _T_348 ? welem[23] : _GEN_3416; // @[Execute.scala 117:10]
  assign _GEN_3418 = 6'h18 == _T_348 ? welem[24] : _GEN_3417; // @[Execute.scala 117:10]
  assign _GEN_3419 = 6'h19 == _T_348 ? welem[25] : _GEN_3418; // @[Execute.scala 117:10]
  assign _GEN_3420 = 6'h1a == _T_348 ? welem[26] : _GEN_3419; // @[Execute.scala 117:10]
  assign _GEN_3421 = 6'h1b == _T_348 ? welem[27] : _GEN_3420; // @[Execute.scala 117:10]
  assign _GEN_3422 = 6'h1c == _T_348 ? welem[28] : _GEN_3421; // @[Execute.scala 117:10]
  assign _GEN_3423 = 6'h1d == _T_348 ? welem[29] : _GEN_3422; // @[Execute.scala 117:10]
  assign _GEN_3424 = 6'h1e == _T_348 ? welem[30] : _GEN_3423; // @[Execute.scala 117:10]
  assign _GEN_3425 = 6'h1f == _T_348 ? welem[31] : _GEN_3424; // @[Execute.scala 117:10]
  assign _GEN_3426 = 6'h20 == _T_348 ? welem[32] : _GEN_3425; // @[Execute.scala 117:10]
  assign _GEN_3427 = 6'h21 == _T_348 ? welem[33] : _GEN_3426; // @[Execute.scala 117:10]
  assign _GEN_3428 = 6'h22 == _T_348 ? welem[34] : _GEN_3427; // @[Execute.scala 117:10]
  assign _GEN_3429 = 6'h23 == _T_348 ? welem[35] : _GEN_3428; // @[Execute.scala 117:10]
  assign _GEN_3430 = 6'h24 == _T_348 ? welem[36] : _GEN_3429; // @[Execute.scala 117:10]
  assign _GEN_3431 = 6'h25 == _T_348 ? welem[37] : _GEN_3430; // @[Execute.scala 117:10]
  assign _GEN_3432 = 6'h26 == _T_348 ? welem[38] : _GEN_3431; // @[Execute.scala 117:10]
  assign _GEN_3433 = 6'h27 == _T_348 ? welem[39] : _GEN_3432; // @[Execute.scala 117:10]
  assign _GEN_3434 = 6'h28 == _T_348 ? welem[40] : _GEN_3433; // @[Execute.scala 117:10]
  assign _GEN_3435 = 6'h29 == _T_348 ? welem[41] : _GEN_3434; // @[Execute.scala 117:10]
  assign _GEN_3436 = 6'h2a == _T_348 ? welem[42] : _GEN_3435; // @[Execute.scala 117:10]
  assign _GEN_3437 = 6'h2b == _T_348 ? welem[43] : _GEN_3436; // @[Execute.scala 117:10]
  assign _GEN_3438 = 6'h2c == _T_348 ? welem[44] : _GEN_3437; // @[Execute.scala 117:10]
  assign _GEN_3439 = 6'h2d == _T_348 ? welem[45] : _GEN_3438; // @[Execute.scala 117:10]
  assign _GEN_3440 = 6'h2e == _T_348 ? welem[46] : _GEN_3439; // @[Execute.scala 117:10]
  assign _GEN_3441 = 6'h2f == _T_348 ? welem[47] : _GEN_3440; // @[Execute.scala 117:10]
  assign _GEN_3442 = 6'h30 == _T_348 ? welem[48] : _GEN_3441; // @[Execute.scala 117:10]
  assign _GEN_3443 = 6'h31 == _T_348 ? welem[49] : _GEN_3442; // @[Execute.scala 117:10]
  assign _GEN_3444 = 6'h32 == _T_348 ? welem[50] : _GEN_3443; // @[Execute.scala 117:10]
  assign _GEN_3445 = 6'h33 == _T_348 ? welem[51] : _GEN_3444; // @[Execute.scala 117:10]
  assign _GEN_3446 = 6'h34 == _T_348 ? welem[52] : _GEN_3445; // @[Execute.scala 117:10]
  assign _GEN_3447 = 6'h35 == _T_348 ? welem[53] : _GEN_3446; // @[Execute.scala 117:10]
  assign _GEN_3448 = 6'h36 == _T_348 ? welem[54] : _GEN_3447; // @[Execute.scala 117:10]
  assign _GEN_3449 = 6'h37 == _T_348 ? welem[55] : _GEN_3448; // @[Execute.scala 117:10]
  assign _GEN_3450 = 6'h38 == _T_348 ? welem[56] : _GEN_3449; // @[Execute.scala 117:10]
  assign _GEN_3451 = 6'h39 == _T_348 ? welem[57] : _GEN_3450; // @[Execute.scala 117:10]
  assign _GEN_3452 = 6'h3a == _T_348 ? welem[58] : _GEN_3451; // @[Execute.scala 117:10]
  assign _GEN_3453 = 6'h3b == _T_348 ? welem[59] : _GEN_3452; // @[Execute.scala 117:10]
  assign _GEN_3454 = 6'h3c == _T_348 ? welem[60] : _GEN_3453; // @[Execute.scala 117:10]
  assign _GEN_3455 = 6'h3d == _T_348 ? welem[61] : _GEN_3454; // @[Execute.scala 117:10]
  assign _GEN_3456 = 6'h3e == _T_348 ? welem[62] : _GEN_3455; // @[Execute.scala 117:10]
  assign _GEN_3457 = 6'h3f == _T_348 ? welem[63] : _GEN_3456; // @[Execute.scala 117:10]
  assign _T_351 = _T_342 ? _GEN_3393 : _GEN_3457; // @[Execute.scala 117:10]
  assign _T_352 = r < 6'h26; // @[Execute.scala 117:15]
  assign _T_354 = r - 6'h26; // @[Execute.scala 117:37]
  assign _T_358 = 6'h1a + r; // @[Execute.scala 117:60]
  assign _GEN_3459 = 6'h1 == _T_354 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3460 = 6'h2 == _T_354 ? welem[2] : _GEN_3459; // @[Execute.scala 117:10]
  assign _GEN_3461 = 6'h3 == _T_354 ? welem[3] : _GEN_3460; // @[Execute.scala 117:10]
  assign _GEN_3462 = 6'h4 == _T_354 ? welem[4] : _GEN_3461; // @[Execute.scala 117:10]
  assign _GEN_3463 = 6'h5 == _T_354 ? welem[5] : _GEN_3462; // @[Execute.scala 117:10]
  assign _GEN_3464 = 6'h6 == _T_354 ? welem[6] : _GEN_3463; // @[Execute.scala 117:10]
  assign _GEN_3465 = 6'h7 == _T_354 ? welem[7] : _GEN_3464; // @[Execute.scala 117:10]
  assign _GEN_3466 = 6'h8 == _T_354 ? welem[8] : _GEN_3465; // @[Execute.scala 117:10]
  assign _GEN_3467 = 6'h9 == _T_354 ? welem[9] : _GEN_3466; // @[Execute.scala 117:10]
  assign _GEN_3468 = 6'ha == _T_354 ? welem[10] : _GEN_3467; // @[Execute.scala 117:10]
  assign _GEN_3469 = 6'hb == _T_354 ? welem[11] : _GEN_3468; // @[Execute.scala 117:10]
  assign _GEN_3470 = 6'hc == _T_354 ? welem[12] : _GEN_3469; // @[Execute.scala 117:10]
  assign _GEN_3471 = 6'hd == _T_354 ? welem[13] : _GEN_3470; // @[Execute.scala 117:10]
  assign _GEN_3472 = 6'he == _T_354 ? welem[14] : _GEN_3471; // @[Execute.scala 117:10]
  assign _GEN_3473 = 6'hf == _T_354 ? welem[15] : _GEN_3472; // @[Execute.scala 117:10]
  assign _GEN_3474 = 6'h10 == _T_354 ? welem[16] : _GEN_3473; // @[Execute.scala 117:10]
  assign _GEN_3475 = 6'h11 == _T_354 ? welem[17] : _GEN_3474; // @[Execute.scala 117:10]
  assign _GEN_3476 = 6'h12 == _T_354 ? welem[18] : _GEN_3475; // @[Execute.scala 117:10]
  assign _GEN_3477 = 6'h13 == _T_354 ? welem[19] : _GEN_3476; // @[Execute.scala 117:10]
  assign _GEN_3478 = 6'h14 == _T_354 ? welem[20] : _GEN_3477; // @[Execute.scala 117:10]
  assign _GEN_3479 = 6'h15 == _T_354 ? welem[21] : _GEN_3478; // @[Execute.scala 117:10]
  assign _GEN_3480 = 6'h16 == _T_354 ? welem[22] : _GEN_3479; // @[Execute.scala 117:10]
  assign _GEN_3481 = 6'h17 == _T_354 ? welem[23] : _GEN_3480; // @[Execute.scala 117:10]
  assign _GEN_3482 = 6'h18 == _T_354 ? welem[24] : _GEN_3481; // @[Execute.scala 117:10]
  assign _GEN_3483 = 6'h19 == _T_354 ? welem[25] : _GEN_3482; // @[Execute.scala 117:10]
  assign _GEN_3484 = 6'h1a == _T_354 ? welem[26] : _GEN_3483; // @[Execute.scala 117:10]
  assign _GEN_3485 = 6'h1b == _T_354 ? welem[27] : _GEN_3484; // @[Execute.scala 117:10]
  assign _GEN_3486 = 6'h1c == _T_354 ? welem[28] : _GEN_3485; // @[Execute.scala 117:10]
  assign _GEN_3487 = 6'h1d == _T_354 ? welem[29] : _GEN_3486; // @[Execute.scala 117:10]
  assign _GEN_3488 = 6'h1e == _T_354 ? welem[30] : _GEN_3487; // @[Execute.scala 117:10]
  assign _GEN_3489 = 6'h1f == _T_354 ? welem[31] : _GEN_3488; // @[Execute.scala 117:10]
  assign _GEN_3490 = 6'h20 == _T_354 ? welem[32] : _GEN_3489; // @[Execute.scala 117:10]
  assign _GEN_3491 = 6'h21 == _T_354 ? welem[33] : _GEN_3490; // @[Execute.scala 117:10]
  assign _GEN_3492 = 6'h22 == _T_354 ? welem[34] : _GEN_3491; // @[Execute.scala 117:10]
  assign _GEN_3493 = 6'h23 == _T_354 ? welem[35] : _GEN_3492; // @[Execute.scala 117:10]
  assign _GEN_3494 = 6'h24 == _T_354 ? welem[36] : _GEN_3493; // @[Execute.scala 117:10]
  assign _GEN_3495 = 6'h25 == _T_354 ? welem[37] : _GEN_3494; // @[Execute.scala 117:10]
  assign _GEN_3496 = 6'h26 == _T_354 ? welem[38] : _GEN_3495; // @[Execute.scala 117:10]
  assign _GEN_3497 = 6'h27 == _T_354 ? welem[39] : _GEN_3496; // @[Execute.scala 117:10]
  assign _GEN_3498 = 6'h28 == _T_354 ? welem[40] : _GEN_3497; // @[Execute.scala 117:10]
  assign _GEN_3499 = 6'h29 == _T_354 ? welem[41] : _GEN_3498; // @[Execute.scala 117:10]
  assign _GEN_3500 = 6'h2a == _T_354 ? welem[42] : _GEN_3499; // @[Execute.scala 117:10]
  assign _GEN_3501 = 6'h2b == _T_354 ? welem[43] : _GEN_3500; // @[Execute.scala 117:10]
  assign _GEN_3502 = 6'h2c == _T_354 ? welem[44] : _GEN_3501; // @[Execute.scala 117:10]
  assign _GEN_3503 = 6'h2d == _T_354 ? welem[45] : _GEN_3502; // @[Execute.scala 117:10]
  assign _GEN_3504 = 6'h2e == _T_354 ? welem[46] : _GEN_3503; // @[Execute.scala 117:10]
  assign _GEN_3505 = 6'h2f == _T_354 ? welem[47] : _GEN_3504; // @[Execute.scala 117:10]
  assign _GEN_3506 = 6'h30 == _T_354 ? welem[48] : _GEN_3505; // @[Execute.scala 117:10]
  assign _GEN_3507 = 6'h31 == _T_354 ? welem[49] : _GEN_3506; // @[Execute.scala 117:10]
  assign _GEN_3508 = 6'h32 == _T_354 ? welem[50] : _GEN_3507; // @[Execute.scala 117:10]
  assign _GEN_3509 = 6'h33 == _T_354 ? welem[51] : _GEN_3508; // @[Execute.scala 117:10]
  assign _GEN_3510 = 6'h34 == _T_354 ? welem[52] : _GEN_3509; // @[Execute.scala 117:10]
  assign _GEN_3511 = 6'h35 == _T_354 ? welem[53] : _GEN_3510; // @[Execute.scala 117:10]
  assign _GEN_3512 = 6'h36 == _T_354 ? welem[54] : _GEN_3511; // @[Execute.scala 117:10]
  assign _GEN_3513 = 6'h37 == _T_354 ? welem[55] : _GEN_3512; // @[Execute.scala 117:10]
  assign _GEN_3514 = 6'h38 == _T_354 ? welem[56] : _GEN_3513; // @[Execute.scala 117:10]
  assign _GEN_3515 = 6'h39 == _T_354 ? welem[57] : _GEN_3514; // @[Execute.scala 117:10]
  assign _GEN_3516 = 6'h3a == _T_354 ? welem[58] : _GEN_3515; // @[Execute.scala 117:10]
  assign _GEN_3517 = 6'h3b == _T_354 ? welem[59] : _GEN_3516; // @[Execute.scala 117:10]
  assign _GEN_3518 = 6'h3c == _T_354 ? welem[60] : _GEN_3517; // @[Execute.scala 117:10]
  assign _GEN_3519 = 6'h3d == _T_354 ? welem[61] : _GEN_3518; // @[Execute.scala 117:10]
  assign _GEN_3520 = 6'h3e == _T_354 ? welem[62] : _GEN_3519; // @[Execute.scala 117:10]
  assign _GEN_3521 = 6'h3f == _T_354 ? welem[63] : _GEN_3520; // @[Execute.scala 117:10]
  assign _GEN_3523 = 6'h1 == _T_358 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3524 = 6'h2 == _T_358 ? welem[2] : _GEN_3523; // @[Execute.scala 117:10]
  assign _GEN_3525 = 6'h3 == _T_358 ? welem[3] : _GEN_3524; // @[Execute.scala 117:10]
  assign _GEN_3526 = 6'h4 == _T_358 ? welem[4] : _GEN_3525; // @[Execute.scala 117:10]
  assign _GEN_3527 = 6'h5 == _T_358 ? welem[5] : _GEN_3526; // @[Execute.scala 117:10]
  assign _GEN_3528 = 6'h6 == _T_358 ? welem[6] : _GEN_3527; // @[Execute.scala 117:10]
  assign _GEN_3529 = 6'h7 == _T_358 ? welem[7] : _GEN_3528; // @[Execute.scala 117:10]
  assign _GEN_3530 = 6'h8 == _T_358 ? welem[8] : _GEN_3529; // @[Execute.scala 117:10]
  assign _GEN_3531 = 6'h9 == _T_358 ? welem[9] : _GEN_3530; // @[Execute.scala 117:10]
  assign _GEN_3532 = 6'ha == _T_358 ? welem[10] : _GEN_3531; // @[Execute.scala 117:10]
  assign _GEN_3533 = 6'hb == _T_358 ? welem[11] : _GEN_3532; // @[Execute.scala 117:10]
  assign _GEN_3534 = 6'hc == _T_358 ? welem[12] : _GEN_3533; // @[Execute.scala 117:10]
  assign _GEN_3535 = 6'hd == _T_358 ? welem[13] : _GEN_3534; // @[Execute.scala 117:10]
  assign _GEN_3536 = 6'he == _T_358 ? welem[14] : _GEN_3535; // @[Execute.scala 117:10]
  assign _GEN_3537 = 6'hf == _T_358 ? welem[15] : _GEN_3536; // @[Execute.scala 117:10]
  assign _GEN_3538 = 6'h10 == _T_358 ? welem[16] : _GEN_3537; // @[Execute.scala 117:10]
  assign _GEN_3539 = 6'h11 == _T_358 ? welem[17] : _GEN_3538; // @[Execute.scala 117:10]
  assign _GEN_3540 = 6'h12 == _T_358 ? welem[18] : _GEN_3539; // @[Execute.scala 117:10]
  assign _GEN_3541 = 6'h13 == _T_358 ? welem[19] : _GEN_3540; // @[Execute.scala 117:10]
  assign _GEN_3542 = 6'h14 == _T_358 ? welem[20] : _GEN_3541; // @[Execute.scala 117:10]
  assign _GEN_3543 = 6'h15 == _T_358 ? welem[21] : _GEN_3542; // @[Execute.scala 117:10]
  assign _GEN_3544 = 6'h16 == _T_358 ? welem[22] : _GEN_3543; // @[Execute.scala 117:10]
  assign _GEN_3545 = 6'h17 == _T_358 ? welem[23] : _GEN_3544; // @[Execute.scala 117:10]
  assign _GEN_3546 = 6'h18 == _T_358 ? welem[24] : _GEN_3545; // @[Execute.scala 117:10]
  assign _GEN_3547 = 6'h19 == _T_358 ? welem[25] : _GEN_3546; // @[Execute.scala 117:10]
  assign _GEN_3548 = 6'h1a == _T_358 ? welem[26] : _GEN_3547; // @[Execute.scala 117:10]
  assign _GEN_3549 = 6'h1b == _T_358 ? welem[27] : _GEN_3548; // @[Execute.scala 117:10]
  assign _GEN_3550 = 6'h1c == _T_358 ? welem[28] : _GEN_3549; // @[Execute.scala 117:10]
  assign _GEN_3551 = 6'h1d == _T_358 ? welem[29] : _GEN_3550; // @[Execute.scala 117:10]
  assign _GEN_3552 = 6'h1e == _T_358 ? welem[30] : _GEN_3551; // @[Execute.scala 117:10]
  assign _GEN_3553 = 6'h1f == _T_358 ? welem[31] : _GEN_3552; // @[Execute.scala 117:10]
  assign _GEN_3554 = 6'h20 == _T_358 ? welem[32] : _GEN_3553; // @[Execute.scala 117:10]
  assign _GEN_3555 = 6'h21 == _T_358 ? welem[33] : _GEN_3554; // @[Execute.scala 117:10]
  assign _GEN_3556 = 6'h22 == _T_358 ? welem[34] : _GEN_3555; // @[Execute.scala 117:10]
  assign _GEN_3557 = 6'h23 == _T_358 ? welem[35] : _GEN_3556; // @[Execute.scala 117:10]
  assign _GEN_3558 = 6'h24 == _T_358 ? welem[36] : _GEN_3557; // @[Execute.scala 117:10]
  assign _GEN_3559 = 6'h25 == _T_358 ? welem[37] : _GEN_3558; // @[Execute.scala 117:10]
  assign _GEN_3560 = 6'h26 == _T_358 ? welem[38] : _GEN_3559; // @[Execute.scala 117:10]
  assign _GEN_3561 = 6'h27 == _T_358 ? welem[39] : _GEN_3560; // @[Execute.scala 117:10]
  assign _GEN_3562 = 6'h28 == _T_358 ? welem[40] : _GEN_3561; // @[Execute.scala 117:10]
  assign _GEN_3563 = 6'h29 == _T_358 ? welem[41] : _GEN_3562; // @[Execute.scala 117:10]
  assign _GEN_3564 = 6'h2a == _T_358 ? welem[42] : _GEN_3563; // @[Execute.scala 117:10]
  assign _GEN_3565 = 6'h2b == _T_358 ? welem[43] : _GEN_3564; // @[Execute.scala 117:10]
  assign _GEN_3566 = 6'h2c == _T_358 ? welem[44] : _GEN_3565; // @[Execute.scala 117:10]
  assign _GEN_3567 = 6'h2d == _T_358 ? welem[45] : _GEN_3566; // @[Execute.scala 117:10]
  assign _GEN_3568 = 6'h2e == _T_358 ? welem[46] : _GEN_3567; // @[Execute.scala 117:10]
  assign _GEN_3569 = 6'h2f == _T_358 ? welem[47] : _GEN_3568; // @[Execute.scala 117:10]
  assign _GEN_3570 = 6'h30 == _T_358 ? welem[48] : _GEN_3569; // @[Execute.scala 117:10]
  assign _GEN_3571 = 6'h31 == _T_358 ? welem[49] : _GEN_3570; // @[Execute.scala 117:10]
  assign _GEN_3572 = 6'h32 == _T_358 ? welem[50] : _GEN_3571; // @[Execute.scala 117:10]
  assign _GEN_3573 = 6'h33 == _T_358 ? welem[51] : _GEN_3572; // @[Execute.scala 117:10]
  assign _GEN_3574 = 6'h34 == _T_358 ? welem[52] : _GEN_3573; // @[Execute.scala 117:10]
  assign _GEN_3575 = 6'h35 == _T_358 ? welem[53] : _GEN_3574; // @[Execute.scala 117:10]
  assign _GEN_3576 = 6'h36 == _T_358 ? welem[54] : _GEN_3575; // @[Execute.scala 117:10]
  assign _GEN_3577 = 6'h37 == _T_358 ? welem[55] : _GEN_3576; // @[Execute.scala 117:10]
  assign _GEN_3578 = 6'h38 == _T_358 ? welem[56] : _GEN_3577; // @[Execute.scala 117:10]
  assign _GEN_3579 = 6'h39 == _T_358 ? welem[57] : _GEN_3578; // @[Execute.scala 117:10]
  assign _GEN_3580 = 6'h3a == _T_358 ? welem[58] : _GEN_3579; // @[Execute.scala 117:10]
  assign _GEN_3581 = 6'h3b == _T_358 ? welem[59] : _GEN_3580; // @[Execute.scala 117:10]
  assign _GEN_3582 = 6'h3c == _T_358 ? welem[60] : _GEN_3581; // @[Execute.scala 117:10]
  assign _GEN_3583 = 6'h3d == _T_358 ? welem[61] : _GEN_3582; // @[Execute.scala 117:10]
  assign _GEN_3584 = 6'h3e == _T_358 ? welem[62] : _GEN_3583; // @[Execute.scala 117:10]
  assign _GEN_3585 = 6'h3f == _T_358 ? welem[63] : _GEN_3584; // @[Execute.scala 117:10]
  assign _T_361 = _T_352 ? _GEN_3521 : _GEN_3585; // @[Execute.scala 117:10]
  assign _T_362 = r < 6'h25; // @[Execute.scala 117:15]
  assign _T_364 = r - 6'h25; // @[Execute.scala 117:37]
  assign _T_368 = 6'h1b + r; // @[Execute.scala 117:60]
  assign _GEN_3587 = 6'h1 == _T_364 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3588 = 6'h2 == _T_364 ? welem[2] : _GEN_3587; // @[Execute.scala 117:10]
  assign _GEN_3589 = 6'h3 == _T_364 ? welem[3] : _GEN_3588; // @[Execute.scala 117:10]
  assign _GEN_3590 = 6'h4 == _T_364 ? welem[4] : _GEN_3589; // @[Execute.scala 117:10]
  assign _GEN_3591 = 6'h5 == _T_364 ? welem[5] : _GEN_3590; // @[Execute.scala 117:10]
  assign _GEN_3592 = 6'h6 == _T_364 ? welem[6] : _GEN_3591; // @[Execute.scala 117:10]
  assign _GEN_3593 = 6'h7 == _T_364 ? welem[7] : _GEN_3592; // @[Execute.scala 117:10]
  assign _GEN_3594 = 6'h8 == _T_364 ? welem[8] : _GEN_3593; // @[Execute.scala 117:10]
  assign _GEN_3595 = 6'h9 == _T_364 ? welem[9] : _GEN_3594; // @[Execute.scala 117:10]
  assign _GEN_3596 = 6'ha == _T_364 ? welem[10] : _GEN_3595; // @[Execute.scala 117:10]
  assign _GEN_3597 = 6'hb == _T_364 ? welem[11] : _GEN_3596; // @[Execute.scala 117:10]
  assign _GEN_3598 = 6'hc == _T_364 ? welem[12] : _GEN_3597; // @[Execute.scala 117:10]
  assign _GEN_3599 = 6'hd == _T_364 ? welem[13] : _GEN_3598; // @[Execute.scala 117:10]
  assign _GEN_3600 = 6'he == _T_364 ? welem[14] : _GEN_3599; // @[Execute.scala 117:10]
  assign _GEN_3601 = 6'hf == _T_364 ? welem[15] : _GEN_3600; // @[Execute.scala 117:10]
  assign _GEN_3602 = 6'h10 == _T_364 ? welem[16] : _GEN_3601; // @[Execute.scala 117:10]
  assign _GEN_3603 = 6'h11 == _T_364 ? welem[17] : _GEN_3602; // @[Execute.scala 117:10]
  assign _GEN_3604 = 6'h12 == _T_364 ? welem[18] : _GEN_3603; // @[Execute.scala 117:10]
  assign _GEN_3605 = 6'h13 == _T_364 ? welem[19] : _GEN_3604; // @[Execute.scala 117:10]
  assign _GEN_3606 = 6'h14 == _T_364 ? welem[20] : _GEN_3605; // @[Execute.scala 117:10]
  assign _GEN_3607 = 6'h15 == _T_364 ? welem[21] : _GEN_3606; // @[Execute.scala 117:10]
  assign _GEN_3608 = 6'h16 == _T_364 ? welem[22] : _GEN_3607; // @[Execute.scala 117:10]
  assign _GEN_3609 = 6'h17 == _T_364 ? welem[23] : _GEN_3608; // @[Execute.scala 117:10]
  assign _GEN_3610 = 6'h18 == _T_364 ? welem[24] : _GEN_3609; // @[Execute.scala 117:10]
  assign _GEN_3611 = 6'h19 == _T_364 ? welem[25] : _GEN_3610; // @[Execute.scala 117:10]
  assign _GEN_3612 = 6'h1a == _T_364 ? welem[26] : _GEN_3611; // @[Execute.scala 117:10]
  assign _GEN_3613 = 6'h1b == _T_364 ? welem[27] : _GEN_3612; // @[Execute.scala 117:10]
  assign _GEN_3614 = 6'h1c == _T_364 ? welem[28] : _GEN_3613; // @[Execute.scala 117:10]
  assign _GEN_3615 = 6'h1d == _T_364 ? welem[29] : _GEN_3614; // @[Execute.scala 117:10]
  assign _GEN_3616 = 6'h1e == _T_364 ? welem[30] : _GEN_3615; // @[Execute.scala 117:10]
  assign _GEN_3617 = 6'h1f == _T_364 ? welem[31] : _GEN_3616; // @[Execute.scala 117:10]
  assign _GEN_3618 = 6'h20 == _T_364 ? welem[32] : _GEN_3617; // @[Execute.scala 117:10]
  assign _GEN_3619 = 6'h21 == _T_364 ? welem[33] : _GEN_3618; // @[Execute.scala 117:10]
  assign _GEN_3620 = 6'h22 == _T_364 ? welem[34] : _GEN_3619; // @[Execute.scala 117:10]
  assign _GEN_3621 = 6'h23 == _T_364 ? welem[35] : _GEN_3620; // @[Execute.scala 117:10]
  assign _GEN_3622 = 6'h24 == _T_364 ? welem[36] : _GEN_3621; // @[Execute.scala 117:10]
  assign _GEN_3623 = 6'h25 == _T_364 ? welem[37] : _GEN_3622; // @[Execute.scala 117:10]
  assign _GEN_3624 = 6'h26 == _T_364 ? welem[38] : _GEN_3623; // @[Execute.scala 117:10]
  assign _GEN_3625 = 6'h27 == _T_364 ? welem[39] : _GEN_3624; // @[Execute.scala 117:10]
  assign _GEN_3626 = 6'h28 == _T_364 ? welem[40] : _GEN_3625; // @[Execute.scala 117:10]
  assign _GEN_3627 = 6'h29 == _T_364 ? welem[41] : _GEN_3626; // @[Execute.scala 117:10]
  assign _GEN_3628 = 6'h2a == _T_364 ? welem[42] : _GEN_3627; // @[Execute.scala 117:10]
  assign _GEN_3629 = 6'h2b == _T_364 ? welem[43] : _GEN_3628; // @[Execute.scala 117:10]
  assign _GEN_3630 = 6'h2c == _T_364 ? welem[44] : _GEN_3629; // @[Execute.scala 117:10]
  assign _GEN_3631 = 6'h2d == _T_364 ? welem[45] : _GEN_3630; // @[Execute.scala 117:10]
  assign _GEN_3632 = 6'h2e == _T_364 ? welem[46] : _GEN_3631; // @[Execute.scala 117:10]
  assign _GEN_3633 = 6'h2f == _T_364 ? welem[47] : _GEN_3632; // @[Execute.scala 117:10]
  assign _GEN_3634 = 6'h30 == _T_364 ? welem[48] : _GEN_3633; // @[Execute.scala 117:10]
  assign _GEN_3635 = 6'h31 == _T_364 ? welem[49] : _GEN_3634; // @[Execute.scala 117:10]
  assign _GEN_3636 = 6'h32 == _T_364 ? welem[50] : _GEN_3635; // @[Execute.scala 117:10]
  assign _GEN_3637 = 6'h33 == _T_364 ? welem[51] : _GEN_3636; // @[Execute.scala 117:10]
  assign _GEN_3638 = 6'h34 == _T_364 ? welem[52] : _GEN_3637; // @[Execute.scala 117:10]
  assign _GEN_3639 = 6'h35 == _T_364 ? welem[53] : _GEN_3638; // @[Execute.scala 117:10]
  assign _GEN_3640 = 6'h36 == _T_364 ? welem[54] : _GEN_3639; // @[Execute.scala 117:10]
  assign _GEN_3641 = 6'h37 == _T_364 ? welem[55] : _GEN_3640; // @[Execute.scala 117:10]
  assign _GEN_3642 = 6'h38 == _T_364 ? welem[56] : _GEN_3641; // @[Execute.scala 117:10]
  assign _GEN_3643 = 6'h39 == _T_364 ? welem[57] : _GEN_3642; // @[Execute.scala 117:10]
  assign _GEN_3644 = 6'h3a == _T_364 ? welem[58] : _GEN_3643; // @[Execute.scala 117:10]
  assign _GEN_3645 = 6'h3b == _T_364 ? welem[59] : _GEN_3644; // @[Execute.scala 117:10]
  assign _GEN_3646 = 6'h3c == _T_364 ? welem[60] : _GEN_3645; // @[Execute.scala 117:10]
  assign _GEN_3647 = 6'h3d == _T_364 ? welem[61] : _GEN_3646; // @[Execute.scala 117:10]
  assign _GEN_3648 = 6'h3e == _T_364 ? welem[62] : _GEN_3647; // @[Execute.scala 117:10]
  assign _GEN_3649 = 6'h3f == _T_364 ? welem[63] : _GEN_3648; // @[Execute.scala 117:10]
  assign _GEN_3651 = 6'h1 == _T_368 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3652 = 6'h2 == _T_368 ? welem[2] : _GEN_3651; // @[Execute.scala 117:10]
  assign _GEN_3653 = 6'h3 == _T_368 ? welem[3] : _GEN_3652; // @[Execute.scala 117:10]
  assign _GEN_3654 = 6'h4 == _T_368 ? welem[4] : _GEN_3653; // @[Execute.scala 117:10]
  assign _GEN_3655 = 6'h5 == _T_368 ? welem[5] : _GEN_3654; // @[Execute.scala 117:10]
  assign _GEN_3656 = 6'h6 == _T_368 ? welem[6] : _GEN_3655; // @[Execute.scala 117:10]
  assign _GEN_3657 = 6'h7 == _T_368 ? welem[7] : _GEN_3656; // @[Execute.scala 117:10]
  assign _GEN_3658 = 6'h8 == _T_368 ? welem[8] : _GEN_3657; // @[Execute.scala 117:10]
  assign _GEN_3659 = 6'h9 == _T_368 ? welem[9] : _GEN_3658; // @[Execute.scala 117:10]
  assign _GEN_3660 = 6'ha == _T_368 ? welem[10] : _GEN_3659; // @[Execute.scala 117:10]
  assign _GEN_3661 = 6'hb == _T_368 ? welem[11] : _GEN_3660; // @[Execute.scala 117:10]
  assign _GEN_3662 = 6'hc == _T_368 ? welem[12] : _GEN_3661; // @[Execute.scala 117:10]
  assign _GEN_3663 = 6'hd == _T_368 ? welem[13] : _GEN_3662; // @[Execute.scala 117:10]
  assign _GEN_3664 = 6'he == _T_368 ? welem[14] : _GEN_3663; // @[Execute.scala 117:10]
  assign _GEN_3665 = 6'hf == _T_368 ? welem[15] : _GEN_3664; // @[Execute.scala 117:10]
  assign _GEN_3666 = 6'h10 == _T_368 ? welem[16] : _GEN_3665; // @[Execute.scala 117:10]
  assign _GEN_3667 = 6'h11 == _T_368 ? welem[17] : _GEN_3666; // @[Execute.scala 117:10]
  assign _GEN_3668 = 6'h12 == _T_368 ? welem[18] : _GEN_3667; // @[Execute.scala 117:10]
  assign _GEN_3669 = 6'h13 == _T_368 ? welem[19] : _GEN_3668; // @[Execute.scala 117:10]
  assign _GEN_3670 = 6'h14 == _T_368 ? welem[20] : _GEN_3669; // @[Execute.scala 117:10]
  assign _GEN_3671 = 6'h15 == _T_368 ? welem[21] : _GEN_3670; // @[Execute.scala 117:10]
  assign _GEN_3672 = 6'h16 == _T_368 ? welem[22] : _GEN_3671; // @[Execute.scala 117:10]
  assign _GEN_3673 = 6'h17 == _T_368 ? welem[23] : _GEN_3672; // @[Execute.scala 117:10]
  assign _GEN_3674 = 6'h18 == _T_368 ? welem[24] : _GEN_3673; // @[Execute.scala 117:10]
  assign _GEN_3675 = 6'h19 == _T_368 ? welem[25] : _GEN_3674; // @[Execute.scala 117:10]
  assign _GEN_3676 = 6'h1a == _T_368 ? welem[26] : _GEN_3675; // @[Execute.scala 117:10]
  assign _GEN_3677 = 6'h1b == _T_368 ? welem[27] : _GEN_3676; // @[Execute.scala 117:10]
  assign _GEN_3678 = 6'h1c == _T_368 ? welem[28] : _GEN_3677; // @[Execute.scala 117:10]
  assign _GEN_3679 = 6'h1d == _T_368 ? welem[29] : _GEN_3678; // @[Execute.scala 117:10]
  assign _GEN_3680 = 6'h1e == _T_368 ? welem[30] : _GEN_3679; // @[Execute.scala 117:10]
  assign _GEN_3681 = 6'h1f == _T_368 ? welem[31] : _GEN_3680; // @[Execute.scala 117:10]
  assign _GEN_3682 = 6'h20 == _T_368 ? welem[32] : _GEN_3681; // @[Execute.scala 117:10]
  assign _GEN_3683 = 6'h21 == _T_368 ? welem[33] : _GEN_3682; // @[Execute.scala 117:10]
  assign _GEN_3684 = 6'h22 == _T_368 ? welem[34] : _GEN_3683; // @[Execute.scala 117:10]
  assign _GEN_3685 = 6'h23 == _T_368 ? welem[35] : _GEN_3684; // @[Execute.scala 117:10]
  assign _GEN_3686 = 6'h24 == _T_368 ? welem[36] : _GEN_3685; // @[Execute.scala 117:10]
  assign _GEN_3687 = 6'h25 == _T_368 ? welem[37] : _GEN_3686; // @[Execute.scala 117:10]
  assign _GEN_3688 = 6'h26 == _T_368 ? welem[38] : _GEN_3687; // @[Execute.scala 117:10]
  assign _GEN_3689 = 6'h27 == _T_368 ? welem[39] : _GEN_3688; // @[Execute.scala 117:10]
  assign _GEN_3690 = 6'h28 == _T_368 ? welem[40] : _GEN_3689; // @[Execute.scala 117:10]
  assign _GEN_3691 = 6'h29 == _T_368 ? welem[41] : _GEN_3690; // @[Execute.scala 117:10]
  assign _GEN_3692 = 6'h2a == _T_368 ? welem[42] : _GEN_3691; // @[Execute.scala 117:10]
  assign _GEN_3693 = 6'h2b == _T_368 ? welem[43] : _GEN_3692; // @[Execute.scala 117:10]
  assign _GEN_3694 = 6'h2c == _T_368 ? welem[44] : _GEN_3693; // @[Execute.scala 117:10]
  assign _GEN_3695 = 6'h2d == _T_368 ? welem[45] : _GEN_3694; // @[Execute.scala 117:10]
  assign _GEN_3696 = 6'h2e == _T_368 ? welem[46] : _GEN_3695; // @[Execute.scala 117:10]
  assign _GEN_3697 = 6'h2f == _T_368 ? welem[47] : _GEN_3696; // @[Execute.scala 117:10]
  assign _GEN_3698 = 6'h30 == _T_368 ? welem[48] : _GEN_3697; // @[Execute.scala 117:10]
  assign _GEN_3699 = 6'h31 == _T_368 ? welem[49] : _GEN_3698; // @[Execute.scala 117:10]
  assign _GEN_3700 = 6'h32 == _T_368 ? welem[50] : _GEN_3699; // @[Execute.scala 117:10]
  assign _GEN_3701 = 6'h33 == _T_368 ? welem[51] : _GEN_3700; // @[Execute.scala 117:10]
  assign _GEN_3702 = 6'h34 == _T_368 ? welem[52] : _GEN_3701; // @[Execute.scala 117:10]
  assign _GEN_3703 = 6'h35 == _T_368 ? welem[53] : _GEN_3702; // @[Execute.scala 117:10]
  assign _GEN_3704 = 6'h36 == _T_368 ? welem[54] : _GEN_3703; // @[Execute.scala 117:10]
  assign _GEN_3705 = 6'h37 == _T_368 ? welem[55] : _GEN_3704; // @[Execute.scala 117:10]
  assign _GEN_3706 = 6'h38 == _T_368 ? welem[56] : _GEN_3705; // @[Execute.scala 117:10]
  assign _GEN_3707 = 6'h39 == _T_368 ? welem[57] : _GEN_3706; // @[Execute.scala 117:10]
  assign _GEN_3708 = 6'h3a == _T_368 ? welem[58] : _GEN_3707; // @[Execute.scala 117:10]
  assign _GEN_3709 = 6'h3b == _T_368 ? welem[59] : _GEN_3708; // @[Execute.scala 117:10]
  assign _GEN_3710 = 6'h3c == _T_368 ? welem[60] : _GEN_3709; // @[Execute.scala 117:10]
  assign _GEN_3711 = 6'h3d == _T_368 ? welem[61] : _GEN_3710; // @[Execute.scala 117:10]
  assign _GEN_3712 = 6'h3e == _T_368 ? welem[62] : _GEN_3711; // @[Execute.scala 117:10]
  assign _GEN_3713 = 6'h3f == _T_368 ? welem[63] : _GEN_3712; // @[Execute.scala 117:10]
  assign _T_371 = _T_362 ? _GEN_3649 : _GEN_3713; // @[Execute.scala 117:10]
  assign _T_372 = r < 6'h24; // @[Execute.scala 117:15]
  assign _T_374 = r - 6'h24; // @[Execute.scala 117:37]
  assign _T_378 = 6'h1c + r; // @[Execute.scala 117:60]
  assign _GEN_3715 = 6'h1 == _T_374 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3716 = 6'h2 == _T_374 ? welem[2] : _GEN_3715; // @[Execute.scala 117:10]
  assign _GEN_3717 = 6'h3 == _T_374 ? welem[3] : _GEN_3716; // @[Execute.scala 117:10]
  assign _GEN_3718 = 6'h4 == _T_374 ? welem[4] : _GEN_3717; // @[Execute.scala 117:10]
  assign _GEN_3719 = 6'h5 == _T_374 ? welem[5] : _GEN_3718; // @[Execute.scala 117:10]
  assign _GEN_3720 = 6'h6 == _T_374 ? welem[6] : _GEN_3719; // @[Execute.scala 117:10]
  assign _GEN_3721 = 6'h7 == _T_374 ? welem[7] : _GEN_3720; // @[Execute.scala 117:10]
  assign _GEN_3722 = 6'h8 == _T_374 ? welem[8] : _GEN_3721; // @[Execute.scala 117:10]
  assign _GEN_3723 = 6'h9 == _T_374 ? welem[9] : _GEN_3722; // @[Execute.scala 117:10]
  assign _GEN_3724 = 6'ha == _T_374 ? welem[10] : _GEN_3723; // @[Execute.scala 117:10]
  assign _GEN_3725 = 6'hb == _T_374 ? welem[11] : _GEN_3724; // @[Execute.scala 117:10]
  assign _GEN_3726 = 6'hc == _T_374 ? welem[12] : _GEN_3725; // @[Execute.scala 117:10]
  assign _GEN_3727 = 6'hd == _T_374 ? welem[13] : _GEN_3726; // @[Execute.scala 117:10]
  assign _GEN_3728 = 6'he == _T_374 ? welem[14] : _GEN_3727; // @[Execute.scala 117:10]
  assign _GEN_3729 = 6'hf == _T_374 ? welem[15] : _GEN_3728; // @[Execute.scala 117:10]
  assign _GEN_3730 = 6'h10 == _T_374 ? welem[16] : _GEN_3729; // @[Execute.scala 117:10]
  assign _GEN_3731 = 6'h11 == _T_374 ? welem[17] : _GEN_3730; // @[Execute.scala 117:10]
  assign _GEN_3732 = 6'h12 == _T_374 ? welem[18] : _GEN_3731; // @[Execute.scala 117:10]
  assign _GEN_3733 = 6'h13 == _T_374 ? welem[19] : _GEN_3732; // @[Execute.scala 117:10]
  assign _GEN_3734 = 6'h14 == _T_374 ? welem[20] : _GEN_3733; // @[Execute.scala 117:10]
  assign _GEN_3735 = 6'h15 == _T_374 ? welem[21] : _GEN_3734; // @[Execute.scala 117:10]
  assign _GEN_3736 = 6'h16 == _T_374 ? welem[22] : _GEN_3735; // @[Execute.scala 117:10]
  assign _GEN_3737 = 6'h17 == _T_374 ? welem[23] : _GEN_3736; // @[Execute.scala 117:10]
  assign _GEN_3738 = 6'h18 == _T_374 ? welem[24] : _GEN_3737; // @[Execute.scala 117:10]
  assign _GEN_3739 = 6'h19 == _T_374 ? welem[25] : _GEN_3738; // @[Execute.scala 117:10]
  assign _GEN_3740 = 6'h1a == _T_374 ? welem[26] : _GEN_3739; // @[Execute.scala 117:10]
  assign _GEN_3741 = 6'h1b == _T_374 ? welem[27] : _GEN_3740; // @[Execute.scala 117:10]
  assign _GEN_3742 = 6'h1c == _T_374 ? welem[28] : _GEN_3741; // @[Execute.scala 117:10]
  assign _GEN_3743 = 6'h1d == _T_374 ? welem[29] : _GEN_3742; // @[Execute.scala 117:10]
  assign _GEN_3744 = 6'h1e == _T_374 ? welem[30] : _GEN_3743; // @[Execute.scala 117:10]
  assign _GEN_3745 = 6'h1f == _T_374 ? welem[31] : _GEN_3744; // @[Execute.scala 117:10]
  assign _GEN_3746 = 6'h20 == _T_374 ? welem[32] : _GEN_3745; // @[Execute.scala 117:10]
  assign _GEN_3747 = 6'h21 == _T_374 ? welem[33] : _GEN_3746; // @[Execute.scala 117:10]
  assign _GEN_3748 = 6'h22 == _T_374 ? welem[34] : _GEN_3747; // @[Execute.scala 117:10]
  assign _GEN_3749 = 6'h23 == _T_374 ? welem[35] : _GEN_3748; // @[Execute.scala 117:10]
  assign _GEN_3750 = 6'h24 == _T_374 ? welem[36] : _GEN_3749; // @[Execute.scala 117:10]
  assign _GEN_3751 = 6'h25 == _T_374 ? welem[37] : _GEN_3750; // @[Execute.scala 117:10]
  assign _GEN_3752 = 6'h26 == _T_374 ? welem[38] : _GEN_3751; // @[Execute.scala 117:10]
  assign _GEN_3753 = 6'h27 == _T_374 ? welem[39] : _GEN_3752; // @[Execute.scala 117:10]
  assign _GEN_3754 = 6'h28 == _T_374 ? welem[40] : _GEN_3753; // @[Execute.scala 117:10]
  assign _GEN_3755 = 6'h29 == _T_374 ? welem[41] : _GEN_3754; // @[Execute.scala 117:10]
  assign _GEN_3756 = 6'h2a == _T_374 ? welem[42] : _GEN_3755; // @[Execute.scala 117:10]
  assign _GEN_3757 = 6'h2b == _T_374 ? welem[43] : _GEN_3756; // @[Execute.scala 117:10]
  assign _GEN_3758 = 6'h2c == _T_374 ? welem[44] : _GEN_3757; // @[Execute.scala 117:10]
  assign _GEN_3759 = 6'h2d == _T_374 ? welem[45] : _GEN_3758; // @[Execute.scala 117:10]
  assign _GEN_3760 = 6'h2e == _T_374 ? welem[46] : _GEN_3759; // @[Execute.scala 117:10]
  assign _GEN_3761 = 6'h2f == _T_374 ? welem[47] : _GEN_3760; // @[Execute.scala 117:10]
  assign _GEN_3762 = 6'h30 == _T_374 ? welem[48] : _GEN_3761; // @[Execute.scala 117:10]
  assign _GEN_3763 = 6'h31 == _T_374 ? welem[49] : _GEN_3762; // @[Execute.scala 117:10]
  assign _GEN_3764 = 6'h32 == _T_374 ? welem[50] : _GEN_3763; // @[Execute.scala 117:10]
  assign _GEN_3765 = 6'h33 == _T_374 ? welem[51] : _GEN_3764; // @[Execute.scala 117:10]
  assign _GEN_3766 = 6'h34 == _T_374 ? welem[52] : _GEN_3765; // @[Execute.scala 117:10]
  assign _GEN_3767 = 6'h35 == _T_374 ? welem[53] : _GEN_3766; // @[Execute.scala 117:10]
  assign _GEN_3768 = 6'h36 == _T_374 ? welem[54] : _GEN_3767; // @[Execute.scala 117:10]
  assign _GEN_3769 = 6'h37 == _T_374 ? welem[55] : _GEN_3768; // @[Execute.scala 117:10]
  assign _GEN_3770 = 6'h38 == _T_374 ? welem[56] : _GEN_3769; // @[Execute.scala 117:10]
  assign _GEN_3771 = 6'h39 == _T_374 ? welem[57] : _GEN_3770; // @[Execute.scala 117:10]
  assign _GEN_3772 = 6'h3a == _T_374 ? welem[58] : _GEN_3771; // @[Execute.scala 117:10]
  assign _GEN_3773 = 6'h3b == _T_374 ? welem[59] : _GEN_3772; // @[Execute.scala 117:10]
  assign _GEN_3774 = 6'h3c == _T_374 ? welem[60] : _GEN_3773; // @[Execute.scala 117:10]
  assign _GEN_3775 = 6'h3d == _T_374 ? welem[61] : _GEN_3774; // @[Execute.scala 117:10]
  assign _GEN_3776 = 6'h3e == _T_374 ? welem[62] : _GEN_3775; // @[Execute.scala 117:10]
  assign _GEN_3777 = 6'h3f == _T_374 ? welem[63] : _GEN_3776; // @[Execute.scala 117:10]
  assign _GEN_3779 = 6'h1 == _T_378 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3780 = 6'h2 == _T_378 ? welem[2] : _GEN_3779; // @[Execute.scala 117:10]
  assign _GEN_3781 = 6'h3 == _T_378 ? welem[3] : _GEN_3780; // @[Execute.scala 117:10]
  assign _GEN_3782 = 6'h4 == _T_378 ? welem[4] : _GEN_3781; // @[Execute.scala 117:10]
  assign _GEN_3783 = 6'h5 == _T_378 ? welem[5] : _GEN_3782; // @[Execute.scala 117:10]
  assign _GEN_3784 = 6'h6 == _T_378 ? welem[6] : _GEN_3783; // @[Execute.scala 117:10]
  assign _GEN_3785 = 6'h7 == _T_378 ? welem[7] : _GEN_3784; // @[Execute.scala 117:10]
  assign _GEN_3786 = 6'h8 == _T_378 ? welem[8] : _GEN_3785; // @[Execute.scala 117:10]
  assign _GEN_3787 = 6'h9 == _T_378 ? welem[9] : _GEN_3786; // @[Execute.scala 117:10]
  assign _GEN_3788 = 6'ha == _T_378 ? welem[10] : _GEN_3787; // @[Execute.scala 117:10]
  assign _GEN_3789 = 6'hb == _T_378 ? welem[11] : _GEN_3788; // @[Execute.scala 117:10]
  assign _GEN_3790 = 6'hc == _T_378 ? welem[12] : _GEN_3789; // @[Execute.scala 117:10]
  assign _GEN_3791 = 6'hd == _T_378 ? welem[13] : _GEN_3790; // @[Execute.scala 117:10]
  assign _GEN_3792 = 6'he == _T_378 ? welem[14] : _GEN_3791; // @[Execute.scala 117:10]
  assign _GEN_3793 = 6'hf == _T_378 ? welem[15] : _GEN_3792; // @[Execute.scala 117:10]
  assign _GEN_3794 = 6'h10 == _T_378 ? welem[16] : _GEN_3793; // @[Execute.scala 117:10]
  assign _GEN_3795 = 6'h11 == _T_378 ? welem[17] : _GEN_3794; // @[Execute.scala 117:10]
  assign _GEN_3796 = 6'h12 == _T_378 ? welem[18] : _GEN_3795; // @[Execute.scala 117:10]
  assign _GEN_3797 = 6'h13 == _T_378 ? welem[19] : _GEN_3796; // @[Execute.scala 117:10]
  assign _GEN_3798 = 6'h14 == _T_378 ? welem[20] : _GEN_3797; // @[Execute.scala 117:10]
  assign _GEN_3799 = 6'h15 == _T_378 ? welem[21] : _GEN_3798; // @[Execute.scala 117:10]
  assign _GEN_3800 = 6'h16 == _T_378 ? welem[22] : _GEN_3799; // @[Execute.scala 117:10]
  assign _GEN_3801 = 6'h17 == _T_378 ? welem[23] : _GEN_3800; // @[Execute.scala 117:10]
  assign _GEN_3802 = 6'h18 == _T_378 ? welem[24] : _GEN_3801; // @[Execute.scala 117:10]
  assign _GEN_3803 = 6'h19 == _T_378 ? welem[25] : _GEN_3802; // @[Execute.scala 117:10]
  assign _GEN_3804 = 6'h1a == _T_378 ? welem[26] : _GEN_3803; // @[Execute.scala 117:10]
  assign _GEN_3805 = 6'h1b == _T_378 ? welem[27] : _GEN_3804; // @[Execute.scala 117:10]
  assign _GEN_3806 = 6'h1c == _T_378 ? welem[28] : _GEN_3805; // @[Execute.scala 117:10]
  assign _GEN_3807 = 6'h1d == _T_378 ? welem[29] : _GEN_3806; // @[Execute.scala 117:10]
  assign _GEN_3808 = 6'h1e == _T_378 ? welem[30] : _GEN_3807; // @[Execute.scala 117:10]
  assign _GEN_3809 = 6'h1f == _T_378 ? welem[31] : _GEN_3808; // @[Execute.scala 117:10]
  assign _GEN_3810 = 6'h20 == _T_378 ? welem[32] : _GEN_3809; // @[Execute.scala 117:10]
  assign _GEN_3811 = 6'h21 == _T_378 ? welem[33] : _GEN_3810; // @[Execute.scala 117:10]
  assign _GEN_3812 = 6'h22 == _T_378 ? welem[34] : _GEN_3811; // @[Execute.scala 117:10]
  assign _GEN_3813 = 6'h23 == _T_378 ? welem[35] : _GEN_3812; // @[Execute.scala 117:10]
  assign _GEN_3814 = 6'h24 == _T_378 ? welem[36] : _GEN_3813; // @[Execute.scala 117:10]
  assign _GEN_3815 = 6'h25 == _T_378 ? welem[37] : _GEN_3814; // @[Execute.scala 117:10]
  assign _GEN_3816 = 6'h26 == _T_378 ? welem[38] : _GEN_3815; // @[Execute.scala 117:10]
  assign _GEN_3817 = 6'h27 == _T_378 ? welem[39] : _GEN_3816; // @[Execute.scala 117:10]
  assign _GEN_3818 = 6'h28 == _T_378 ? welem[40] : _GEN_3817; // @[Execute.scala 117:10]
  assign _GEN_3819 = 6'h29 == _T_378 ? welem[41] : _GEN_3818; // @[Execute.scala 117:10]
  assign _GEN_3820 = 6'h2a == _T_378 ? welem[42] : _GEN_3819; // @[Execute.scala 117:10]
  assign _GEN_3821 = 6'h2b == _T_378 ? welem[43] : _GEN_3820; // @[Execute.scala 117:10]
  assign _GEN_3822 = 6'h2c == _T_378 ? welem[44] : _GEN_3821; // @[Execute.scala 117:10]
  assign _GEN_3823 = 6'h2d == _T_378 ? welem[45] : _GEN_3822; // @[Execute.scala 117:10]
  assign _GEN_3824 = 6'h2e == _T_378 ? welem[46] : _GEN_3823; // @[Execute.scala 117:10]
  assign _GEN_3825 = 6'h2f == _T_378 ? welem[47] : _GEN_3824; // @[Execute.scala 117:10]
  assign _GEN_3826 = 6'h30 == _T_378 ? welem[48] : _GEN_3825; // @[Execute.scala 117:10]
  assign _GEN_3827 = 6'h31 == _T_378 ? welem[49] : _GEN_3826; // @[Execute.scala 117:10]
  assign _GEN_3828 = 6'h32 == _T_378 ? welem[50] : _GEN_3827; // @[Execute.scala 117:10]
  assign _GEN_3829 = 6'h33 == _T_378 ? welem[51] : _GEN_3828; // @[Execute.scala 117:10]
  assign _GEN_3830 = 6'h34 == _T_378 ? welem[52] : _GEN_3829; // @[Execute.scala 117:10]
  assign _GEN_3831 = 6'h35 == _T_378 ? welem[53] : _GEN_3830; // @[Execute.scala 117:10]
  assign _GEN_3832 = 6'h36 == _T_378 ? welem[54] : _GEN_3831; // @[Execute.scala 117:10]
  assign _GEN_3833 = 6'h37 == _T_378 ? welem[55] : _GEN_3832; // @[Execute.scala 117:10]
  assign _GEN_3834 = 6'h38 == _T_378 ? welem[56] : _GEN_3833; // @[Execute.scala 117:10]
  assign _GEN_3835 = 6'h39 == _T_378 ? welem[57] : _GEN_3834; // @[Execute.scala 117:10]
  assign _GEN_3836 = 6'h3a == _T_378 ? welem[58] : _GEN_3835; // @[Execute.scala 117:10]
  assign _GEN_3837 = 6'h3b == _T_378 ? welem[59] : _GEN_3836; // @[Execute.scala 117:10]
  assign _GEN_3838 = 6'h3c == _T_378 ? welem[60] : _GEN_3837; // @[Execute.scala 117:10]
  assign _GEN_3839 = 6'h3d == _T_378 ? welem[61] : _GEN_3838; // @[Execute.scala 117:10]
  assign _GEN_3840 = 6'h3e == _T_378 ? welem[62] : _GEN_3839; // @[Execute.scala 117:10]
  assign _GEN_3841 = 6'h3f == _T_378 ? welem[63] : _GEN_3840; // @[Execute.scala 117:10]
  assign _T_381 = _T_372 ? _GEN_3777 : _GEN_3841; // @[Execute.scala 117:10]
  assign _T_382 = r < 6'h23; // @[Execute.scala 117:15]
  assign _T_384 = r - 6'h23; // @[Execute.scala 117:37]
  assign _T_388 = 6'h1d + r; // @[Execute.scala 117:60]
  assign _GEN_3843 = 6'h1 == _T_384 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3844 = 6'h2 == _T_384 ? welem[2] : _GEN_3843; // @[Execute.scala 117:10]
  assign _GEN_3845 = 6'h3 == _T_384 ? welem[3] : _GEN_3844; // @[Execute.scala 117:10]
  assign _GEN_3846 = 6'h4 == _T_384 ? welem[4] : _GEN_3845; // @[Execute.scala 117:10]
  assign _GEN_3847 = 6'h5 == _T_384 ? welem[5] : _GEN_3846; // @[Execute.scala 117:10]
  assign _GEN_3848 = 6'h6 == _T_384 ? welem[6] : _GEN_3847; // @[Execute.scala 117:10]
  assign _GEN_3849 = 6'h7 == _T_384 ? welem[7] : _GEN_3848; // @[Execute.scala 117:10]
  assign _GEN_3850 = 6'h8 == _T_384 ? welem[8] : _GEN_3849; // @[Execute.scala 117:10]
  assign _GEN_3851 = 6'h9 == _T_384 ? welem[9] : _GEN_3850; // @[Execute.scala 117:10]
  assign _GEN_3852 = 6'ha == _T_384 ? welem[10] : _GEN_3851; // @[Execute.scala 117:10]
  assign _GEN_3853 = 6'hb == _T_384 ? welem[11] : _GEN_3852; // @[Execute.scala 117:10]
  assign _GEN_3854 = 6'hc == _T_384 ? welem[12] : _GEN_3853; // @[Execute.scala 117:10]
  assign _GEN_3855 = 6'hd == _T_384 ? welem[13] : _GEN_3854; // @[Execute.scala 117:10]
  assign _GEN_3856 = 6'he == _T_384 ? welem[14] : _GEN_3855; // @[Execute.scala 117:10]
  assign _GEN_3857 = 6'hf == _T_384 ? welem[15] : _GEN_3856; // @[Execute.scala 117:10]
  assign _GEN_3858 = 6'h10 == _T_384 ? welem[16] : _GEN_3857; // @[Execute.scala 117:10]
  assign _GEN_3859 = 6'h11 == _T_384 ? welem[17] : _GEN_3858; // @[Execute.scala 117:10]
  assign _GEN_3860 = 6'h12 == _T_384 ? welem[18] : _GEN_3859; // @[Execute.scala 117:10]
  assign _GEN_3861 = 6'h13 == _T_384 ? welem[19] : _GEN_3860; // @[Execute.scala 117:10]
  assign _GEN_3862 = 6'h14 == _T_384 ? welem[20] : _GEN_3861; // @[Execute.scala 117:10]
  assign _GEN_3863 = 6'h15 == _T_384 ? welem[21] : _GEN_3862; // @[Execute.scala 117:10]
  assign _GEN_3864 = 6'h16 == _T_384 ? welem[22] : _GEN_3863; // @[Execute.scala 117:10]
  assign _GEN_3865 = 6'h17 == _T_384 ? welem[23] : _GEN_3864; // @[Execute.scala 117:10]
  assign _GEN_3866 = 6'h18 == _T_384 ? welem[24] : _GEN_3865; // @[Execute.scala 117:10]
  assign _GEN_3867 = 6'h19 == _T_384 ? welem[25] : _GEN_3866; // @[Execute.scala 117:10]
  assign _GEN_3868 = 6'h1a == _T_384 ? welem[26] : _GEN_3867; // @[Execute.scala 117:10]
  assign _GEN_3869 = 6'h1b == _T_384 ? welem[27] : _GEN_3868; // @[Execute.scala 117:10]
  assign _GEN_3870 = 6'h1c == _T_384 ? welem[28] : _GEN_3869; // @[Execute.scala 117:10]
  assign _GEN_3871 = 6'h1d == _T_384 ? welem[29] : _GEN_3870; // @[Execute.scala 117:10]
  assign _GEN_3872 = 6'h1e == _T_384 ? welem[30] : _GEN_3871; // @[Execute.scala 117:10]
  assign _GEN_3873 = 6'h1f == _T_384 ? welem[31] : _GEN_3872; // @[Execute.scala 117:10]
  assign _GEN_3874 = 6'h20 == _T_384 ? welem[32] : _GEN_3873; // @[Execute.scala 117:10]
  assign _GEN_3875 = 6'h21 == _T_384 ? welem[33] : _GEN_3874; // @[Execute.scala 117:10]
  assign _GEN_3876 = 6'h22 == _T_384 ? welem[34] : _GEN_3875; // @[Execute.scala 117:10]
  assign _GEN_3877 = 6'h23 == _T_384 ? welem[35] : _GEN_3876; // @[Execute.scala 117:10]
  assign _GEN_3878 = 6'h24 == _T_384 ? welem[36] : _GEN_3877; // @[Execute.scala 117:10]
  assign _GEN_3879 = 6'h25 == _T_384 ? welem[37] : _GEN_3878; // @[Execute.scala 117:10]
  assign _GEN_3880 = 6'h26 == _T_384 ? welem[38] : _GEN_3879; // @[Execute.scala 117:10]
  assign _GEN_3881 = 6'h27 == _T_384 ? welem[39] : _GEN_3880; // @[Execute.scala 117:10]
  assign _GEN_3882 = 6'h28 == _T_384 ? welem[40] : _GEN_3881; // @[Execute.scala 117:10]
  assign _GEN_3883 = 6'h29 == _T_384 ? welem[41] : _GEN_3882; // @[Execute.scala 117:10]
  assign _GEN_3884 = 6'h2a == _T_384 ? welem[42] : _GEN_3883; // @[Execute.scala 117:10]
  assign _GEN_3885 = 6'h2b == _T_384 ? welem[43] : _GEN_3884; // @[Execute.scala 117:10]
  assign _GEN_3886 = 6'h2c == _T_384 ? welem[44] : _GEN_3885; // @[Execute.scala 117:10]
  assign _GEN_3887 = 6'h2d == _T_384 ? welem[45] : _GEN_3886; // @[Execute.scala 117:10]
  assign _GEN_3888 = 6'h2e == _T_384 ? welem[46] : _GEN_3887; // @[Execute.scala 117:10]
  assign _GEN_3889 = 6'h2f == _T_384 ? welem[47] : _GEN_3888; // @[Execute.scala 117:10]
  assign _GEN_3890 = 6'h30 == _T_384 ? welem[48] : _GEN_3889; // @[Execute.scala 117:10]
  assign _GEN_3891 = 6'h31 == _T_384 ? welem[49] : _GEN_3890; // @[Execute.scala 117:10]
  assign _GEN_3892 = 6'h32 == _T_384 ? welem[50] : _GEN_3891; // @[Execute.scala 117:10]
  assign _GEN_3893 = 6'h33 == _T_384 ? welem[51] : _GEN_3892; // @[Execute.scala 117:10]
  assign _GEN_3894 = 6'h34 == _T_384 ? welem[52] : _GEN_3893; // @[Execute.scala 117:10]
  assign _GEN_3895 = 6'h35 == _T_384 ? welem[53] : _GEN_3894; // @[Execute.scala 117:10]
  assign _GEN_3896 = 6'h36 == _T_384 ? welem[54] : _GEN_3895; // @[Execute.scala 117:10]
  assign _GEN_3897 = 6'h37 == _T_384 ? welem[55] : _GEN_3896; // @[Execute.scala 117:10]
  assign _GEN_3898 = 6'h38 == _T_384 ? welem[56] : _GEN_3897; // @[Execute.scala 117:10]
  assign _GEN_3899 = 6'h39 == _T_384 ? welem[57] : _GEN_3898; // @[Execute.scala 117:10]
  assign _GEN_3900 = 6'h3a == _T_384 ? welem[58] : _GEN_3899; // @[Execute.scala 117:10]
  assign _GEN_3901 = 6'h3b == _T_384 ? welem[59] : _GEN_3900; // @[Execute.scala 117:10]
  assign _GEN_3902 = 6'h3c == _T_384 ? welem[60] : _GEN_3901; // @[Execute.scala 117:10]
  assign _GEN_3903 = 6'h3d == _T_384 ? welem[61] : _GEN_3902; // @[Execute.scala 117:10]
  assign _GEN_3904 = 6'h3e == _T_384 ? welem[62] : _GEN_3903; // @[Execute.scala 117:10]
  assign _GEN_3905 = 6'h3f == _T_384 ? welem[63] : _GEN_3904; // @[Execute.scala 117:10]
  assign _GEN_3907 = 6'h1 == _T_388 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3908 = 6'h2 == _T_388 ? welem[2] : _GEN_3907; // @[Execute.scala 117:10]
  assign _GEN_3909 = 6'h3 == _T_388 ? welem[3] : _GEN_3908; // @[Execute.scala 117:10]
  assign _GEN_3910 = 6'h4 == _T_388 ? welem[4] : _GEN_3909; // @[Execute.scala 117:10]
  assign _GEN_3911 = 6'h5 == _T_388 ? welem[5] : _GEN_3910; // @[Execute.scala 117:10]
  assign _GEN_3912 = 6'h6 == _T_388 ? welem[6] : _GEN_3911; // @[Execute.scala 117:10]
  assign _GEN_3913 = 6'h7 == _T_388 ? welem[7] : _GEN_3912; // @[Execute.scala 117:10]
  assign _GEN_3914 = 6'h8 == _T_388 ? welem[8] : _GEN_3913; // @[Execute.scala 117:10]
  assign _GEN_3915 = 6'h9 == _T_388 ? welem[9] : _GEN_3914; // @[Execute.scala 117:10]
  assign _GEN_3916 = 6'ha == _T_388 ? welem[10] : _GEN_3915; // @[Execute.scala 117:10]
  assign _GEN_3917 = 6'hb == _T_388 ? welem[11] : _GEN_3916; // @[Execute.scala 117:10]
  assign _GEN_3918 = 6'hc == _T_388 ? welem[12] : _GEN_3917; // @[Execute.scala 117:10]
  assign _GEN_3919 = 6'hd == _T_388 ? welem[13] : _GEN_3918; // @[Execute.scala 117:10]
  assign _GEN_3920 = 6'he == _T_388 ? welem[14] : _GEN_3919; // @[Execute.scala 117:10]
  assign _GEN_3921 = 6'hf == _T_388 ? welem[15] : _GEN_3920; // @[Execute.scala 117:10]
  assign _GEN_3922 = 6'h10 == _T_388 ? welem[16] : _GEN_3921; // @[Execute.scala 117:10]
  assign _GEN_3923 = 6'h11 == _T_388 ? welem[17] : _GEN_3922; // @[Execute.scala 117:10]
  assign _GEN_3924 = 6'h12 == _T_388 ? welem[18] : _GEN_3923; // @[Execute.scala 117:10]
  assign _GEN_3925 = 6'h13 == _T_388 ? welem[19] : _GEN_3924; // @[Execute.scala 117:10]
  assign _GEN_3926 = 6'h14 == _T_388 ? welem[20] : _GEN_3925; // @[Execute.scala 117:10]
  assign _GEN_3927 = 6'h15 == _T_388 ? welem[21] : _GEN_3926; // @[Execute.scala 117:10]
  assign _GEN_3928 = 6'h16 == _T_388 ? welem[22] : _GEN_3927; // @[Execute.scala 117:10]
  assign _GEN_3929 = 6'h17 == _T_388 ? welem[23] : _GEN_3928; // @[Execute.scala 117:10]
  assign _GEN_3930 = 6'h18 == _T_388 ? welem[24] : _GEN_3929; // @[Execute.scala 117:10]
  assign _GEN_3931 = 6'h19 == _T_388 ? welem[25] : _GEN_3930; // @[Execute.scala 117:10]
  assign _GEN_3932 = 6'h1a == _T_388 ? welem[26] : _GEN_3931; // @[Execute.scala 117:10]
  assign _GEN_3933 = 6'h1b == _T_388 ? welem[27] : _GEN_3932; // @[Execute.scala 117:10]
  assign _GEN_3934 = 6'h1c == _T_388 ? welem[28] : _GEN_3933; // @[Execute.scala 117:10]
  assign _GEN_3935 = 6'h1d == _T_388 ? welem[29] : _GEN_3934; // @[Execute.scala 117:10]
  assign _GEN_3936 = 6'h1e == _T_388 ? welem[30] : _GEN_3935; // @[Execute.scala 117:10]
  assign _GEN_3937 = 6'h1f == _T_388 ? welem[31] : _GEN_3936; // @[Execute.scala 117:10]
  assign _GEN_3938 = 6'h20 == _T_388 ? welem[32] : _GEN_3937; // @[Execute.scala 117:10]
  assign _GEN_3939 = 6'h21 == _T_388 ? welem[33] : _GEN_3938; // @[Execute.scala 117:10]
  assign _GEN_3940 = 6'h22 == _T_388 ? welem[34] : _GEN_3939; // @[Execute.scala 117:10]
  assign _GEN_3941 = 6'h23 == _T_388 ? welem[35] : _GEN_3940; // @[Execute.scala 117:10]
  assign _GEN_3942 = 6'h24 == _T_388 ? welem[36] : _GEN_3941; // @[Execute.scala 117:10]
  assign _GEN_3943 = 6'h25 == _T_388 ? welem[37] : _GEN_3942; // @[Execute.scala 117:10]
  assign _GEN_3944 = 6'h26 == _T_388 ? welem[38] : _GEN_3943; // @[Execute.scala 117:10]
  assign _GEN_3945 = 6'h27 == _T_388 ? welem[39] : _GEN_3944; // @[Execute.scala 117:10]
  assign _GEN_3946 = 6'h28 == _T_388 ? welem[40] : _GEN_3945; // @[Execute.scala 117:10]
  assign _GEN_3947 = 6'h29 == _T_388 ? welem[41] : _GEN_3946; // @[Execute.scala 117:10]
  assign _GEN_3948 = 6'h2a == _T_388 ? welem[42] : _GEN_3947; // @[Execute.scala 117:10]
  assign _GEN_3949 = 6'h2b == _T_388 ? welem[43] : _GEN_3948; // @[Execute.scala 117:10]
  assign _GEN_3950 = 6'h2c == _T_388 ? welem[44] : _GEN_3949; // @[Execute.scala 117:10]
  assign _GEN_3951 = 6'h2d == _T_388 ? welem[45] : _GEN_3950; // @[Execute.scala 117:10]
  assign _GEN_3952 = 6'h2e == _T_388 ? welem[46] : _GEN_3951; // @[Execute.scala 117:10]
  assign _GEN_3953 = 6'h2f == _T_388 ? welem[47] : _GEN_3952; // @[Execute.scala 117:10]
  assign _GEN_3954 = 6'h30 == _T_388 ? welem[48] : _GEN_3953; // @[Execute.scala 117:10]
  assign _GEN_3955 = 6'h31 == _T_388 ? welem[49] : _GEN_3954; // @[Execute.scala 117:10]
  assign _GEN_3956 = 6'h32 == _T_388 ? welem[50] : _GEN_3955; // @[Execute.scala 117:10]
  assign _GEN_3957 = 6'h33 == _T_388 ? welem[51] : _GEN_3956; // @[Execute.scala 117:10]
  assign _GEN_3958 = 6'h34 == _T_388 ? welem[52] : _GEN_3957; // @[Execute.scala 117:10]
  assign _GEN_3959 = 6'h35 == _T_388 ? welem[53] : _GEN_3958; // @[Execute.scala 117:10]
  assign _GEN_3960 = 6'h36 == _T_388 ? welem[54] : _GEN_3959; // @[Execute.scala 117:10]
  assign _GEN_3961 = 6'h37 == _T_388 ? welem[55] : _GEN_3960; // @[Execute.scala 117:10]
  assign _GEN_3962 = 6'h38 == _T_388 ? welem[56] : _GEN_3961; // @[Execute.scala 117:10]
  assign _GEN_3963 = 6'h39 == _T_388 ? welem[57] : _GEN_3962; // @[Execute.scala 117:10]
  assign _GEN_3964 = 6'h3a == _T_388 ? welem[58] : _GEN_3963; // @[Execute.scala 117:10]
  assign _GEN_3965 = 6'h3b == _T_388 ? welem[59] : _GEN_3964; // @[Execute.scala 117:10]
  assign _GEN_3966 = 6'h3c == _T_388 ? welem[60] : _GEN_3965; // @[Execute.scala 117:10]
  assign _GEN_3967 = 6'h3d == _T_388 ? welem[61] : _GEN_3966; // @[Execute.scala 117:10]
  assign _GEN_3968 = 6'h3e == _T_388 ? welem[62] : _GEN_3967; // @[Execute.scala 117:10]
  assign _GEN_3969 = 6'h3f == _T_388 ? welem[63] : _GEN_3968; // @[Execute.scala 117:10]
  assign _T_391 = _T_382 ? _GEN_3905 : _GEN_3969; // @[Execute.scala 117:10]
  assign _T_392 = r < 6'h22; // @[Execute.scala 117:15]
  assign _T_394 = r - 6'h22; // @[Execute.scala 117:37]
  assign _T_398 = 6'h1e + r; // @[Execute.scala 117:60]
  assign _GEN_3971 = 6'h1 == _T_394 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_3972 = 6'h2 == _T_394 ? welem[2] : _GEN_3971; // @[Execute.scala 117:10]
  assign _GEN_3973 = 6'h3 == _T_394 ? welem[3] : _GEN_3972; // @[Execute.scala 117:10]
  assign _GEN_3974 = 6'h4 == _T_394 ? welem[4] : _GEN_3973; // @[Execute.scala 117:10]
  assign _GEN_3975 = 6'h5 == _T_394 ? welem[5] : _GEN_3974; // @[Execute.scala 117:10]
  assign _GEN_3976 = 6'h6 == _T_394 ? welem[6] : _GEN_3975; // @[Execute.scala 117:10]
  assign _GEN_3977 = 6'h7 == _T_394 ? welem[7] : _GEN_3976; // @[Execute.scala 117:10]
  assign _GEN_3978 = 6'h8 == _T_394 ? welem[8] : _GEN_3977; // @[Execute.scala 117:10]
  assign _GEN_3979 = 6'h9 == _T_394 ? welem[9] : _GEN_3978; // @[Execute.scala 117:10]
  assign _GEN_3980 = 6'ha == _T_394 ? welem[10] : _GEN_3979; // @[Execute.scala 117:10]
  assign _GEN_3981 = 6'hb == _T_394 ? welem[11] : _GEN_3980; // @[Execute.scala 117:10]
  assign _GEN_3982 = 6'hc == _T_394 ? welem[12] : _GEN_3981; // @[Execute.scala 117:10]
  assign _GEN_3983 = 6'hd == _T_394 ? welem[13] : _GEN_3982; // @[Execute.scala 117:10]
  assign _GEN_3984 = 6'he == _T_394 ? welem[14] : _GEN_3983; // @[Execute.scala 117:10]
  assign _GEN_3985 = 6'hf == _T_394 ? welem[15] : _GEN_3984; // @[Execute.scala 117:10]
  assign _GEN_3986 = 6'h10 == _T_394 ? welem[16] : _GEN_3985; // @[Execute.scala 117:10]
  assign _GEN_3987 = 6'h11 == _T_394 ? welem[17] : _GEN_3986; // @[Execute.scala 117:10]
  assign _GEN_3988 = 6'h12 == _T_394 ? welem[18] : _GEN_3987; // @[Execute.scala 117:10]
  assign _GEN_3989 = 6'h13 == _T_394 ? welem[19] : _GEN_3988; // @[Execute.scala 117:10]
  assign _GEN_3990 = 6'h14 == _T_394 ? welem[20] : _GEN_3989; // @[Execute.scala 117:10]
  assign _GEN_3991 = 6'h15 == _T_394 ? welem[21] : _GEN_3990; // @[Execute.scala 117:10]
  assign _GEN_3992 = 6'h16 == _T_394 ? welem[22] : _GEN_3991; // @[Execute.scala 117:10]
  assign _GEN_3993 = 6'h17 == _T_394 ? welem[23] : _GEN_3992; // @[Execute.scala 117:10]
  assign _GEN_3994 = 6'h18 == _T_394 ? welem[24] : _GEN_3993; // @[Execute.scala 117:10]
  assign _GEN_3995 = 6'h19 == _T_394 ? welem[25] : _GEN_3994; // @[Execute.scala 117:10]
  assign _GEN_3996 = 6'h1a == _T_394 ? welem[26] : _GEN_3995; // @[Execute.scala 117:10]
  assign _GEN_3997 = 6'h1b == _T_394 ? welem[27] : _GEN_3996; // @[Execute.scala 117:10]
  assign _GEN_3998 = 6'h1c == _T_394 ? welem[28] : _GEN_3997; // @[Execute.scala 117:10]
  assign _GEN_3999 = 6'h1d == _T_394 ? welem[29] : _GEN_3998; // @[Execute.scala 117:10]
  assign _GEN_4000 = 6'h1e == _T_394 ? welem[30] : _GEN_3999; // @[Execute.scala 117:10]
  assign _GEN_4001 = 6'h1f == _T_394 ? welem[31] : _GEN_4000; // @[Execute.scala 117:10]
  assign _GEN_4002 = 6'h20 == _T_394 ? welem[32] : _GEN_4001; // @[Execute.scala 117:10]
  assign _GEN_4003 = 6'h21 == _T_394 ? welem[33] : _GEN_4002; // @[Execute.scala 117:10]
  assign _GEN_4004 = 6'h22 == _T_394 ? welem[34] : _GEN_4003; // @[Execute.scala 117:10]
  assign _GEN_4005 = 6'h23 == _T_394 ? welem[35] : _GEN_4004; // @[Execute.scala 117:10]
  assign _GEN_4006 = 6'h24 == _T_394 ? welem[36] : _GEN_4005; // @[Execute.scala 117:10]
  assign _GEN_4007 = 6'h25 == _T_394 ? welem[37] : _GEN_4006; // @[Execute.scala 117:10]
  assign _GEN_4008 = 6'h26 == _T_394 ? welem[38] : _GEN_4007; // @[Execute.scala 117:10]
  assign _GEN_4009 = 6'h27 == _T_394 ? welem[39] : _GEN_4008; // @[Execute.scala 117:10]
  assign _GEN_4010 = 6'h28 == _T_394 ? welem[40] : _GEN_4009; // @[Execute.scala 117:10]
  assign _GEN_4011 = 6'h29 == _T_394 ? welem[41] : _GEN_4010; // @[Execute.scala 117:10]
  assign _GEN_4012 = 6'h2a == _T_394 ? welem[42] : _GEN_4011; // @[Execute.scala 117:10]
  assign _GEN_4013 = 6'h2b == _T_394 ? welem[43] : _GEN_4012; // @[Execute.scala 117:10]
  assign _GEN_4014 = 6'h2c == _T_394 ? welem[44] : _GEN_4013; // @[Execute.scala 117:10]
  assign _GEN_4015 = 6'h2d == _T_394 ? welem[45] : _GEN_4014; // @[Execute.scala 117:10]
  assign _GEN_4016 = 6'h2e == _T_394 ? welem[46] : _GEN_4015; // @[Execute.scala 117:10]
  assign _GEN_4017 = 6'h2f == _T_394 ? welem[47] : _GEN_4016; // @[Execute.scala 117:10]
  assign _GEN_4018 = 6'h30 == _T_394 ? welem[48] : _GEN_4017; // @[Execute.scala 117:10]
  assign _GEN_4019 = 6'h31 == _T_394 ? welem[49] : _GEN_4018; // @[Execute.scala 117:10]
  assign _GEN_4020 = 6'h32 == _T_394 ? welem[50] : _GEN_4019; // @[Execute.scala 117:10]
  assign _GEN_4021 = 6'h33 == _T_394 ? welem[51] : _GEN_4020; // @[Execute.scala 117:10]
  assign _GEN_4022 = 6'h34 == _T_394 ? welem[52] : _GEN_4021; // @[Execute.scala 117:10]
  assign _GEN_4023 = 6'h35 == _T_394 ? welem[53] : _GEN_4022; // @[Execute.scala 117:10]
  assign _GEN_4024 = 6'h36 == _T_394 ? welem[54] : _GEN_4023; // @[Execute.scala 117:10]
  assign _GEN_4025 = 6'h37 == _T_394 ? welem[55] : _GEN_4024; // @[Execute.scala 117:10]
  assign _GEN_4026 = 6'h38 == _T_394 ? welem[56] : _GEN_4025; // @[Execute.scala 117:10]
  assign _GEN_4027 = 6'h39 == _T_394 ? welem[57] : _GEN_4026; // @[Execute.scala 117:10]
  assign _GEN_4028 = 6'h3a == _T_394 ? welem[58] : _GEN_4027; // @[Execute.scala 117:10]
  assign _GEN_4029 = 6'h3b == _T_394 ? welem[59] : _GEN_4028; // @[Execute.scala 117:10]
  assign _GEN_4030 = 6'h3c == _T_394 ? welem[60] : _GEN_4029; // @[Execute.scala 117:10]
  assign _GEN_4031 = 6'h3d == _T_394 ? welem[61] : _GEN_4030; // @[Execute.scala 117:10]
  assign _GEN_4032 = 6'h3e == _T_394 ? welem[62] : _GEN_4031; // @[Execute.scala 117:10]
  assign _GEN_4033 = 6'h3f == _T_394 ? welem[63] : _GEN_4032; // @[Execute.scala 117:10]
  assign _GEN_4035 = 6'h1 == _T_398 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4036 = 6'h2 == _T_398 ? welem[2] : _GEN_4035; // @[Execute.scala 117:10]
  assign _GEN_4037 = 6'h3 == _T_398 ? welem[3] : _GEN_4036; // @[Execute.scala 117:10]
  assign _GEN_4038 = 6'h4 == _T_398 ? welem[4] : _GEN_4037; // @[Execute.scala 117:10]
  assign _GEN_4039 = 6'h5 == _T_398 ? welem[5] : _GEN_4038; // @[Execute.scala 117:10]
  assign _GEN_4040 = 6'h6 == _T_398 ? welem[6] : _GEN_4039; // @[Execute.scala 117:10]
  assign _GEN_4041 = 6'h7 == _T_398 ? welem[7] : _GEN_4040; // @[Execute.scala 117:10]
  assign _GEN_4042 = 6'h8 == _T_398 ? welem[8] : _GEN_4041; // @[Execute.scala 117:10]
  assign _GEN_4043 = 6'h9 == _T_398 ? welem[9] : _GEN_4042; // @[Execute.scala 117:10]
  assign _GEN_4044 = 6'ha == _T_398 ? welem[10] : _GEN_4043; // @[Execute.scala 117:10]
  assign _GEN_4045 = 6'hb == _T_398 ? welem[11] : _GEN_4044; // @[Execute.scala 117:10]
  assign _GEN_4046 = 6'hc == _T_398 ? welem[12] : _GEN_4045; // @[Execute.scala 117:10]
  assign _GEN_4047 = 6'hd == _T_398 ? welem[13] : _GEN_4046; // @[Execute.scala 117:10]
  assign _GEN_4048 = 6'he == _T_398 ? welem[14] : _GEN_4047; // @[Execute.scala 117:10]
  assign _GEN_4049 = 6'hf == _T_398 ? welem[15] : _GEN_4048; // @[Execute.scala 117:10]
  assign _GEN_4050 = 6'h10 == _T_398 ? welem[16] : _GEN_4049; // @[Execute.scala 117:10]
  assign _GEN_4051 = 6'h11 == _T_398 ? welem[17] : _GEN_4050; // @[Execute.scala 117:10]
  assign _GEN_4052 = 6'h12 == _T_398 ? welem[18] : _GEN_4051; // @[Execute.scala 117:10]
  assign _GEN_4053 = 6'h13 == _T_398 ? welem[19] : _GEN_4052; // @[Execute.scala 117:10]
  assign _GEN_4054 = 6'h14 == _T_398 ? welem[20] : _GEN_4053; // @[Execute.scala 117:10]
  assign _GEN_4055 = 6'h15 == _T_398 ? welem[21] : _GEN_4054; // @[Execute.scala 117:10]
  assign _GEN_4056 = 6'h16 == _T_398 ? welem[22] : _GEN_4055; // @[Execute.scala 117:10]
  assign _GEN_4057 = 6'h17 == _T_398 ? welem[23] : _GEN_4056; // @[Execute.scala 117:10]
  assign _GEN_4058 = 6'h18 == _T_398 ? welem[24] : _GEN_4057; // @[Execute.scala 117:10]
  assign _GEN_4059 = 6'h19 == _T_398 ? welem[25] : _GEN_4058; // @[Execute.scala 117:10]
  assign _GEN_4060 = 6'h1a == _T_398 ? welem[26] : _GEN_4059; // @[Execute.scala 117:10]
  assign _GEN_4061 = 6'h1b == _T_398 ? welem[27] : _GEN_4060; // @[Execute.scala 117:10]
  assign _GEN_4062 = 6'h1c == _T_398 ? welem[28] : _GEN_4061; // @[Execute.scala 117:10]
  assign _GEN_4063 = 6'h1d == _T_398 ? welem[29] : _GEN_4062; // @[Execute.scala 117:10]
  assign _GEN_4064 = 6'h1e == _T_398 ? welem[30] : _GEN_4063; // @[Execute.scala 117:10]
  assign _GEN_4065 = 6'h1f == _T_398 ? welem[31] : _GEN_4064; // @[Execute.scala 117:10]
  assign _GEN_4066 = 6'h20 == _T_398 ? welem[32] : _GEN_4065; // @[Execute.scala 117:10]
  assign _GEN_4067 = 6'h21 == _T_398 ? welem[33] : _GEN_4066; // @[Execute.scala 117:10]
  assign _GEN_4068 = 6'h22 == _T_398 ? welem[34] : _GEN_4067; // @[Execute.scala 117:10]
  assign _GEN_4069 = 6'h23 == _T_398 ? welem[35] : _GEN_4068; // @[Execute.scala 117:10]
  assign _GEN_4070 = 6'h24 == _T_398 ? welem[36] : _GEN_4069; // @[Execute.scala 117:10]
  assign _GEN_4071 = 6'h25 == _T_398 ? welem[37] : _GEN_4070; // @[Execute.scala 117:10]
  assign _GEN_4072 = 6'h26 == _T_398 ? welem[38] : _GEN_4071; // @[Execute.scala 117:10]
  assign _GEN_4073 = 6'h27 == _T_398 ? welem[39] : _GEN_4072; // @[Execute.scala 117:10]
  assign _GEN_4074 = 6'h28 == _T_398 ? welem[40] : _GEN_4073; // @[Execute.scala 117:10]
  assign _GEN_4075 = 6'h29 == _T_398 ? welem[41] : _GEN_4074; // @[Execute.scala 117:10]
  assign _GEN_4076 = 6'h2a == _T_398 ? welem[42] : _GEN_4075; // @[Execute.scala 117:10]
  assign _GEN_4077 = 6'h2b == _T_398 ? welem[43] : _GEN_4076; // @[Execute.scala 117:10]
  assign _GEN_4078 = 6'h2c == _T_398 ? welem[44] : _GEN_4077; // @[Execute.scala 117:10]
  assign _GEN_4079 = 6'h2d == _T_398 ? welem[45] : _GEN_4078; // @[Execute.scala 117:10]
  assign _GEN_4080 = 6'h2e == _T_398 ? welem[46] : _GEN_4079; // @[Execute.scala 117:10]
  assign _GEN_4081 = 6'h2f == _T_398 ? welem[47] : _GEN_4080; // @[Execute.scala 117:10]
  assign _GEN_4082 = 6'h30 == _T_398 ? welem[48] : _GEN_4081; // @[Execute.scala 117:10]
  assign _GEN_4083 = 6'h31 == _T_398 ? welem[49] : _GEN_4082; // @[Execute.scala 117:10]
  assign _GEN_4084 = 6'h32 == _T_398 ? welem[50] : _GEN_4083; // @[Execute.scala 117:10]
  assign _GEN_4085 = 6'h33 == _T_398 ? welem[51] : _GEN_4084; // @[Execute.scala 117:10]
  assign _GEN_4086 = 6'h34 == _T_398 ? welem[52] : _GEN_4085; // @[Execute.scala 117:10]
  assign _GEN_4087 = 6'h35 == _T_398 ? welem[53] : _GEN_4086; // @[Execute.scala 117:10]
  assign _GEN_4088 = 6'h36 == _T_398 ? welem[54] : _GEN_4087; // @[Execute.scala 117:10]
  assign _GEN_4089 = 6'h37 == _T_398 ? welem[55] : _GEN_4088; // @[Execute.scala 117:10]
  assign _GEN_4090 = 6'h38 == _T_398 ? welem[56] : _GEN_4089; // @[Execute.scala 117:10]
  assign _GEN_4091 = 6'h39 == _T_398 ? welem[57] : _GEN_4090; // @[Execute.scala 117:10]
  assign _GEN_4092 = 6'h3a == _T_398 ? welem[58] : _GEN_4091; // @[Execute.scala 117:10]
  assign _GEN_4093 = 6'h3b == _T_398 ? welem[59] : _GEN_4092; // @[Execute.scala 117:10]
  assign _GEN_4094 = 6'h3c == _T_398 ? welem[60] : _GEN_4093; // @[Execute.scala 117:10]
  assign _GEN_4095 = 6'h3d == _T_398 ? welem[61] : _GEN_4094; // @[Execute.scala 117:10]
  assign _GEN_4096 = 6'h3e == _T_398 ? welem[62] : _GEN_4095; // @[Execute.scala 117:10]
  assign _GEN_4097 = 6'h3f == _T_398 ? welem[63] : _GEN_4096; // @[Execute.scala 117:10]
  assign _T_401 = _T_392 ? _GEN_4033 : _GEN_4097; // @[Execute.scala 117:10]
  assign _T_402 = r < 6'h21; // @[Execute.scala 117:15]
  assign _T_404 = r - 6'h21; // @[Execute.scala 117:37]
  assign _T_408 = 6'h1f + r; // @[Execute.scala 117:60]
  assign _GEN_4099 = 6'h1 == _T_404 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4100 = 6'h2 == _T_404 ? welem[2] : _GEN_4099; // @[Execute.scala 117:10]
  assign _GEN_4101 = 6'h3 == _T_404 ? welem[3] : _GEN_4100; // @[Execute.scala 117:10]
  assign _GEN_4102 = 6'h4 == _T_404 ? welem[4] : _GEN_4101; // @[Execute.scala 117:10]
  assign _GEN_4103 = 6'h5 == _T_404 ? welem[5] : _GEN_4102; // @[Execute.scala 117:10]
  assign _GEN_4104 = 6'h6 == _T_404 ? welem[6] : _GEN_4103; // @[Execute.scala 117:10]
  assign _GEN_4105 = 6'h7 == _T_404 ? welem[7] : _GEN_4104; // @[Execute.scala 117:10]
  assign _GEN_4106 = 6'h8 == _T_404 ? welem[8] : _GEN_4105; // @[Execute.scala 117:10]
  assign _GEN_4107 = 6'h9 == _T_404 ? welem[9] : _GEN_4106; // @[Execute.scala 117:10]
  assign _GEN_4108 = 6'ha == _T_404 ? welem[10] : _GEN_4107; // @[Execute.scala 117:10]
  assign _GEN_4109 = 6'hb == _T_404 ? welem[11] : _GEN_4108; // @[Execute.scala 117:10]
  assign _GEN_4110 = 6'hc == _T_404 ? welem[12] : _GEN_4109; // @[Execute.scala 117:10]
  assign _GEN_4111 = 6'hd == _T_404 ? welem[13] : _GEN_4110; // @[Execute.scala 117:10]
  assign _GEN_4112 = 6'he == _T_404 ? welem[14] : _GEN_4111; // @[Execute.scala 117:10]
  assign _GEN_4113 = 6'hf == _T_404 ? welem[15] : _GEN_4112; // @[Execute.scala 117:10]
  assign _GEN_4114 = 6'h10 == _T_404 ? welem[16] : _GEN_4113; // @[Execute.scala 117:10]
  assign _GEN_4115 = 6'h11 == _T_404 ? welem[17] : _GEN_4114; // @[Execute.scala 117:10]
  assign _GEN_4116 = 6'h12 == _T_404 ? welem[18] : _GEN_4115; // @[Execute.scala 117:10]
  assign _GEN_4117 = 6'h13 == _T_404 ? welem[19] : _GEN_4116; // @[Execute.scala 117:10]
  assign _GEN_4118 = 6'h14 == _T_404 ? welem[20] : _GEN_4117; // @[Execute.scala 117:10]
  assign _GEN_4119 = 6'h15 == _T_404 ? welem[21] : _GEN_4118; // @[Execute.scala 117:10]
  assign _GEN_4120 = 6'h16 == _T_404 ? welem[22] : _GEN_4119; // @[Execute.scala 117:10]
  assign _GEN_4121 = 6'h17 == _T_404 ? welem[23] : _GEN_4120; // @[Execute.scala 117:10]
  assign _GEN_4122 = 6'h18 == _T_404 ? welem[24] : _GEN_4121; // @[Execute.scala 117:10]
  assign _GEN_4123 = 6'h19 == _T_404 ? welem[25] : _GEN_4122; // @[Execute.scala 117:10]
  assign _GEN_4124 = 6'h1a == _T_404 ? welem[26] : _GEN_4123; // @[Execute.scala 117:10]
  assign _GEN_4125 = 6'h1b == _T_404 ? welem[27] : _GEN_4124; // @[Execute.scala 117:10]
  assign _GEN_4126 = 6'h1c == _T_404 ? welem[28] : _GEN_4125; // @[Execute.scala 117:10]
  assign _GEN_4127 = 6'h1d == _T_404 ? welem[29] : _GEN_4126; // @[Execute.scala 117:10]
  assign _GEN_4128 = 6'h1e == _T_404 ? welem[30] : _GEN_4127; // @[Execute.scala 117:10]
  assign _GEN_4129 = 6'h1f == _T_404 ? welem[31] : _GEN_4128; // @[Execute.scala 117:10]
  assign _GEN_4130 = 6'h20 == _T_404 ? welem[32] : _GEN_4129; // @[Execute.scala 117:10]
  assign _GEN_4131 = 6'h21 == _T_404 ? welem[33] : _GEN_4130; // @[Execute.scala 117:10]
  assign _GEN_4132 = 6'h22 == _T_404 ? welem[34] : _GEN_4131; // @[Execute.scala 117:10]
  assign _GEN_4133 = 6'h23 == _T_404 ? welem[35] : _GEN_4132; // @[Execute.scala 117:10]
  assign _GEN_4134 = 6'h24 == _T_404 ? welem[36] : _GEN_4133; // @[Execute.scala 117:10]
  assign _GEN_4135 = 6'h25 == _T_404 ? welem[37] : _GEN_4134; // @[Execute.scala 117:10]
  assign _GEN_4136 = 6'h26 == _T_404 ? welem[38] : _GEN_4135; // @[Execute.scala 117:10]
  assign _GEN_4137 = 6'h27 == _T_404 ? welem[39] : _GEN_4136; // @[Execute.scala 117:10]
  assign _GEN_4138 = 6'h28 == _T_404 ? welem[40] : _GEN_4137; // @[Execute.scala 117:10]
  assign _GEN_4139 = 6'h29 == _T_404 ? welem[41] : _GEN_4138; // @[Execute.scala 117:10]
  assign _GEN_4140 = 6'h2a == _T_404 ? welem[42] : _GEN_4139; // @[Execute.scala 117:10]
  assign _GEN_4141 = 6'h2b == _T_404 ? welem[43] : _GEN_4140; // @[Execute.scala 117:10]
  assign _GEN_4142 = 6'h2c == _T_404 ? welem[44] : _GEN_4141; // @[Execute.scala 117:10]
  assign _GEN_4143 = 6'h2d == _T_404 ? welem[45] : _GEN_4142; // @[Execute.scala 117:10]
  assign _GEN_4144 = 6'h2e == _T_404 ? welem[46] : _GEN_4143; // @[Execute.scala 117:10]
  assign _GEN_4145 = 6'h2f == _T_404 ? welem[47] : _GEN_4144; // @[Execute.scala 117:10]
  assign _GEN_4146 = 6'h30 == _T_404 ? welem[48] : _GEN_4145; // @[Execute.scala 117:10]
  assign _GEN_4147 = 6'h31 == _T_404 ? welem[49] : _GEN_4146; // @[Execute.scala 117:10]
  assign _GEN_4148 = 6'h32 == _T_404 ? welem[50] : _GEN_4147; // @[Execute.scala 117:10]
  assign _GEN_4149 = 6'h33 == _T_404 ? welem[51] : _GEN_4148; // @[Execute.scala 117:10]
  assign _GEN_4150 = 6'h34 == _T_404 ? welem[52] : _GEN_4149; // @[Execute.scala 117:10]
  assign _GEN_4151 = 6'h35 == _T_404 ? welem[53] : _GEN_4150; // @[Execute.scala 117:10]
  assign _GEN_4152 = 6'h36 == _T_404 ? welem[54] : _GEN_4151; // @[Execute.scala 117:10]
  assign _GEN_4153 = 6'h37 == _T_404 ? welem[55] : _GEN_4152; // @[Execute.scala 117:10]
  assign _GEN_4154 = 6'h38 == _T_404 ? welem[56] : _GEN_4153; // @[Execute.scala 117:10]
  assign _GEN_4155 = 6'h39 == _T_404 ? welem[57] : _GEN_4154; // @[Execute.scala 117:10]
  assign _GEN_4156 = 6'h3a == _T_404 ? welem[58] : _GEN_4155; // @[Execute.scala 117:10]
  assign _GEN_4157 = 6'h3b == _T_404 ? welem[59] : _GEN_4156; // @[Execute.scala 117:10]
  assign _GEN_4158 = 6'h3c == _T_404 ? welem[60] : _GEN_4157; // @[Execute.scala 117:10]
  assign _GEN_4159 = 6'h3d == _T_404 ? welem[61] : _GEN_4158; // @[Execute.scala 117:10]
  assign _GEN_4160 = 6'h3e == _T_404 ? welem[62] : _GEN_4159; // @[Execute.scala 117:10]
  assign _GEN_4161 = 6'h3f == _T_404 ? welem[63] : _GEN_4160; // @[Execute.scala 117:10]
  assign _GEN_4163 = 6'h1 == _T_408 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4164 = 6'h2 == _T_408 ? welem[2] : _GEN_4163; // @[Execute.scala 117:10]
  assign _GEN_4165 = 6'h3 == _T_408 ? welem[3] : _GEN_4164; // @[Execute.scala 117:10]
  assign _GEN_4166 = 6'h4 == _T_408 ? welem[4] : _GEN_4165; // @[Execute.scala 117:10]
  assign _GEN_4167 = 6'h5 == _T_408 ? welem[5] : _GEN_4166; // @[Execute.scala 117:10]
  assign _GEN_4168 = 6'h6 == _T_408 ? welem[6] : _GEN_4167; // @[Execute.scala 117:10]
  assign _GEN_4169 = 6'h7 == _T_408 ? welem[7] : _GEN_4168; // @[Execute.scala 117:10]
  assign _GEN_4170 = 6'h8 == _T_408 ? welem[8] : _GEN_4169; // @[Execute.scala 117:10]
  assign _GEN_4171 = 6'h9 == _T_408 ? welem[9] : _GEN_4170; // @[Execute.scala 117:10]
  assign _GEN_4172 = 6'ha == _T_408 ? welem[10] : _GEN_4171; // @[Execute.scala 117:10]
  assign _GEN_4173 = 6'hb == _T_408 ? welem[11] : _GEN_4172; // @[Execute.scala 117:10]
  assign _GEN_4174 = 6'hc == _T_408 ? welem[12] : _GEN_4173; // @[Execute.scala 117:10]
  assign _GEN_4175 = 6'hd == _T_408 ? welem[13] : _GEN_4174; // @[Execute.scala 117:10]
  assign _GEN_4176 = 6'he == _T_408 ? welem[14] : _GEN_4175; // @[Execute.scala 117:10]
  assign _GEN_4177 = 6'hf == _T_408 ? welem[15] : _GEN_4176; // @[Execute.scala 117:10]
  assign _GEN_4178 = 6'h10 == _T_408 ? welem[16] : _GEN_4177; // @[Execute.scala 117:10]
  assign _GEN_4179 = 6'h11 == _T_408 ? welem[17] : _GEN_4178; // @[Execute.scala 117:10]
  assign _GEN_4180 = 6'h12 == _T_408 ? welem[18] : _GEN_4179; // @[Execute.scala 117:10]
  assign _GEN_4181 = 6'h13 == _T_408 ? welem[19] : _GEN_4180; // @[Execute.scala 117:10]
  assign _GEN_4182 = 6'h14 == _T_408 ? welem[20] : _GEN_4181; // @[Execute.scala 117:10]
  assign _GEN_4183 = 6'h15 == _T_408 ? welem[21] : _GEN_4182; // @[Execute.scala 117:10]
  assign _GEN_4184 = 6'h16 == _T_408 ? welem[22] : _GEN_4183; // @[Execute.scala 117:10]
  assign _GEN_4185 = 6'h17 == _T_408 ? welem[23] : _GEN_4184; // @[Execute.scala 117:10]
  assign _GEN_4186 = 6'h18 == _T_408 ? welem[24] : _GEN_4185; // @[Execute.scala 117:10]
  assign _GEN_4187 = 6'h19 == _T_408 ? welem[25] : _GEN_4186; // @[Execute.scala 117:10]
  assign _GEN_4188 = 6'h1a == _T_408 ? welem[26] : _GEN_4187; // @[Execute.scala 117:10]
  assign _GEN_4189 = 6'h1b == _T_408 ? welem[27] : _GEN_4188; // @[Execute.scala 117:10]
  assign _GEN_4190 = 6'h1c == _T_408 ? welem[28] : _GEN_4189; // @[Execute.scala 117:10]
  assign _GEN_4191 = 6'h1d == _T_408 ? welem[29] : _GEN_4190; // @[Execute.scala 117:10]
  assign _GEN_4192 = 6'h1e == _T_408 ? welem[30] : _GEN_4191; // @[Execute.scala 117:10]
  assign _GEN_4193 = 6'h1f == _T_408 ? welem[31] : _GEN_4192; // @[Execute.scala 117:10]
  assign _GEN_4194 = 6'h20 == _T_408 ? welem[32] : _GEN_4193; // @[Execute.scala 117:10]
  assign _GEN_4195 = 6'h21 == _T_408 ? welem[33] : _GEN_4194; // @[Execute.scala 117:10]
  assign _GEN_4196 = 6'h22 == _T_408 ? welem[34] : _GEN_4195; // @[Execute.scala 117:10]
  assign _GEN_4197 = 6'h23 == _T_408 ? welem[35] : _GEN_4196; // @[Execute.scala 117:10]
  assign _GEN_4198 = 6'h24 == _T_408 ? welem[36] : _GEN_4197; // @[Execute.scala 117:10]
  assign _GEN_4199 = 6'h25 == _T_408 ? welem[37] : _GEN_4198; // @[Execute.scala 117:10]
  assign _GEN_4200 = 6'h26 == _T_408 ? welem[38] : _GEN_4199; // @[Execute.scala 117:10]
  assign _GEN_4201 = 6'h27 == _T_408 ? welem[39] : _GEN_4200; // @[Execute.scala 117:10]
  assign _GEN_4202 = 6'h28 == _T_408 ? welem[40] : _GEN_4201; // @[Execute.scala 117:10]
  assign _GEN_4203 = 6'h29 == _T_408 ? welem[41] : _GEN_4202; // @[Execute.scala 117:10]
  assign _GEN_4204 = 6'h2a == _T_408 ? welem[42] : _GEN_4203; // @[Execute.scala 117:10]
  assign _GEN_4205 = 6'h2b == _T_408 ? welem[43] : _GEN_4204; // @[Execute.scala 117:10]
  assign _GEN_4206 = 6'h2c == _T_408 ? welem[44] : _GEN_4205; // @[Execute.scala 117:10]
  assign _GEN_4207 = 6'h2d == _T_408 ? welem[45] : _GEN_4206; // @[Execute.scala 117:10]
  assign _GEN_4208 = 6'h2e == _T_408 ? welem[46] : _GEN_4207; // @[Execute.scala 117:10]
  assign _GEN_4209 = 6'h2f == _T_408 ? welem[47] : _GEN_4208; // @[Execute.scala 117:10]
  assign _GEN_4210 = 6'h30 == _T_408 ? welem[48] : _GEN_4209; // @[Execute.scala 117:10]
  assign _GEN_4211 = 6'h31 == _T_408 ? welem[49] : _GEN_4210; // @[Execute.scala 117:10]
  assign _GEN_4212 = 6'h32 == _T_408 ? welem[50] : _GEN_4211; // @[Execute.scala 117:10]
  assign _GEN_4213 = 6'h33 == _T_408 ? welem[51] : _GEN_4212; // @[Execute.scala 117:10]
  assign _GEN_4214 = 6'h34 == _T_408 ? welem[52] : _GEN_4213; // @[Execute.scala 117:10]
  assign _GEN_4215 = 6'h35 == _T_408 ? welem[53] : _GEN_4214; // @[Execute.scala 117:10]
  assign _GEN_4216 = 6'h36 == _T_408 ? welem[54] : _GEN_4215; // @[Execute.scala 117:10]
  assign _GEN_4217 = 6'h37 == _T_408 ? welem[55] : _GEN_4216; // @[Execute.scala 117:10]
  assign _GEN_4218 = 6'h38 == _T_408 ? welem[56] : _GEN_4217; // @[Execute.scala 117:10]
  assign _GEN_4219 = 6'h39 == _T_408 ? welem[57] : _GEN_4218; // @[Execute.scala 117:10]
  assign _GEN_4220 = 6'h3a == _T_408 ? welem[58] : _GEN_4219; // @[Execute.scala 117:10]
  assign _GEN_4221 = 6'h3b == _T_408 ? welem[59] : _GEN_4220; // @[Execute.scala 117:10]
  assign _GEN_4222 = 6'h3c == _T_408 ? welem[60] : _GEN_4221; // @[Execute.scala 117:10]
  assign _GEN_4223 = 6'h3d == _T_408 ? welem[61] : _GEN_4222; // @[Execute.scala 117:10]
  assign _GEN_4224 = 6'h3e == _T_408 ? welem[62] : _GEN_4223; // @[Execute.scala 117:10]
  assign _GEN_4225 = 6'h3f == _T_408 ? welem[63] : _GEN_4224; // @[Execute.scala 117:10]
  assign _T_411 = _T_402 ? _GEN_4161 : _GEN_4225; // @[Execute.scala 117:10]
  assign _T_412 = r < 6'h20; // @[Execute.scala 117:15]
  assign _T_414 = r - 6'h20; // @[Execute.scala 117:37]
  assign _T_418 = 6'h20 + r; // @[Execute.scala 117:60]
  assign _GEN_4227 = 6'h1 == _T_414 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4228 = 6'h2 == _T_414 ? welem[2] : _GEN_4227; // @[Execute.scala 117:10]
  assign _GEN_4229 = 6'h3 == _T_414 ? welem[3] : _GEN_4228; // @[Execute.scala 117:10]
  assign _GEN_4230 = 6'h4 == _T_414 ? welem[4] : _GEN_4229; // @[Execute.scala 117:10]
  assign _GEN_4231 = 6'h5 == _T_414 ? welem[5] : _GEN_4230; // @[Execute.scala 117:10]
  assign _GEN_4232 = 6'h6 == _T_414 ? welem[6] : _GEN_4231; // @[Execute.scala 117:10]
  assign _GEN_4233 = 6'h7 == _T_414 ? welem[7] : _GEN_4232; // @[Execute.scala 117:10]
  assign _GEN_4234 = 6'h8 == _T_414 ? welem[8] : _GEN_4233; // @[Execute.scala 117:10]
  assign _GEN_4235 = 6'h9 == _T_414 ? welem[9] : _GEN_4234; // @[Execute.scala 117:10]
  assign _GEN_4236 = 6'ha == _T_414 ? welem[10] : _GEN_4235; // @[Execute.scala 117:10]
  assign _GEN_4237 = 6'hb == _T_414 ? welem[11] : _GEN_4236; // @[Execute.scala 117:10]
  assign _GEN_4238 = 6'hc == _T_414 ? welem[12] : _GEN_4237; // @[Execute.scala 117:10]
  assign _GEN_4239 = 6'hd == _T_414 ? welem[13] : _GEN_4238; // @[Execute.scala 117:10]
  assign _GEN_4240 = 6'he == _T_414 ? welem[14] : _GEN_4239; // @[Execute.scala 117:10]
  assign _GEN_4241 = 6'hf == _T_414 ? welem[15] : _GEN_4240; // @[Execute.scala 117:10]
  assign _GEN_4242 = 6'h10 == _T_414 ? welem[16] : _GEN_4241; // @[Execute.scala 117:10]
  assign _GEN_4243 = 6'h11 == _T_414 ? welem[17] : _GEN_4242; // @[Execute.scala 117:10]
  assign _GEN_4244 = 6'h12 == _T_414 ? welem[18] : _GEN_4243; // @[Execute.scala 117:10]
  assign _GEN_4245 = 6'h13 == _T_414 ? welem[19] : _GEN_4244; // @[Execute.scala 117:10]
  assign _GEN_4246 = 6'h14 == _T_414 ? welem[20] : _GEN_4245; // @[Execute.scala 117:10]
  assign _GEN_4247 = 6'h15 == _T_414 ? welem[21] : _GEN_4246; // @[Execute.scala 117:10]
  assign _GEN_4248 = 6'h16 == _T_414 ? welem[22] : _GEN_4247; // @[Execute.scala 117:10]
  assign _GEN_4249 = 6'h17 == _T_414 ? welem[23] : _GEN_4248; // @[Execute.scala 117:10]
  assign _GEN_4250 = 6'h18 == _T_414 ? welem[24] : _GEN_4249; // @[Execute.scala 117:10]
  assign _GEN_4251 = 6'h19 == _T_414 ? welem[25] : _GEN_4250; // @[Execute.scala 117:10]
  assign _GEN_4252 = 6'h1a == _T_414 ? welem[26] : _GEN_4251; // @[Execute.scala 117:10]
  assign _GEN_4253 = 6'h1b == _T_414 ? welem[27] : _GEN_4252; // @[Execute.scala 117:10]
  assign _GEN_4254 = 6'h1c == _T_414 ? welem[28] : _GEN_4253; // @[Execute.scala 117:10]
  assign _GEN_4255 = 6'h1d == _T_414 ? welem[29] : _GEN_4254; // @[Execute.scala 117:10]
  assign _GEN_4256 = 6'h1e == _T_414 ? welem[30] : _GEN_4255; // @[Execute.scala 117:10]
  assign _GEN_4257 = 6'h1f == _T_414 ? welem[31] : _GEN_4256; // @[Execute.scala 117:10]
  assign _GEN_4258 = 6'h20 == _T_414 ? welem[32] : _GEN_4257; // @[Execute.scala 117:10]
  assign _GEN_4259 = 6'h21 == _T_414 ? welem[33] : _GEN_4258; // @[Execute.scala 117:10]
  assign _GEN_4260 = 6'h22 == _T_414 ? welem[34] : _GEN_4259; // @[Execute.scala 117:10]
  assign _GEN_4261 = 6'h23 == _T_414 ? welem[35] : _GEN_4260; // @[Execute.scala 117:10]
  assign _GEN_4262 = 6'h24 == _T_414 ? welem[36] : _GEN_4261; // @[Execute.scala 117:10]
  assign _GEN_4263 = 6'h25 == _T_414 ? welem[37] : _GEN_4262; // @[Execute.scala 117:10]
  assign _GEN_4264 = 6'h26 == _T_414 ? welem[38] : _GEN_4263; // @[Execute.scala 117:10]
  assign _GEN_4265 = 6'h27 == _T_414 ? welem[39] : _GEN_4264; // @[Execute.scala 117:10]
  assign _GEN_4266 = 6'h28 == _T_414 ? welem[40] : _GEN_4265; // @[Execute.scala 117:10]
  assign _GEN_4267 = 6'h29 == _T_414 ? welem[41] : _GEN_4266; // @[Execute.scala 117:10]
  assign _GEN_4268 = 6'h2a == _T_414 ? welem[42] : _GEN_4267; // @[Execute.scala 117:10]
  assign _GEN_4269 = 6'h2b == _T_414 ? welem[43] : _GEN_4268; // @[Execute.scala 117:10]
  assign _GEN_4270 = 6'h2c == _T_414 ? welem[44] : _GEN_4269; // @[Execute.scala 117:10]
  assign _GEN_4271 = 6'h2d == _T_414 ? welem[45] : _GEN_4270; // @[Execute.scala 117:10]
  assign _GEN_4272 = 6'h2e == _T_414 ? welem[46] : _GEN_4271; // @[Execute.scala 117:10]
  assign _GEN_4273 = 6'h2f == _T_414 ? welem[47] : _GEN_4272; // @[Execute.scala 117:10]
  assign _GEN_4274 = 6'h30 == _T_414 ? welem[48] : _GEN_4273; // @[Execute.scala 117:10]
  assign _GEN_4275 = 6'h31 == _T_414 ? welem[49] : _GEN_4274; // @[Execute.scala 117:10]
  assign _GEN_4276 = 6'h32 == _T_414 ? welem[50] : _GEN_4275; // @[Execute.scala 117:10]
  assign _GEN_4277 = 6'h33 == _T_414 ? welem[51] : _GEN_4276; // @[Execute.scala 117:10]
  assign _GEN_4278 = 6'h34 == _T_414 ? welem[52] : _GEN_4277; // @[Execute.scala 117:10]
  assign _GEN_4279 = 6'h35 == _T_414 ? welem[53] : _GEN_4278; // @[Execute.scala 117:10]
  assign _GEN_4280 = 6'h36 == _T_414 ? welem[54] : _GEN_4279; // @[Execute.scala 117:10]
  assign _GEN_4281 = 6'h37 == _T_414 ? welem[55] : _GEN_4280; // @[Execute.scala 117:10]
  assign _GEN_4282 = 6'h38 == _T_414 ? welem[56] : _GEN_4281; // @[Execute.scala 117:10]
  assign _GEN_4283 = 6'h39 == _T_414 ? welem[57] : _GEN_4282; // @[Execute.scala 117:10]
  assign _GEN_4284 = 6'h3a == _T_414 ? welem[58] : _GEN_4283; // @[Execute.scala 117:10]
  assign _GEN_4285 = 6'h3b == _T_414 ? welem[59] : _GEN_4284; // @[Execute.scala 117:10]
  assign _GEN_4286 = 6'h3c == _T_414 ? welem[60] : _GEN_4285; // @[Execute.scala 117:10]
  assign _GEN_4287 = 6'h3d == _T_414 ? welem[61] : _GEN_4286; // @[Execute.scala 117:10]
  assign _GEN_4288 = 6'h3e == _T_414 ? welem[62] : _GEN_4287; // @[Execute.scala 117:10]
  assign _GEN_4289 = 6'h3f == _T_414 ? welem[63] : _GEN_4288; // @[Execute.scala 117:10]
  assign _GEN_4291 = 6'h1 == _T_418 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4292 = 6'h2 == _T_418 ? welem[2] : _GEN_4291; // @[Execute.scala 117:10]
  assign _GEN_4293 = 6'h3 == _T_418 ? welem[3] : _GEN_4292; // @[Execute.scala 117:10]
  assign _GEN_4294 = 6'h4 == _T_418 ? welem[4] : _GEN_4293; // @[Execute.scala 117:10]
  assign _GEN_4295 = 6'h5 == _T_418 ? welem[5] : _GEN_4294; // @[Execute.scala 117:10]
  assign _GEN_4296 = 6'h6 == _T_418 ? welem[6] : _GEN_4295; // @[Execute.scala 117:10]
  assign _GEN_4297 = 6'h7 == _T_418 ? welem[7] : _GEN_4296; // @[Execute.scala 117:10]
  assign _GEN_4298 = 6'h8 == _T_418 ? welem[8] : _GEN_4297; // @[Execute.scala 117:10]
  assign _GEN_4299 = 6'h9 == _T_418 ? welem[9] : _GEN_4298; // @[Execute.scala 117:10]
  assign _GEN_4300 = 6'ha == _T_418 ? welem[10] : _GEN_4299; // @[Execute.scala 117:10]
  assign _GEN_4301 = 6'hb == _T_418 ? welem[11] : _GEN_4300; // @[Execute.scala 117:10]
  assign _GEN_4302 = 6'hc == _T_418 ? welem[12] : _GEN_4301; // @[Execute.scala 117:10]
  assign _GEN_4303 = 6'hd == _T_418 ? welem[13] : _GEN_4302; // @[Execute.scala 117:10]
  assign _GEN_4304 = 6'he == _T_418 ? welem[14] : _GEN_4303; // @[Execute.scala 117:10]
  assign _GEN_4305 = 6'hf == _T_418 ? welem[15] : _GEN_4304; // @[Execute.scala 117:10]
  assign _GEN_4306 = 6'h10 == _T_418 ? welem[16] : _GEN_4305; // @[Execute.scala 117:10]
  assign _GEN_4307 = 6'h11 == _T_418 ? welem[17] : _GEN_4306; // @[Execute.scala 117:10]
  assign _GEN_4308 = 6'h12 == _T_418 ? welem[18] : _GEN_4307; // @[Execute.scala 117:10]
  assign _GEN_4309 = 6'h13 == _T_418 ? welem[19] : _GEN_4308; // @[Execute.scala 117:10]
  assign _GEN_4310 = 6'h14 == _T_418 ? welem[20] : _GEN_4309; // @[Execute.scala 117:10]
  assign _GEN_4311 = 6'h15 == _T_418 ? welem[21] : _GEN_4310; // @[Execute.scala 117:10]
  assign _GEN_4312 = 6'h16 == _T_418 ? welem[22] : _GEN_4311; // @[Execute.scala 117:10]
  assign _GEN_4313 = 6'h17 == _T_418 ? welem[23] : _GEN_4312; // @[Execute.scala 117:10]
  assign _GEN_4314 = 6'h18 == _T_418 ? welem[24] : _GEN_4313; // @[Execute.scala 117:10]
  assign _GEN_4315 = 6'h19 == _T_418 ? welem[25] : _GEN_4314; // @[Execute.scala 117:10]
  assign _GEN_4316 = 6'h1a == _T_418 ? welem[26] : _GEN_4315; // @[Execute.scala 117:10]
  assign _GEN_4317 = 6'h1b == _T_418 ? welem[27] : _GEN_4316; // @[Execute.scala 117:10]
  assign _GEN_4318 = 6'h1c == _T_418 ? welem[28] : _GEN_4317; // @[Execute.scala 117:10]
  assign _GEN_4319 = 6'h1d == _T_418 ? welem[29] : _GEN_4318; // @[Execute.scala 117:10]
  assign _GEN_4320 = 6'h1e == _T_418 ? welem[30] : _GEN_4319; // @[Execute.scala 117:10]
  assign _GEN_4321 = 6'h1f == _T_418 ? welem[31] : _GEN_4320; // @[Execute.scala 117:10]
  assign _GEN_4322 = 6'h20 == _T_418 ? welem[32] : _GEN_4321; // @[Execute.scala 117:10]
  assign _GEN_4323 = 6'h21 == _T_418 ? welem[33] : _GEN_4322; // @[Execute.scala 117:10]
  assign _GEN_4324 = 6'h22 == _T_418 ? welem[34] : _GEN_4323; // @[Execute.scala 117:10]
  assign _GEN_4325 = 6'h23 == _T_418 ? welem[35] : _GEN_4324; // @[Execute.scala 117:10]
  assign _GEN_4326 = 6'h24 == _T_418 ? welem[36] : _GEN_4325; // @[Execute.scala 117:10]
  assign _GEN_4327 = 6'h25 == _T_418 ? welem[37] : _GEN_4326; // @[Execute.scala 117:10]
  assign _GEN_4328 = 6'h26 == _T_418 ? welem[38] : _GEN_4327; // @[Execute.scala 117:10]
  assign _GEN_4329 = 6'h27 == _T_418 ? welem[39] : _GEN_4328; // @[Execute.scala 117:10]
  assign _GEN_4330 = 6'h28 == _T_418 ? welem[40] : _GEN_4329; // @[Execute.scala 117:10]
  assign _GEN_4331 = 6'h29 == _T_418 ? welem[41] : _GEN_4330; // @[Execute.scala 117:10]
  assign _GEN_4332 = 6'h2a == _T_418 ? welem[42] : _GEN_4331; // @[Execute.scala 117:10]
  assign _GEN_4333 = 6'h2b == _T_418 ? welem[43] : _GEN_4332; // @[Execute.scala 117:10]
  assign _GEN_4334 = 6'h2c == _T_418 ? welem[44] : _GEN_4333; // @[Execute.scala 117:10]
  assign _GEN_4335 = 6'h2d == _T_418 ? welem[45] : _GEN_4334; // @[Execute.scala 117:10]
  assign _GEN_4336 = 6'h2e == _T_418 ? welem[46] : _GEN_4335; // @[Execute.scala 117:10]
  assign _GEN_4337 = 6'h2f == _T_418 ? welem[47] : _GEN_4336; // @[Execute.scala 117:10]
  assign _GEN_4338 = 6'h30 == _T_418 ? welem[48] : _GEN_4337; // @[Execute.scala 117:10]
  assign _GEN_4339 = 6'h31 == _T_418 ? welem[49] : _GEN_4338; // @[Execute.scala 117:10]
  assign _GEN_4340 = 6'h32 == _T_418 ? welem[50] : _GEN_4339; // @[Execute.scala 117:10]
  assign _GEN_4341 = 6'h33 == _T_418 ? welem[51] : _GEN_4340; // @[Execute.scala 117:10]
  assign _GEN_4342 = 6'h34 == _T_418 ? welem[52] : _GEN_4341; // @[Execute.scala 117:10]
  assign _GEN_4343 = 6'h35 == _T_418 ? welem[53] : _GEN_4342; // @[Execute.scala 117:10]
  assign _GEN_4344 = 6'h36 == _T_418 ? welem[54] : _GEN_4343; // @[Execute.scala 117:10]
  assign _GEN_4345 = 6'h37 == _T_418 ? welem[55] : _GEN_4344; // @[Execute.scala 117:10]
  assign _GEN_4346 = 6'h38 == _T_418 ? welem[56] : _GEN_4345; // @[Execute.scala 117:10]
  assign _GEN_4347 = 6'h39 == _T_418 ? welem[57] : _GEN_4346; // @[Execute.scala 117:10]
  assign _GEN_4348 = 6'h3a == _T_418 ? welem[58] : _GEN_4347; // @[Execute.scala 117:10]
  assign _GEN_4349 = 6'h3b == _T_418 ? welem[59] : _GEN_4348; // @[Execute.scala 117:10]
  assign _GEN_4350 = 6'h3c == _T_418 ? welem[60] : _GEN_4349; // @[Execute.scala 117:10]
  assign _GEN_4351 = 6'h3d == _T_418 ? welem[61] : _GEN_4350; // @[Execute.scala 117:10]
  assign _GEN_4352 = 6'h3e == _T_418 ? welem[62] : _GEN_4351; // @[Execute.scala 117:10]
  assign _GEN_4353 = 6'h3f == _T_418 ? welem[63] : _GEN_4352; // @[Execute.scala 117:10]
  assign _T_421 = _T_412 ? _GEN_4289 : _GEN_4353; // @[Execute.scala 117:10]
  assign _T_422 = r < 6'h1f; // @[Execute.scala 117:15]
  assign _T_424 = r - 6'h1f; // @[Execute.scala 117:37]
  assign _T_428 = 6'h21 + r; // @[Execute.scala 117:60]
  assign _GEN_4355 = 6'h1 == _T_424 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4356 = 6'h2 == _T_424 ? welem[2] : _GEN_4355; // @[Execute.scala 117:10]
  assign _GEN_4357 = 6'h3 == _T_424 ? welem[3] : _GEN_4356; // @[Execute.scala 117:10]
  assign _GEN_4358 = 6'h4 == _T_424 ? welem[4] : _GEN_4357; // @[Execute.scala 117:10]
  assign _GEN_4359 = 6'h5 == _T_424 ? welem[5] : _GEN_4358; // @[Execute.scala 117:10]
  assign _GEN_4360 = 6'h6 == _T_424 ? welem[6] : _GEN_4359; // @[Execute.scala 117:10]
  assign _GEN_4361 = 6'h7 == _T_424 ? welem[7] : _GEN_4360; // @[Execute.scala 117:10]
  assign _GEN_4362 = 6'h8 == _T_424 ? welem[8] : _GEN_4361; // @[Execute.scala 117:10]
  assign _GEN_4363 = 6'h9 == _T_424 ? welem[9] : _GEN_4362; // @[Execute.scala 117:10]
  assign _GEN_4364 = 6'ha == _T_424 ? welem[10] : _GEN_4363; // @[Execute.scala 117:10]
  assign _GEN_4365 = 6'hb == _T_424 ? welem[11] : _GEN_4364; // @[Execute.scala 117:10]
  assign _GEN_4366 = 6'hc == _T_424 ? welem[12] : _GEN_4365; // @[Execute.scala 117:10]
  assign _GEN_4367 = 6'hd == _T_424 ? welem[13] : _GEN_4366; // @[Execute.scala 117:10]
  assign _GEN_4368 = 6'he == _T_424 ? welem[14] : _GEN_4367; // @[Execute.scala 117:10]
  assign _GEN_4369 = 6'hf == _T_424 ? welem[15] : _GEN_4368; // @[Execute.scala 117:10]
  assign _GEN_4370 = 6'h10 == _T_424 ? welem[16] : _GEN_4369; // @[Execute.scala 117:10]
  assign _GEN_4371 = 6'h11 == _T_424 ? welem[17] : _GEN_4370; // @[Execute.scala 117:10]
  assign _GEN_4372 = 6'h12 == _T_424 ? welem[18] : _GEN_4371; // @[Execute.scala 117:10]
  assign _GEN_4373 = 6'h13 == _T_424 ? welem[19] : _GEN_4372; // @[Execute.scala 117:10]
  assign _GEN_4374 = 6'h14 == _T_424 ? welem[20] : _GEN_4373; // @[Execute.scala 117:10]
  assign _GEN_4375 = 6'h15 == _T_424 ? welem[21] : _GEN_4374; // @[Execute.scala 117:10]
  assign _GEN_4376 = 6'h16 == _T_424 ? welem[22] : _GEN_4375; // @[Execute.scala 117:10]
  assign _GEN_4377 = 6'h17 == _T_424 ? welem[23] : _GEN_4376; // @[Execute.scala 117:10]
  assign _GEN_4378 = 6'h18 == _T_424 ? welem[24] : _GEN_4377; // @[Execute.scala 117:10]
  assign _GEN_4379 = 6'h19 == _T_424 ? welem[25] : _GEN_4378; // @[Execute.scala 117:10]
  assign _GEN_4380 = 6'h1a == _T_424 ? welem[26] : _GEN_4379; // @[Execute.scala 117:10]
  assign _GEN_4381 = 6'h1b == _T_424 ? welem[27] : _GEN_4380; // @[Execute.scala 117:10]
  assign _GEN_4382 = 6'h1c == _T_424 ? welem[28] : _GEN_4381; // @[Execute.scala 117:10]
  assign _GEN_4383 = 6'h1d == _T_424 ? welem[29] : _GEN_4382; // @[Execute.scala 117:10]
  assign _GEN_4384 = 6'h1e == _T_424 ? welem[30] : _GEN_4383; // @[Execute.scala 117:10]
  assign _GEN_4385 = 6'h1f == _T_424 ? welem[31] : _GEN_4384; // @[Execute.scala 117:10]
  assign _GEN_4386 = 6'h20 == _T_424 ? welem[32] : _GEN_4385; // @[Execute.scala 117:10]
  assign _GEN_4387 = 6'h21 == _T_424 ? welem[33] : _GEN_4386; // @[Execute.scala 117:10]
  assign _GEN_4388 = 6'h22 == _T_424 ? welem[34] : _GEN_4387; // @[Execute.scala 117:10]
  assign _GEN_4389 = 6'h23 == _T_424 ? welem[35] : _GEN_4388; // @[Execute.scala 117:10]
  assign _GEN_4390 = 6'h24 == _T_424 ? welem[36] : _GEN_4389; // @[Execute.scala 117:10]
  assign _GEN_4391 = 6'h25 == _T_424 ? welem[37] : _GEN_4390; // @[Execute.scala 117:10]
  assign _GEN_4392 = 6'h26 == _T_424 ? welem[38] : _GEN_4391; // @[Execute.scala 117:10]
  assign _GEN_4393 = 6'h27 == _T_424 ? welem[39] : _GEN_4392; // @[Execute.scala 117:10]
  assign _GEN_4394 = 6'h28 == _T_424 ? welem[40] : _GEN_4393; // @[Execute.scala 117:10]
  assign _GEN_4395 = 6'h29 == _T_424 ? welem[41] : _GEN_4394; // @[Execute.scala 117:10]
  assign _GEN_4396 = 6'h2a == _T_424 ? welem[42] : _GEN_4395; // @[Execute.scala 117:10]
  assign _GEN_4397 = 6'h2b == _T_424 ? welem[43] : _GEN_4396; // @[Execute.scala 117:10]
  assign _GEN_4398 = 6'h2c == _T_424 ? welem[44] : _GEN_4397; // @[Execute.scala 117:10]
  assign _GEN_4399 = 6'h2d == _T_424 ? welem[45] : _GEN_4398; // @[Execute.scala 117:10]
  assign _GEN_4400 = 6'h2e == _T_424 ? welem[46] : _GEN_4399; // @[Execute.scala 117:10]
  assign _GEN_4401 = 6'h2f == _T_424 ? welem[47] : _GEN_4400; // @[Execute.scala 117:10]
  assign _GEN_4402 = 6'h30 == _T_424 ? welem[48] : _GEN_4401; // @[Execute.scala 117:10]
  assign _GEN_4403 = 6'h31 == _T_424 ? welem[49] : _GEN_4402; // @[Execute.scala 117:10]
  assign _GEN_4404 = 6'h32 == _T_424 ? welem[50] : _GEN_4403; // @[Execute.scala 117:10]
  assign _GEN_4405 = 6'h33 == _T_424 ? welem[51] : _GEN_4404; // @[Execute.scala 117:10]
  assign _GEN_4406 = 6'h34 == _T_424 ? welem[52] : _GEN_4405; // @[Execute.scala 117:10]
  assign _GEN_4407 = 6'h35 == _T_424 ? welem[53] : _GEN_4406; // @[Execute.scala 117:10]
  assign _GEN_4408 = 6'h36 == _T_424 ? welem[54] : _GEN_4407; // @[Execute.scala 117:10]
  assign _GEN_4409 = 6'h37 == _T_424 ? welem[55] : _GEN_4408; // @[Execute.scala 117:10]
  assign _GEN_4410 = 6'h38 == _T_424 ? welem[56] : _GEN_4409; // @[Execute.scala 117:10]
  assign _GEN_4411 = 6'h39 == _T_424 ? welem[57] : _GEN_4410; // @[Execute.scala 117:10]
  assign _GEN_4412 = 6'h3a == _T_424 ? welem[58] : _GEN_4411; // @[Execute.scala 117:10]
  assign _GEN_4413 = 6'h3b == _T_424 ? welem[59] : _GEN_4412; // @[Execute.scala 117:10]
  assign _GEN_4414 = 6'h3c == _T_424 ? welem[60] : _GEN_4413; // @[Execute.scala 117:10]
  assign _GEN_4415 = 6'h3d == _T_424 ? welem[61] : _GEN_4414; // @[Execute.scala 117:10]
  assign _GEN_4416 = 6'h3e == _T_424 ? welem[62] : _GEN_4415; // @[Execute.scala 117:10]
  assign _GEN_4417 = 6'h3f == _T_424 ? welem[63] : _GEN_4416; // @[Execute.scala 117:10]
  assign _GEN_4419 = 6'h1 == _T_428 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4420 = 6'h2 == _T_428 ? welem[2] : _GEN_4419; // @[Execute.scala 117:10]
  assign _GEN_4421 = 6'h3 == _T_428 ? welem[3] : _GEN_4420; // @[Execute.scala 117:10]
  assign _GEN_4422 = 6'h4 == _T_428 ? welem[4] : _GEN_4421; // @[Execute.scala 117:10]
  assign _GEN_4423 = 6'h5 == _T_428 ? welem[5] : _GEN_4422; // @[Execute.scala 117:10]
  assign _GEN_4424 = 6'h6 == _T_428 ? welem[6] : _GEN_4423; // @[Execute.scala 117:10]
  assign _GEN_4425 = 6'h7 == _T_428 ? welem[7] : _GEN_4424; // @[Execute.scala 117:10]
  assign _GEN_4426 = 6'h8 == _T_428 ? welem[8] : _GEN_4425; // @[Execute.scala 117:10]
  assign _GEN_4427 = 6'h9 == _T_428 ? welem[9] : _GEN_4426; // @[Execute.scala 117:10]
  assign _GEN_4428 = 6'ha == _T_428 ? welem[10] : _GEN_4427; // @[Execute.scala 117:10]
  assign _GEN_4429 = 6'hb == _T_428 ? welem[11] : _GEN_4428; // @[Execute.scala 117:10]
  assign _GEN_4430 = 6'hc == _T_428 ? welem[12] : _GEN_4429; // @[Execute.scala 117:10]
  assign _GEN_4431 = 6'hd == _T_428 ? welem[13] : _GEN_4430; // @[Execute.scala 117:10]
  assign _GEN_4432 = 6'he == _T_428 ? welem[14] : _GEN_4431; // @[Execute.scala 117:10]
  assign _GEN_4433 = 6'hf == _T_428 ? welem[15] : _GEN_4432; // @[Execute.scala 117:10]
  assign _GEN_4434 = 6'h10 == _T_428 ? welem[16] : _GEN_4433; // @[Execute.scala 117:10]
  assign _GEN_4435 = 6'h11 == _T_428 ? welem[17] : _GEN_4434; // @[Execute.scala 117:10]
  assign _GEN_4436 = 6'h12 == _T_428 ? welem[18] : _GEN_4435; // @[Execute.scala 117:10]
  assign _GEN_4437 = 6'h13 == _T_428 ? welem[19] : _GEN_4436; // @[Execute.scala 117:10]
  assign _GEN_4438 = 6'h14 == _T_428 ? welem[20] : _GEN_4437; // @[Execute.scala 117:10]
  assign _GEN_4439 = 6'h15 == _T_428 ? welem[21] : _GEN_4438; // @[Execute.scala 117:10]
  assign _GEN_4440 = 6'h16 == _T_428 ? welem[22] : _GEN_4439; // @[Execute.scala 117:10]
  assign _GEN_4441 = 6'h17 == _T_428 ? welem[23] : _GEN_4440; // @[Execute.scala 117:10]
  assign _GEN_4442 = 6'h18 == _T_428 ? welem[24] : _GEN_4441; // @[Execute.scala 117:10]
  assign _GEN_4443 = 6'h19 == _T_428 ? welem[25] : _GEN_4442; // @[Execute.scala 117:10]
  assign _GEN_4444 = 6'h1a == _T_428 ? welem[26] : _GEN_4443; // @[Execute.scala 117:10]
  assign _GEN_4445 = 6'h1b == _T_428 ? welem[27] : _GEN_4444; // @[Execute.scala 117:10]
  assign _GEN_4446 = 6'h1c == _T_428 ? welem[28] : _GEN_4445; // @[Execute.scala 117:10]
  assign _GEN_4447 = 6'h1d == _T_428 ? welem[29] : _GEN_4446; // @[Execute.scala 117:10]
  assign _GEN_4448 = 6'h1e == _T_428 ? welem[30] : _GEN_4447; // @[Execute.scala 117:10]
  assign _GEN_4449 = 6'h1f == _T_428 ? welem[31] : _GEN_4448; // @[Execute.scala 117:10]
  assign _GEN_4450 = 6'h20 == _T_428 ? welem[32] : _GEN_4449; // @[Execute.scala 117:10]
  assign _GEN_4451 = 6'h21 == _T_428 ? welem[33] : _GEN_4450; // @[Execute.scala 117:10]
  assign _GEN_4452 = 6'h22 == _T_428 ? welem[34] : _GEN_4451; // @[Execute.scala 117:10]
  assign _GEN_4453 = 6'h23 == _T_428 ? welem[35] : _GEN_4452; // @[Execute.scala 117:10]
  assign _GEN_4454 = 6'h24 == _T_428 ? welem[36] : _GEN_4453; // @[Execute.scala 117:10]
  assign _GEN_4455 = 6'h25 == _T_428 ? welem[37] : _GEN_4454; // @[Execute.scala 117:10]
  assign _GEN_4456 = 6'h26 == _T_428 ? welem[38] : _GEN_4455; // @[Execute.scala 117:10]
  assign _GEN_4457 = 6'h27 == _T_428 ? welem[39] : _GEN_4456; // @[Execute.scala 117:10]
  assign _GEN_4458 = 6'h28 == _T_428 ? welem[40] : _GEN_4457; // @[Execute.scala 117:10]
  assign _GEN_4459 = 6'h29 == _T_428 ? welem[41] : _GEN_4458; // @[Execute.scala 117:10]
  assign _GEN_4460 = 6'h2a == _T_428 ? welem[42] : _GEN_4459; // @[Execute.scala 117:10]
  assign _GEN_4461 = 6'h2b == _T_428 ? welem[43] : _GEN_4460; // @[Execute.scala 117:10]
  assign _GEN_4462 = 6'h2c == _T_428 ? welem[44] : _GEN_4461; // @[Execute.scala 117:10]
  assign _GEN_4463 = 6'h2d == _T_428 ? welem[45] : _GEN_4462; // @[Execute.scala 117:10]
  assign _GEN_4464 = 6'h2e == _T_428 ? welem[46] : _GEN_4463; // @[Execute.scala 117:10]
  assign _GEN_4465 = 6'h2f == _T_428 ? welem[47] : _GEN_4464; // @[Execute.scala 117:10]
  assign _GEN_4466 = 6'h30 == _T_428 ? welem[48] : _GEN_4465; // @[Execute.scala 117:10]
  assign _GEN_4467 = 6'h31 == _T_428 ? welem[49] : _GEN_4466; // @[Execute.scala 117:10]
  assign _GEN_4468 = 6'h32 == _T_428 ? welem[50] : _GEN_4467; // @[Execute.scala 117:10]
  assign _GEN_4469 = 6'h33 == _T_428 ? welem[51] : _GEN_4468; // @[Execute.scala 117:10]
  assign _GEN_4470 = 6'h34 == _T_428 ? welem[52] : _GEN_4469; // @[Execute.scala 117:10]
  assign _GEN_4471 = 6'h35 == _T_428 ? welem[53] : _GEN_4470; // @[Execute.scala 117:10]
  assign _GEN_4472 = 6'h36 == _T_428 ? welem[54] : _GEN_4471; // @[Execute.scala 117:10]
  assign _GEN_4473 = 6'h37 == _T_428 ? welem[55] : _GEN_4472; // @[Execute.scala 117:10]
  assign _GEN_4474 = 6'h38 == _T_428 ? welem[56] : _GEN_4473; // @[Execute.scala 117:10]
  assign _GEN_4475 = 6'h39 == _T_428 ? welem[57] : _GEN_4474; // @[Execute.scala 117:10]
  assign _GEN_4476 = 6'h3a == _T_428 ? welem[58] : _GEN_4475; // @[Execute.scala 117:10]
  assign _GEN_4477 = 6'h3b == _T_428 ? welem[59] : _GEN_4476; // @[Execute.scala 117:10]
  assign _GEN_4478 = 6'h3c == _T_428 ? welem[60] : _GEN_4477; // @[Execute.scala 117:10]
  assign _GEN_4479 = 6'h3d == _T_428 ? welem[61] : _GEN_4478; // @[Execute.scala 117:10]
  assign _GEN_4480 = 6'h3e == _T_428 ? welem[62] : _GEN_4479; // @[Execute.scala 117:10]
  assign _GEN_4481 = 6'h3f == _T_428 ? welem[63] : _GEN_4480; // @[Execute.scala 117:10]
  assign _T_431 = _T_422 ? _GEN_4417 : _GEN_4481; // @[Execute.scala 117:10]
  assign _T_432 = r < 6'h1e; // @[Execute.scala 117:15]
  assign _T_434 = r - 6'h1e; // @[Execute.scala 117:37]
  assign _T_438 = 6'h22 + r; // @[Execute.scala 117:60]
  assign _GEN_4483 = 6'h1 == _T_434 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4484 = 6'h2 == _T_434 ? welem[2] : _GEN_4483; // @[Execute.scala 117:10]
  assign _GEN_4485 = 6'h3 == _T_434 ? welem[3] : _GEN_4484; // @[Execute.scala 117:10]
  assign _GEN_4486 = 6'h4 == _T_434 ? welem[4] : _GEN_4485; // @[Execute.scala 117:10]
  assign _GEN_4487 = 6'h5 == _T_434 ? welem[5] : _GEN_4486; // @[Execute.scala 117:10]
  assign _GEN_4488 = 6'h6 == _T_434 ? welem[6] : _GEN_4487; // @[Execute.scala 117:10]
  assign _GEN_4489 = 6'h7 == _T_434 ? welem[7] : _GEN_4488; // @[Execute.scala 117:10]
  assign _GEN_4490 = 6'h8 == _T_434 ? welem[8] : _GEN_4489; // @[Execute.scala 117:10]
  assign _GEN_4491 = 6'h9 == _T_434 ? welem[9] : _GEN_4490; // @[Execute.scala 117:10]
  assign _GEN_4492 = 6'ha == _T_434 ? welem[10] : _GEN_4491; // @[Execute.scala 117:10]
  assign _GEN_4493 = 6'hb == _T_434 ? welem[11] : _GEN_4492; // @[Execute.scala 117:10]
  assign _GEN_4494 = 6'hc == _T_434 ? welem[12] : _GEN_4493; // @[Execute.scala 117:10]
  assign _GEN_4495 = 6'hd == _T_434 ? welem[13] : _GEN_4494; // @[Execute.scala 117:10]
  assign _GEN_4496 = 6'he == _T_434 ? welem[14] : _GEN_4495; // @[Execute.scala 117:10]
  assign _GEN_4497 = 6'hf == _T_434 ? welem[15] : _GEN_4496; // @[Execute.scala 117:10]
  assign _GEN_4498 = 6'h10 == _T_434 ? welem[16] : _GEN_4497; // @[Execute.scala 117:10]
  assign _GEN_4499 = 6'h11 == _T_434 ? welem[17] : _GEN_4498; // @[Execute.scala 117:10]
  assign _GEN_4500 = 6'h12 == _T_434 ? welem[18] : _GEN_4499; // @[Execute.scala 117:10]
  assign _GEN_4501 = 6'h13 == _T_434 ? welem[19] : _GEN_4500; // @[Execute.scala 117:10]
  assign _GEN_4502 = 6'h14 == _T_434 ? welem[20] : _GEN_4501; // @[Execute.scala 117:10]
  assign _GEN_4503 = 6'h15 == _T_434 ? welem[21] : _GEN_4502; // @[Execute.scala 117:10]
  assign _GEN_4504 = 6'h16 == _T_434 ? welem[22] : _GEN_4503; // @[Execute.scala 117:10]
  assign _GEN_4505 = 6'h17 == _T_434 ? welem[23] : _GEN_4504; // @[Execute.scala 117:10]
  assign _GEN_4506 = 6'h18 == _T_434 ? welem[24] : _GEN_4505; // @[Execute.scala 117:10]
  assign _GEN_4507 = 6'h19 == _T_434 ? welem[25] : _GEN_4506; // @[Execute.scala 117:10]
  assign _GEN_4508 = 6'h1a == _T_434 ? welem[26] : _GEN_4507; // @[Execute.scala 117:10]
  assign _GEN_4509 = 6'h1b == _T_434 ? welem[27] : _GEN_4508; // @[Execute.scala 117:10]
  assign _GEN_4510 = 6'h1c == _T_434 ? welem[28] : _GEN_4509; // @[Execute.scala 117:10]
  assign _GEN_4511 = 6'h1d == _T_434 ? welem[29] : _GEN_4510; // @[Execute.scala 117:10]
  assign _GEN_4512 = 6'h1e == _T_434 ? welem[30] : _GEN_4511; // @[Execute.scala 117:10]
  assign _GEN_4513 = 6'h1f == _T_434 ? welem[31] : _GEN_4512; // @[Execute.scala 117:10]
  assign _GEN_4514 = 6'h20 == _T_434 ? welem[32] : _GEN_4513; // @[Execute.scala 117:10]
  assign _GEN_4515 = 6'h21 == _T_434 ? welem[33] : _GEN_4514; // @[Execute.scala 117:10]
  assign _GEN_4516 = 6'h22 == _T_434 ? welem[34] : _GEN_4515; // @[Execute.scala 117:10]
  assign _GEN_4517 = 6'h23 == _T_434 ? welem[35] : _GEN_4516; // @[Execute.scala 117:10]
  assign _GEN_4518 = 6'h24 == _T_434 ? welem[36] : _GEN_4517; // @[Execute.scala 117:10]
  assign _GEN_4519 = 6'h25 == _T_434 ? welem[37] : _GEN_4518; // @[Execute.scala 117:10]
  assign _GEN_4520 = 6'h26 == _T_434 ? welem[38] : _GEN_4519; // @[Execute.scala 117:10]
  assign _GEN_4521 = 6'h27 == _T_434 ? welem[39] : _GEN_4520; // @[Execute.scala 117:10]
  assign _GEN_4522 = 6'h28 == _T_434 ? welem[40] : _GEN_4521; // @[Execute.scala 117:10]
  assign _GEN_4523 = 6'h29 == _T_434 ? welem[41] : _GEN_4522; // @[Execute.scala 117:10]
  assign _GEN_4524 = 6'h2a == _T_434 ? welem[42] : _GEN_4523; // @[Execute.scala 117:10]
  assign _GEN_4525 = 6'h2b == _T_434 ? welem[43] : _GEN_4524; // @[Execute.scala 117:10]
  assign _GEN_4526 = 6'h2c == _T_434 ? welem[44] : _GEN_4525; // @[Execute.scala 117:10]
  assign _GEN_4527 = 6'h2d == _T_434 ? welem[45] : _GEN_4526; // @[Execute.scala 117:10]
  assign _GEN_4528 = 6'h2e == _T_434 ? welem[46] : _GEN_4527; // @[Execute.scala 117:10]
  assign _GEN_4529 = 6'h2f == _T_434 ? welem[47] : _GEN_4528; // @[Execute.scala 117:10]
  assign _GEN_4530 = 6'h30 == _T_434 ? welem[48] : _GEN_4529; // @[Execute.scala 117:10]
  assign _GEN_4531 = 6'h31 == _T_434 ? welem[49] : _GEN_4530; // @[Execute.scala 117:10]
  assign _GEN_4532 = 6'h32 == _T_434 ? welem[50] : _GEN_4531; // @[Execute.scala 117:10]
  assign _GEN_4533 = 6'h33 == _T_434 ? welem[51] : _GEN_4532; // @[Execute.scala 117:10]
  assign _GEN_4534 = 6'h34 == _T_434 ? welem[52] : _GEN_4533; // @[Execute.scala 117:10]
  assign _GEN_4535 = 6'h35 == _T_434 ? welem[53] : _GEN_4534; // @[Execute.scala 117:10]
  assign _GEN_4536 = 6'h36 == _T_434 ? welem[54] : _GEN_4535; // @[Execute.scala 117:10]
  assign _GEN_4537 = 6'h37 == _T_434 ? welem[55] : _GEN_4536; // @[Execute.scala 117:10]
  assign _GEN_4538 = 6'h38 == _T_434 ? welem[56] : _GEN_4537; // @[Execute.scala 117:10]
  assign _GEN_4539 = 6'h39 == _T_434 ? welem[57] : _GEN_4538; // @[Execute.scala 117:10]
  assign _GEN_4540 = 6'h3a == _T_434 ? welem[58] : _GEN_4539; // @[Execute.scala 117:10]
  assign _GEN_4541 = 6'h3b == _T_434 ? welem[59] : _GEN_4540; // @[Execute.scala 117:10]
  assign _GEN_4542 = 6'h3c == _T_434 ? welem[60] : _GEN_4541; // @[Execute.scala 117:10]
  assign _GEN_4543 = 6'h3d == _T_434 ? welem[61] : _GEN_4542; // @[Execute.scala 117:10]
  assign _GEN_4544 = 6'h3e == _T_434 ? welem[62] : _GEN_4543; // @[Execute.scala 117:10]
  assign _GEN_4545 = 6'h3f == _T_434 ? welem[63] : _GEN_4544; // @[Execute.scala 117:10]
  assign _GEN_4547 = 6'h1 == _T_438 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4548 = 6'h2 == _T_438 ? welem[2] : _GEN_4547; // @[Execute.scala 117:10]
  assign _GEN_4549 = 6'h3 == _T_438 ? welem[3] : _GEN_4548; // @[Execute.scala 117:10]
  assign _GEN_4550 = 6'h4 == _T_438 ? welem[4] : _GEN_4549; // @[Execute.scala 117:10]
  assign _GEN_4551 = 6'h5 == _T_438 ? welem[5] : _GEN_4550; // @[Execute.scala 117:10]
  assign _GEN_4552 = 6'h6 == _T_438 ? welem[6] : _GEN_4551; // @[Execute.scala 117:10]
  assign _GEN_4553 = 6'h7 == _T_438 ? welem[7] : _GEN_4552; // @[Execute.scala 117:10]
  assign _GEN_4554 = 6'h8 == _T_438 ? welem[8] : _GEN_4553; // @[Execute.scala 117:10]
  assign _GEN_4555 = 6'h9 == _T_438 ? welem[9] : _GEN_4554; // @[Execute.scala 117:10]
  assign _GEN_4556 = 6'ha == _T_438 ? welem[10] : _GEN_4555; // @[Execute.scala 117:10]
  assign _GEN_4557 = 6'hb == _T_438 ? welem[11] : _GEN_4556; // @[Execute.scala 117:10]
  assign _GEN_4558 = 6'hc == _T_438 ? welem[12] : _GEN_4557; // @[Execute.scala 117:10]
  assign _GEN_4559 = 6'hd == _T_438 ? welem[13] : _GEN_4558; // @[Execute.scala 117:10]
  assign _GEN_4560 = 6'he == _T_438 ? welem[14] : _GEN_4559; // @[Execute.scala 117:10]
  assign _GEN_4561 = 6'hf == _T_438 ? welem[15] : _GEN_4560; // @[Execute.scala 117:10]
  assign _GEN_4562 = 6'h10 == _T_438 ? welem[16] : _GEN_4561; // @[Execute.scala 117:10]
  assign _GEN_4563 = 6'h11 == _T_438 ? welem[17] : _GEN_4562; // @[Execute.scala 117:10]
  assign _GEN_4564 = 6'h12 == _T_438 ? welem[18] : _GEN_4563; // @[Execute.scala 117:10]
  assign _GEN_4565 = 6'h13 == _T_438 ? welem[19] : _GEN_4564; // @[Execute.scala 117:10]
  assign _GEN_4566 = 6'h14 == _T_438 ? welem[20] : _GEN_4565; // @[Execute.scala 117:10]
  assign _GEN_4567 = 6'h15 == _T_438 ? welem[21] : _GEN_4566; // @[Execute.scala 117:10]
  assign _GEN_4568 = 6'h16 == _T_438 ? welem[22] : _GEN_4567; // @[Execute.scala 117:10]
  assign _GEN_4569 = 6'h17 == _T_438 ? welem[23] : _GEN_4568; // @[Execute.scala 117:10]
  assign _GEN_4570 = 6'h18 == _T_438 ? welem[24] : _GEN_4569; // @[Execute.scala 117:10]
  assign _GEN_4571 = 6'h19 == _T_438 ? welem[25] : _GEN_4570; // @[Execute.scala 117:10]
  assign _GEN_4572 = 6'h1a == _T_438 ? welem[26] : _GEN_4571; // @[Execute.scala 117:10]
  assign _GEN_4573 = 6'h1b == _T_438 ? welem[27] : _GEN_4572; // @[Execute.scala 117:10]
  assign _GEN_4574 = 6'h1c == _T_438 ? welem[28] : _GEN_4573; // @[Execute.scala 117:10]
  assign _GEN_4575 = 6'h1d == _T_438 ? welem[29] : _GEN_4574; // @[Execute.scala 117:10]
  assign _GEN_4576 = 6'h1e == _T_438 ? welem[30] : _GEN_4575; // @[Execute.scala 117:10]
  assign _GEN_4577 = 6'h1f == _T_438 ? welem[31] : _GEN_4576; // @[Execute.scala 117:10]
  assign _GEN_4578 = 6'h20 == _T_438 ? welem[32] : _GEN_4577; // @[Execute.scala 117:10]
  assign _GEN_4579 = 6'h21 == _T_438 ? welem[33] : _GEN_4578; // @[Execute.scala 117:10]
  assign _GEN_4580 = 6'h22 == _T_438 ? welem[34] : _GEN_4579; // @[Execute.scala 117:10]
  assign _GEN_4581 = 6'h23 == _T_438 ? welem[35] : _GEN_4580; // @[Execute.scala 117:10]
  assign _GEN_4582 = 6'h24 == _T_438 ? welem[36] : _GEN_4581; // @[Execute.scala 117:10]
  assign _GEN_4583 = 6'h25 == _T_438 ? welem[37] : _GEN_4582; // @[Execute.scala 117:10]
  assign _GEN_4584 = 6'h26 == _T_438 ? welem[38] : _GEN_4583; // @[Execute.scala 117:10]
  assign _GEN_4585 = 6'h27 == _T_438 ? welem[39] : _GEN_4584; // @[Execute.scala 117:10]
  assign _GEN_4586 = 6'h28 == _T_438 ? welem[40] : _GEN_4585; // @[Execute.scala 117:10]
  assign _GEN_4587 = 6'h29 == _T_438 ? welem[41] : _GEN_4586; // @[Execute.scala 117:10]
  assign _GEN_4588 = 6'h2a == _T_438 ? welem[42] : _GEN_4587; // @[Execute.scala 117:10]
  assign _GEN_4589 = 6'h2b == _T_438 ? welem[43] : _GEN_4588; // @[Execute.scala 117:10]
  assign _GEN_4590 = 6'h2c == _T_438 ? welem[44] : _GEN_4589; // @[Execute.scala 117:10]
  assign _GEN_4591 = 6'h2d == _T_438 ? welem[45] : _GEN_4590; // @[Execute.scala 117:10]
  assign _GEN_4592 = 6'h2e == _T_438 ? welem[46] : _GEN_4591; // @[Execute.scala 117:10]
  assign _GEN_4593 = 6'h2f == _T_438 ? welem[47] : _GEN_4592; // @[Execute.scala 117:10]
  assign _GEN_4594 = 6'h30 == _T_438 ? welem[48] : _GEN_4593; // @[Execute.scala 117:10]
  assign _GEN_4595 = 6'h31 == _T_438 ? welem[49] : _GEN_4594; // @[Execute.scala 117:10]
  assign _GEN_4596 = 6'h32 == _T_438 ? welem[50] : _GEN_4595; // @[Execute.scala 117:10]
  assign _GEN_4597 = 6'h33 == _T_438 ? welem[51] : _GEN_4596; // @[Execute.scala 117:10]
  assign _GEN_4598 = 6'h34 == _T_438 ? welem[52] : _GEN_4597; // @[Execute.scala 117:10]
  assign _GEN_4599 = 6'h35 == _T_438 ? welem[53] : _GEN_4598; // @[Execute.scala 117:10]
  assign _GEN_4600 = 6'h36 == _T_438 ? welem[54] : _GEN_4599; // @[Execute.scala 117:10]
  assign _GEN_4601 = 6'h37 == _T_438 ? welem[55] : _GEN_4600; // @[Execute.scala 117:10]
  assign _GEN_4602 = 6'h38 == _T_438 ? welem[56] : _GEN_4601; // @[Execute.scala 117:10]
  assign _GEN_4603 = 6'h39 == _T_438 ? welem[57] : _GEN_4602; // @[Execute.scala 117:10]
  assign _GEN_4604 = 6'h3a == _T_438 ? welem[58] : _GEN_4603; // @[Execute.scala 117:10]
  assign _GEN_4605 = 6'h3b == _T_438 ? welem[59] : _GEN_4604; // @[Execute.scala 117:10]
  assign _GEN_4606 = 6'h3c == _T_438 ? welem[60] : _GEN_4605; // @[Execute.scala 117:10]
  assign _GEN_4607 = 6'h3d == _T_438 ? welem[61] : _GEN_4606; // @[Execute.scala 117:10]
  assign _GEN_4608 = 6'h3e == _T_438 ? welem[62] : _GEN_4607; // @[Execute.scala 117:10]
  assign _GEN_4609 = 6'h3f == _T_438 ? welem[63] : _GEN_4608; // @[Execute.scala 117:10]
  assign _T_441 = _T_432 ? _GEN_4545 : _GEN_4609; // @[Execute.scala 117:10]
  assign _T_442 = r < 6'h1d; // @[Execute.scala 117:15]
  assign _T_444 = r - 6'h1d; // @[Execute.scala 117:37]
  assign _T_448 = 6'h23 + r; // @[Execute.scala 117:60]
  assign _GEN_4611 = 6'h1 == _T_444 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4612 = 6'h2 == _T_444 ? welem[2] : _GEN_4611; // @[Execute.scala 117:10]
  assign _GEN_4613 = 6'h3 == _T_444 ? welem[3] : _GEN_4612; // @[Execute.scala 117:10]
  assign _GEN_4614 = 6'h4 == _T_444 ? welem[4] : _GEN_4613; // @[Execute.scala 117:10]
  assign _GEN_4615 = 6'h5 == _T_444 ? welem[5] : _GEN_4614; // @[Execute.scala 117:10]
  assign _GEN_4616 = 6'h6 == _T_444 ? welem[6] : _GEN_4615; // @[Execute.scala 117:10]
  assign _GEN_4617 = 6'h7 == _T_444 ? welem[7] : _GEN_4616; // @[Execute.scala 117:10]
  assign _GEN_4618 = 6'h8 == _T_444 ? welem[8] : _GEN_4617; // @[Execute.scala 117:10]
  assign _GEN_4619 = 6'h9 == _T_444 ? welem[9] : _GEN_4618; // @[Execute.scala 117:10]
  assign _GEN_4620 = 6'ha == _T_444 ? welem[10] : _GEN_4619; // @[Execute.scala 117:10]
  assign _GEN_4621 = 6'hb == _T_444 ? welem[11] : _GEN_4620; // @[Execute.scala 117:10]
  assign _GEN_4622 = 6'hc == _T_444 ? welem[12] : _GEN_4621; // @[Execute.scala 117:10]
  assign _GEN_4623 = 6'hd == _T_444 ? welem[13] : _GEN_4622; // @[Execute.scala 117:10]
  assign _GEN_4624 = 6'he == _T_444 ? welem[14] : _GEN_4623; // @[Execute.scala 117:10]
  assign _GEN_4625 = 6'hf == _T_444 ? welem[15] : _GEN_4624; // @[Execute.scala 117:10]
  assign _GEN_4626 = 6'h10 == _T_444 ? welem[16] : _GEN_4625; // @[Execute.scala 117:10]
  assign _GEN_4627 = 6'h11 == _T_444 ? welem[17] : _GEN_4626; // @[Execute.scala 117:10]
  assign _GEN_4628 = 6'h12 == _T_444 ? welem[18] : _GEN_4627; // @[Execute.scala 117:10]
  assign _GEN_4629 = 6'h13 == _T_444 ? welem[19] : _GEN_4628; // @[Execute.scala 117:10]
  assign _GEN_4630 = 6'h14 == _T_444 ? welem[20] : _GEN_4629; // @[Execute.scala 117:10]
  assign _GEN_4631 = 6'h15 == _T_444 ? welem[21] : _GEN_4630; // @[Execute.scala 117:10]
  assign _GEN_4632 = 6'h16 == _T_444 ? welem[22] : _GEN_4631; // @[Execute.scala 117:10]
  assign _GEN_4633 = 6'h17 == _T_444 ? welem[23] : _GEN_4632; // @[Execute.scala 117:10]
  assign _GEN_4634 = 6'h18 == _T_444 ? welem[24] : _GEN_4633; // @[Execute.scala 117:10]
  assign _GEN_4635 = 6'h19 == _T_444 ? welem[25] : _GEN_4634; // @[Execute.scala 117:10]
  assign _GEN_4636 = 6'h1a == _T_444 ? welem[26] : _GEN_4635; // @[Execute.scala 117:10]
  assign _GEN_4637 = 6'h1b == _T_444 ? welem[27] : _GEN_4636; // @[Execute.scala 117:10]
  assign _GEN_4638 = 6'h1c == _T_444 ? welem[28] : _GEN_4637; // @[Execute.scala 117:10]
  assign _GEN_4639 = 6'h1d == _T_444 ? welem[29] : _GEN_4638; // @[Execute.scala 117:10]
  assign _GEN_4640 = 6'h1e == _T_444 ? welem[30] : _GEN_4639; // @[Execute.scala 117:10]
  assign _GEN_4641 = 6'h1f == _T_444 ? welem[31] : _GEN_4640; // @[Execute.scala 117:10]
  assign _GEN_4642 = 6'h20 == _T_444 ? welem[32] : _GEN_4641; // @[Execute.scala 117:10]
  assign _GEN_4643 = 6'h21 == _T_444 ? welem[33] : _GEN_4642; // @[Execute.scala 117:10]
  assign _GEN_4644 = 6'h22 == _T_444 ? welem[34] : _GEN_4643; // @[Execute.scala 117:10]
  assign _GEN_4645 = 6'h23 == _T_444 ? welem[35] : _GEN_4644; // @[Execute.scala 117:10]
  assign _GEN_4646 = 6'h24 == _T_444 ? welem[36] : _GEN_4645; // @[Execute.scala 117:10]
  assign _GEN_4647 = 6'h25 == _T_444 ? welem[37] : _GEN_4646; // @[Execute.scala 117:10]
  assign _GEN_4648 = 6'h26 == _T_444 ? welem[38] : _GEN_4647; // @[Execute.scala 117:10]
  assign _GEN_4649 = 6'h27 == _T_444 ? welem[39] : _GEN_4648; // @[Execute.scala 117:10]
  assign _GEN_4650 = 6'h28 == _T_444 ? welem[40] : _GEN_4649; // @[Execute.scala 117:10]
  assign _GEN_4651 = 6'h29 == _T_444 ? welem[41] : _GEN_4650; // @[Execute.scala 117:10]
  assign _GEN_4652 = 6'h2a == _T_444 ? welem[42] : _GEN_4651; // @[Execute.scala 117:10]
  assign _GEN_4653 = 6'h2b == _T_444 ? welem[43] : _GEN_4652; // @[Execute.scala 117:10]
  assign _GEN_4654 = 6'h2c == _T_444 ? welem[44] : _GEN_4653; // @[Execute.scala 117:10]
  assign _GEN_4655 = 6'h2d == _T_444 ? welem[45] : _GEN_4654; // @[Execute.scala 117:10]
  assign _GEN_4656 = 6'h2e == _T_444 ? welem[46] : _GEN_4655; // @[Execute.scala 117:10]
  assign _GEN_4657 = 6'h2f == _T_444 ? welem[47] : _GEN_4656; // @[Execute.scala 117:10]
  assign _GEN_4658 = 6'h30 == _T_444 ? welem[48] : _GEN_4657; // @[Execute.scala 117:10]
  assign _GEN_4659 = 6'h31 == _T_444 ? welem[49] : _GEN_4658; // @[Execute.scala 117:10]
  assign _GEN_4660 = 6'h32 == _T_444 ? welem[50] : _GEN_4659; // @[Execute.scala 117:10]
  assign _GEN_4661 = 6'h33 == _T_444 ? welem[51] : _GEN_4660; // @[Execute.scala 117:10]
  assign _GEN_4662 = 6'h34 == _T_444 ? welem[52] : _GEN_4661; // @[Execute.scala 117:10]
  assign _GEN_4663 = 6'h35 == _T_444 ? welem[53] : _GEN_4662; // @[Execute.scala 117:10]
  assign _GEN_4664 = 6'h36 == _T_444 ? welem[54] : _GEN_4663; // @[Execute.scala 117:10]
  assign _GEN_4665 = 6'h37 == _T_444 ? welem[55] : _GEN_4664; // @[Execute.scala 117:10]
  assign _GEN_4666 = 6'h38 == _T_444 ? welem[56] : _GEN_4665; // @[Execute.scala 117:10]
  assign _GEN_4667 = 6'h39 == _T_444 ? welem[57] : _GEN_4666; // @[Execute.scala 117:10]
  assign _GEN_4668 = 6'h3a == _T_444 ? welem[58] : _GEN_4667; // @[Execute.scala 117:10]
  assign _GEN_4669 = 6'h3b == _T_444 ? welem[59] : _GEN_4668; // @[Execute.scala 117:10]
  assign _GEN_4670 = 6'h3c == _T_444 ? welem[60] : _GEN_4669; // @[Execute.scala 117:10]
  assign _GEN_4671 = 6'h3d == _T_444 ? welem[61] : _GEN_4670; // @[Execute.scala 117:10]
  assign _GEN_4672 = 6'h3e == _T_444 ? welem[62] : _GEN_4671; // @[Execute.scala 117:10]
  assign _GEN_4673 = 6'h3f == _T_444 ? welem[63] : _GEN_4672; // @[Execute.scala 117:10]
  assign _GEN_4675 = 6'h1 == _T_448 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4676 = 6'h2 == _T_448 ? welem[2] : _GEN_4675; // @[Execute.scala 117:10]
  assign _GEN_4677 = 6'h3 == _T_448 ? welem[3] : _GEN_4676; // @[Execute.scala 117:10]
  assign _GEN_4678 = 6'h4 == _T_448 ? welem[4] : _GEN_4677; // @[Execute.scala 117:10]
  assign _GEN_4679 = 6'h5 == _T_448 ? welem[5] : _GEN_4678; // @[Execute.scala 117:10]
  assign _GEN_4680 = 6'h6 == _T_448 ? welem[6] : _GEN_4679; // @[Execute.scala 117:10]
  assign _GEN_4681 = 6'h7 == _T_448 ? welem[7] : _GEN_4680; // @[Execute.scala 117:10]
  assign _GEN_4682 = 6'h8 == _T_448 ? welem[8] : _GEN_4681; // @[Execute.scala 117:10]
  assign _GEN_4683 = 6'h9 == _T_448 ? welem[9] : _GEN_4682; // @[Execute.scala 117:10]
  assign _GEN_4684 = 6'ha == _T_448 ? welem[10] : _GEN_4683; // @[Execute.scala 117:10]
  assign _GEN_4685 = 6'hb == _T_448 ? welem[11] : _GEN_4684; // @[Execute.scala 117:10]
  assign _GEN_4686 = 6'hc == _T_448 ? welem[12] : _GEN_4685; // @[Execute.scala 117:10]
  assign _GEN_4687 = 6'hd == _T_448 ? welem[13] : _GEN_4686; // @[Execute.scala 117:10]
  assign _GEN_4688 = 6'he == _T_448 ? welem[14] : _GEN_4687; // @[Execute.scala 117:10]
  assign _GEN_4689 = 6'hf == _T_448 ? welem[15] : _GEN_4688; // @[Execute.scala 117:10]
  assign _GEN_4690 = 6'h10 == _T_448 ? welem[16] : _GEN_4689; // @[Execute.scala 117:10]
  assign _GEN_4691 = 6'h11 == _T_448 ? welem[17] : _GEN_4690; // @[Execute.scala 117:10]
  assign _GEN_4692 = 6'h12 == _T_448 ? welem[18] : _GEN_4691; // @[Execute.scala 117:10]
  assign _GEN_4693 = 6'h13 == _T_448 ? welem[19] : _GEN_4692; // @[Execute.scala 117:10]
  assign _GEN_4694 = 6'h14 == _T_448 ? welem[20] : _GEN_4693; // @[Execute.scala 117:10]
  assign _GEN_4695 = 6'h15 == _T_448 ? welem[21] : _GEN_4694; // @[Execute.scala 117:10]
  assign _GEN_4696 = 6'h16 == _T_448 ? welem[22] : _GEN_4695; // @[Execute.scala 117:10]
  assign _GEN_4697 = 6'h17 == _T_448 ? welem[23] : _GEN_4696; // @[Execute.scala 117:10]
  assign _GEN_4698 = 6'h18 == _T_448 ? welem[24] : _GEN_4697; // @[Execute.scala 117:10]
  assign _GEN_4699 = 6'h19 == _T_448 ? welem[25] : _GEN_4698; // @[Execute.scala 117:10]
  assign _GEN_4700 = 6'h1a == _T_448 ? welem[26] : _GEN_4699; // @[Execute.scala 117:10]
  assign _GEN_4701 = 6'h1b == _T_448 ? welem[27] : _GEN_4700; // @[Execute.scala 117:10]
  assign _GEN_4702 = 6'h1c == _T_448 ? welem[28] : _GEN_4701; // @[Execute.scala 117:10]
  assign _GEN_4703 = 6'h1d == _T_448 ? welem[29] : _GEN_4702; // @[Execute.scala 117:10]
  assign _GEN_4704 = 6'h1e == _T_448 ? welem[30] : _GEN_4703; // @[Execute.scala 117:10]
  assign _GEN_4705 = 6'h1f == _T_448 ? welem[31] : _GEN_4704; // @[Execute.scala 117:10]
  assign _GEN_4706 = 6'h20 == _T_448 ? welem[32] : _GEN_4705; // @[Execute.scala 117:10]
  assign _GEN_4707 = 6'h21 == _T_448 ? welem[33] : _GEN_4706; // @[Execute.scala 117:10]
  assign _GEN_4708 = 6'h22 == _T_448 ? welem[34] : _GEN_4707; // @[Execute.scala 117:10]
  assign _GEN_4709 = 6'h23 == _T_448 ? welem[35] : _GEN_4708; // @[Execute.scala 117:10]
  assign _GEN_4710 = 6'h24 == _T_448 ? welem[36] : _GEN_4709; // @[Execute.scala 117:10]
  assign _GEN_4711 = 6'h25 == _T_448 ? welem[37] : _GEN_4710; // @[Execute.scala 117:10]
  assign _GEN_4712 = 6'h26 == _T_448 ? welem[38] : _GEN_4711; // @[Execute.scala 117:10]
  assign _GEN_4713 = 6'h27 == _T_448 ? welem[39] : _GEN_4712; // @[Execute.scala 117:10]
  assign _GEN_4714 = 6'h28 == _T_448 ? welem[40] : _GEN_4713; // @[Execute.scala 117:10]
  assign _GEN_4715 = 6'h29 == _T_448 ? welem[41] : _GEN_4714; // @[Execute.scala 117:10]
  assign _GEN_4716 = 6'h2a == _T_448 ? welem[42] : _GEN_4715; // @[Execute.scala 117:10]
  assign _GEN_4717 = 6'h2b == _T_448 ? welem[43] : _GEN_4716; // @[Execute.scala 117:10]
  assign _GEN_4718 = 6'h2c == _T_448 ? welem[44] : _GEN_4717; // @[Execute.scala 117:10]
  assign _GEN_4719 = 6'h2d == _T_448 ? welem[45] : _GEN_4718; // @[Execute.scala 117:10]
  assign _GEN_4720 = 6'h2e == _T_448 ? welem[46] : _GEN_4719; // @[Execute.scala 117:10]
  assign _GEN_4721 = 6'h2f == _T_448 ? welem[47] : _GEN_4720; // @[Execute.scala 117:10]
  assign _GEN_4722 = 6'h30 == _T_448 ? welem[48] : _GEN_4721; // @[Execute.scala 117:10]
  assign _GEN_4723 = 6'h31 == _T_448 ? welem[49] : _GEN_4722; // @[Execute.scala 117:10]
  assign _GEN_4724 = 6'h32 == _T_448 ? welem[50] : _GEN_4723; // @[Execute.scala 117:10]
  assign _GEN_4725 = 6'h33 == _T_448 ? welem[51] : _GEN_4724; // @[Execute.scala 117:10]
  assign _GEN_4726 = 6'h34 == _T_448 ? welem[52] : _GEN_4725; // @[Execute.scala 117:10]
  assign _GEN_4727 = 6'h35 == _T_448 ? welem[53] : _GEN_4726; // @[Execute.scala 117:10]
  assign _GEN_4728 = 6'h36 == _T_448 ? welem[54] : _GEN_4727; // @[Execute.scala 117:10]
  assign _GEN_4729 = 6'h37 == _T_448 ? welem[55] : _GEN_4728; // @[Execute.scala 117:10]
  assign _GEN_4730 = 6'h38 == _T_448 ? welem[56] : _GEN_4729; // @[Execute.scala 117:10]
  assign _GEN_4731 = 6'h39 == _T_448 ? welem[57] : _GEN_4730; // @[Execute.scala 117:10]
  assign _GEN_4732 = 6'h3a == _T_448 ? welem[58] : _GEN_4731; // @[Execute.scala 117:10]
  assign _GEN_4733 = 6'h3b == _T_448 ? welem[59] : _GEN_4732; // @[Execute.scala 117:10]
  assign _GEN_4734 = 6'h3c == _T_448 ? welem[60] : _GEN_4733; // @[Execute.scala 117:10]
  assign _GEN_4735 = 6'h3d == _T_448 ? welem[61] : _GEN_4734; // @[Execute.scala 117:10]
  assign _GEN_4736 = 6'h3e == _T_448 ? welem[62] : _GEN_4735; // @[Execute.scala 117:10]
  assign _GEN_4737 = 6'h3f == _T_448 ? welem[63] : _GEN_4736; // @[Execute.scala 117:10]
  assign _T_451 = _T_442 ? _GEN_4673 : _GEN_4737; // @[Execute.scala 117:10]
  assign _T_452 = r < 6'h1c; // @[Execute.scala 117:15]
  assign _T_454 = r - 6'h1c; // @[Execute.scala 117:37]
  assign _T_458 = 6'h24 + r; // @[Execute.scala 117:60]
  assign _GEN_4739 = 6'h1 == _T_454 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4740 = 6'h2 == _T_454 ? welem[2] : _GEN_4739; // @[Execute.scala 117:10]
  assign _GEN_4741 = 6'h3 == _T_454 ? welem[3] : _GEN_4740; // @[Execute.scala 117:10]
  assign _GEN_4742 = 6'h4 == _T_454 ? welem[4] : _GEN_4741; // @[Execute.scala 117:10]
  assign _GEN_4743 = 6'h5 == _T_454 ? welem[5] : _GEN_4742; // @[Execute.scala 117:10]
  assign _GEN_4744 = 6'h6 == _T_454 ? welem[6] : _GEN_4743; // @[Execute.scala 117:10]
  assign _GEN_4745 = 6'h7 == _T_454 ? welem[7] : _GEN_4744; // @[Execute.scala 117:10]
  assign _GEN_4746 = 6'h8 == _T_454 ? welem[8] : _GEN_4745; // @[Execute.scala 117:10]
  assign _GEN_4747 = 6'h9 == _T_454 ? welem[9] : _GEN_4746; // @[Execute.scala 117:10]
  assign _GEN_4748 = 6'ha == _T_454 ? welem[10] : _GEN_4747; // @[Execute.scala 117:10]
  assign _GEN_4749 = 6'hb == _T_454 ? welem[11] : _GEN_4748; // @[Execute.scala 117:10]
  assign _GEN_4750 = 6'hc == _T_454 ? welem[12] : _GEN_4749; // @[Execute.scala 117:10]
  assign _GEN_4751 = 6'hd == _T_454 ? welem[13] : _GEN_4750; // @[Execute.scala 117:10]
  assign _GEN_4752 = 6'he == _T_454 ? welem[14] : _GEN_4751; // @[Execute.scala 117:10]
  assign _GEN_4753 = 6'hf == _T_454 ? welem[15] : _GEN_4752; // @[Execute.scala 117:10]
  assign _GEN_4754 = 6'h10 == _T_454 ? welem[16] : _GEN_4753; // @[Execute.scala 117:10]
  assign _GEN_4755 = 6'h11 == _T_454 ? welem[17] : _GEN_4754; // @[Execute.scala 117:10]
  assign _GEN_4756 = 6'h12 == _T_454 ? welem[18] : _GEN_4755; // @[Execute.scala 117:10]
  assign _GEN_4757 = 6'h13 == _T_454 ? welem[19] : _GEN_4756; // @[Execute.scala 117:10]
  assign _GEN_4758 = 6'h14 == _T_454 ? welem[20] : _GEN_4757; // @[Execute.scala 117:10]
  assign _GEN_4759 = 6'h15 == _T_454 ? welem[21] : _GEN_4758; // @[Execute.scala 117:10]
  assign _GEN_4760 = 6'h16 == _T_454 ? welem[22] : _GEN_4759; // @[Execute.scala 117:10]
  assign _GEN_4761 = 6'h17 == _T_454 ? welem[23] : _GEN_4760; // @[Execute.scala 117:10]
  assign _GEN_4762 = 6'h18 == _T_454 ? welem[24] : _GEN_4761; // @[Execute.scala 117:10]
  assign _GEN_4763 = 6'h19 == _T_454 ? welem[25] : _GEN_4762; // @[Execute.scala 117:10]
  assign _GEN_4764 = 6'h1a == _T_454 ? welem[26] : _GEN_4763; // @[Execute.scala 117:10]
  assign _GEN_4765 = 6'h1b == _T_454 ? welem[27] : _GEN_4764; // @[Execute.scala 117:10]
  assign _GEN_4766 = 6'h1c == _T_454 ? welem[28] : _GEN_4765; // @[Execute.scala 117:10]
  assign _GEN_4767 = 6'h1d == _T_454 ? welem[29] : _GEN_4766; // @[Execute.scala 117:10]
  assign _GEN_4768 = 6'h1e == _T_454 ? welem[30] : _GEN_4767; // @[Execute.scala 117:10]
  assign _GEN_4769 = 6'h1f == _T_454 ? welem[31] : _GEN_4768; // @[Execute.scala 117:10]
  assign _GEN_4770 = 6'h20 == _T_454 ? welem[32] : _GEN_4769; // @[Execute.scala 117:10]
  assign _GEN_4771 = 6'h21 == _T_454 ? welem[33] : _GEN_4770; // @[Execute.scala 117:10]
  assign _GEN_4772 = 6'h22 == _T_454 ? welem[34] : _GEN_4771; // @[Execute.scala 117:10]
  assign _GEN_4773 = 6'h23 == _T_454 ? welem[35] : _GEN_4772; // @[Execute.scala 117:10]
  assign _GEN_4774 = 6'h24 == _T_454 ? welem[36] : _GEN_4773; // @[Execute.scala 117:10]
  assign _GEN_4775 = 6'h25 == _T_454 ? welem[37] : _GEN_4774; // @[Execute.scala 117:10]
  assign _GEN_4776 = 6'h26 == _T_454 ? welem[38] : _GEN_4775; // @[Execute.scala 117:10]
  assign _GEN_4777 = 6'h27 == _T_454 ? welem[39] : _GEN_4776; // @[Execute.scala 117:10]
  assign _GEN_4778 = 6'h28 == _T_454 ? welem[40] : _GEN_4777; // @[Execute.scala 117:10]
  assign _GEN_4779 = 6'h29 == _T_454 ? welem[41] : _GEN_4778; // @[Execute.scala 117:10]
  assign _GEN_4780 = 6'h2a == _T_454 ? welem[42] : _GEN_4779; // @[Execute.scala 117:10]
  assign _GEN_4781 = 6'h2b == _T_454 ? welem[43] : _GEN_4780; // @[Execute.scala 117:10]
  assign _GEN_4782 = 6'h2c == _T_454 ? welem[44] : _GEN_4781; // @[Execute.scala 117:10]
  assign _GEN_4783 = 6'h2d == _T_454 ? welem[45] : _GEN_4782; // @[Execute.scala 117:10]
  assign _GEN_4784 = 6'h2e == _T_454 ? welem[46] : _GEN_4783; // @[Execute.scala 117:10]
  assign _GEN_4785 = 6'h2f == _T_454 ? welem[47] : _GEN_4784; // @[Execute.scala 117:10]
  assign _GEN_4786 = 6'h30 == _T_454 ? welem[48] : _GEN_4785; // @[Execute.scala 117:10]
  assign _GEN_4787 = 6'h31 == _T_454 ? welem[49] : _GEN_4786; // @[Execute.scala 117:10]
  assign _GEN_4788 = 6'h32 == _T_454 ? welem[50] : _GEN_4787; // @[Execute.scala 117:10]
  assign _GEN_4789 = 6'h33 == _T_454 ? welem[51] : _GEN_4788; // @[Execute.scala 117:10]
  assign _GEN_4790 = 6'h34 == _T_454 ? welem[52] : _GEN_4789; // @[Execute.scala 117:10]
  assign _GEN_4791 = 6'h35 == _T_454 ? welem[53] : _GEN_4790; // @[Execute.scala 117:10]
  assign _GEN_4792 = 6'h36 == _T_454 ? welem[54] : _GEN_4791; // @[Execute.scala 117:10]
  assign _GEN_4793 = 6'h37 == _T_454 ? welem[55] : _GEN_4792; // @[Execute.scala 117:10]
  assign _GEN_4794 = 6'h38 == _T_454 ? welem[56] : _GEN_4793; // @[Execute.scala 117:10]
  assign _GEN_4795 = 6'h39 == _T_454 ? welem[57] : _GEN_4794; // @[Execute.scala 117:10]
  assign _GEN_4796 = 6'h3a == _T_454 ? welem[58] : _GEN_4795; // @[Execute.scala 117:10]
  assign _GEN_4797 = 6'h3b == _T_454 ? welem[59] : _GEN_4796; // @[Execute.scala 117:10]
  assign _GEN_4798 = 6'h3c == _T_454 ? welem[60] : _GEN_4797; // @[Execute.scala 117:10]
  assign _GEN_4799 = 6'h3d == _T_454 ? welem[61] : _GEN_4798; // @[Execute.scala 117:10]
  assign _GEN_4800 = 6'h3e == _T_454 ? welem[62] : _GEN_4799; // @[Execute.scala 117:10]
  assign _GEN_4801 = 6'h3f == _T_454 ? welem[63] : _GEN_4800; // @[Execute.scala 117:10]
  assign _GEN_4803 = 6'h1 == _T_458 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4804 = 6'h2 == _T_458 ? welem[2] : _GEN_4803; // @[Execute.scala 117:10]
  assign _GEN_4805 = 6'h3 == _T_458 ? welem[3] : _GEN_4804; // @[Execute.scala 117:10]
  assign _GEN_4806 = 6'h4 == _T_458 ? welem[4] : _GEN_4805; // @[Execute.scala 117:10]
  assign _GEN_4807 = 6'h5 == _T_458 ? welem[5] : _GEN_4806; // @[Execute.scala 117:10]
  assign _GEN_4808 = 6'h6 == _T_458 ? welem[6] : _GEN_4807; // @[Execute.scala 117:10]
  assign _GEN_4809 = 6'h7 == _T_458 ? welem[7] : _GEN_4808; // @[Execute.scala 117:10]
  assign _GEN_4810 = 6'h8 == _T_458 ? welem[8] : _GEN_4809; // @[Execute.scala 117:10]
  assign _GEN_4811 = 6'h9 == _T_458 ? welem[9] : _GEN_4810; // @[Execute.scala 117:10]
  assign _GEN_4812 = 6'ha == _T_458 ? welem[10] : _GEN_4811; // @[Execute.scala 117:10]
  assign _GEN_4813 = 6'hb == _T_458 ? welem[11] : _GEN_4812; // @[Execute.scala 117:10]
  assign _GEN_4814 = 6'hc == _T_458 ? welem[12] : _GEN_4813; // @[Execute.scala 117:10]
  assign _GEN_4815 = 6'hd == _T_458 ? welem[13] : _GEN_4814; // @[Execute.scala 117:10]
  assign _GEN_4816 = 6'he == _T_458 ? welem[14] : _GEN_4815; // @[Execute.scala 117:10]
  assign _GEN_4817 = 6'hf == _T_458 ? welem[15] : _GEN_4816; // @[Execute.scala 117:10]
  assign _GEN_4818 = 6'h10 == _T_458 ? welem[16] : _GEN_4817; // @[Execute.scala 117:10]
  assign _GEN_4819 = 6'h11 == _T_458 ? welem[17] : _GEN_4818; // @[Execute.scala 117:10]
  assign _GEN_4820 = 6'h12 == _T_458 ? welem[18] : _GEN_4819; // @[Execute.scala 117:10]
  assign _GEN_4821 = 6'h13 == _T_458 ? welem[19] : _GEN_4820; // @[Execute.scala 117:10]
  assign _GEN_4822 = 6'h14 == _T_458 ? welem[20] : _GEN_4821; // @[Execute.scala 117:10]
  assign _GEN_4823 = 6'h15 == _T_458 ? welem[21] : _GEN_4822; // @[Execute.scala 117:10]
  assign _GEN_4824 = 6'h16 == _T_458 ? welem[22] : _GEN_4823; // @[Execute.scala 117:10]
  assign _GEN_4825 = 6'h17 == _T_458 ? welem[23] : _GEN_4824; // @[Execute.scala 117:10]
  assign _GEN_4826 = 6'h18 == _T_458 ? welem[24] : _GEN_4825; // @[Execute.scala 117:10]
  assign _GEN_4827 = 6'h19 == _T_458 ? welem[25] : _GEN_4826; // @[Execute.scala 117:10]
  assign _GEN_4828 = 6'h1a == _T_458 ? welem[26] : _GEN_4827; // @[Execute.scala 117:10]
  assign _GEN_4829 = 6'h1b == _T_458 ? welem[27] : _GEN_4828; // @[Execute.scala 117:10]
  assign _GEN_4830 = 6'h1c == _T_458 ? welem[28] : _GEN_4829; // @[Execute.scala 117:10]
  assign _GEN_4831 = 6'h1d == _T_458 ? welem[29] : _GEN_4830; // @[Execute.scala 117:10]
  assign _GEN_4832 = 6'h1e == _T_458 ? welem[30] : _GEN_4831; // @[Execute.scala 117:10]
  assign _GEN_4833 = 6'h1f == _T_458 ? welem[31] : _GEN_4832; // @[Execute.scala 117:10]
  assign _GEN_4834 = 6'h20 == _T_458 ? welem[32] : _GEN_4833; // @[Execute.scala 117:10]
  assign _GEN_4835 = 6'h21 == _T_458 ? welem[33] : _GEN_4834; // @[Execute.scala 117:10]
  assign _GEN_4836 = 6'h22 == _T_458 ? welem[34] : _GEN_4835; // @[Execute.scala 117:10]
  assign _GEN_4837 = 6'h23 == _T_458 ? welem[35] : _GEN_4836; // @[Execute.scala 117:10]
  assign _GEN_4838 = 6'h24 == _T_458 ? welem[36] : _GEN_4837; // @[Execute.scala 117:10]
  assign _GEN_4839 = 6'h25 == _T_458 ? welem[37] : _GEN_4838; // @[Execute.scala 117:10]
  assign _GEN_4840 = 6'h26 == _T_458 ? welem[38] : _GEN_4839; // @[Execute.scala 117:10]
  assign _GEN_4841 = 6'h27 == _T_458 ? welem[39] : _GEN_4840; // @[Execute.scala 117:10]
  assign _GEN_4842 = 6'h28 == _T_458 ? welem[40] : _GEN_4841; // @[Execute.scala 117:10]
  assign _GEN_4843 = 6'h29 == _T_458 ? welem[41] : _GEN_4842; // @[Execute.scala 117:10]
  assign _GEN_4844 = 6'h2a == _T_458 ? welem[42] : _GEN_4843; // @[Execute.scala 117:10]
  assign _GEN_4845 = 6'h2b == _T_458 ? welem[43] : _GEN_4844; // @[Execute.scala 117:10]
  assign _GEN_4846 = 6'h2c == _T_458 ? welem[44] : _GEN_4845; // @[Execute.scala 117:10]
  assign _GEN_4847 = 6'h2d == _T_458 ? welem[45] : _GEN_4846; // @[Execute.scala 117:10]
  assign _GEN_4848 = 6'h2e == _T_458 ? welem[46] : _GEN_4847; // @[Execute.scala 117:10]
  assign _GEN_4849 = 6'h2f == _T_458 ? welem[47] : _GEN_4848; // @[Execute.scala 117:10]
  assign _GEN_4850 = 6'h30 == _T_458 ? welem[48] : _GEN_4849; // @[Execute.scala 117:10]
  assign _GEN_4851 = 6'h31 == _T_458 ? welem[49] : _GEN_4850; // @[Execute.scala 117:10]
  assign _GEN_4852 = 6'h32 == _T_458 ? welem[50] : _GEN_4851; // @[Execute.scala 117:10]
  assign _GEN_4853 = 6'h33 == _T_458 ? welem[51] : _GEN_4852; // @[Execute.scala 117:10]
  assign _GEN_4854 = 6'h34 == _T_458 ? welem[52] : _GEN_4853; // @[Execute.scala 117:10]
  assign _GEN_4855 = 6'h35 == _T_458 ? welem[53] : _GEN_4854; // @[Execute.scala 117:10]
  assign _GEN_4856 = 6'h36 == _T_458 ? welem[54] : _GEN_4855; // @[Execute.scala 117:10]
  assign _GEN_4857 = 6'h37 == _T_458 ? welem[55] : _GEN_4856; // @[Execute.scala 117:10]
  assign _GEN_4858 = 6'h38 == _T_458 ? welem[56] : _GEN_4857; // @[Execute.scala 117:10]
  assign _GEN_4859 = 6'h39 == _T_458 ? welem[57] : _GEN_4858; // @[Execute.scala 117:10]
  assign _GEN_4860 = 6'h3a == _T_458 ? welem[58] : _GEN_4859; // @[Execute.scala 117:10]
  assign _GEN_4861 = 6'h3b == _T_458 ? welem[59] : _GEN_4860; // @[Execute.scala 117:10]
  assign _GEN_4862 = 6'h3c == _T_458 ? welem[60] : _GEN_4861; // @[Execute.scala 117:10]
  assign _GEN_4863 = 6'h3d == _T_458 ? welem[61] : _GEN_4862; // @[Execute.scala 117:10]
  assign _GEN_4864 = 6'h3e == _T_458 ? welem[62] : _GEN_4863; // @[Execute.scala 117:10]
  assign _GEN_4865 = 6'h3f == _T_458 ? welem[63] : _GEN_4864; // @[Execute.scala 117:10]
  assign _T_461 = _T_452 ? _GEN_4801 : _GEN_4865; // @[Execute.scala 117:10]
  assign _T_462 = r < 6'h1b; // @[Execute.scala 117:15]
  assign _T_464 = r - 6'h1b; // @[Execute.scala 117:37]
  assign _T_468 = 6'h25 + r; // @[Execute.scala 117:60]
  assign _GEN_4867 = 6'h1 == _T_464 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4868 = 6'h2 == _T_464 ? welem[2] : _GEN_4867; // @[Execute.scala 117:10]
  assign _GEN_4869 = 6'h3 == _T_464 ? welem[3] : _GEN_4868; // @[Execute.scala 117:10]
  assign _GEN_4870 = 6'h4 == _T_464 ? welem[4] : _GEN_4869; // @[Execute.scala 117:10]
  assign _GEN_4871 = 6'h5 == _T_464 ? welem[5] : _GEN_4870; // @[Execute.scala 117:10]
  assign _GEN_4872 = 6'h6 == _T_464 ? welem[6] : _GEN_4871; // @[Execute.scala 117:10]
  assign _GEN_4873 = 6'h7 == _T_464 ? welem[7] : _GEN_4872; // @[Execute.scala 117:10]
  assign _GEN_4874 = 6'h8 == _T_464 ? welem[8] : _GEN_4873; // @[Execute.scala 117:10]
  assign _GEN_4875 = 6'h9 == _T_464 ? welem[9] : _GEN_4874; // @[Execute.scala 117:10]
  assign _GEN_4876 = 6'ha == _T_464 ? welem[10] : _GEN_4875; // @[Execute.scala 117:10]
  assign _GEN_4877 = 6'hb == _T_464 ? welem[11] : _GEN_4876; // @[Execute.scala 117:10]
  assign _GEN_4878 = 6'hc == _T_464 ? welem[12] : _GEN_4877; // @[Execute.scala 117:10]
  assign _GEN_4879 = 6'hd == _T_464 ? welem[13] : _GEN_4878; // @[Execute.scala 117:10]
  assign _GEN_4880 = 6'he == _T_464 ? welem[14] : _GEN_4879; // @[Execute.scala 117:10]
  assign _GEN_4881 = 6'hf == _T_464 ? welem[15] : _GEN_4880; // @[Execute.scala 117:10]
  assign _GEN_4882 = 6'h10 == _T_464 ? welem[16] : _GEN_4881; // @[Execute.scala 117:10]
  assign _GEN_4883 = 6'h11 == _T_464 ? welem[17] : _GEN_4882; // @[Execute.scala 117:10]
  assign _GEN_4884 = 6'h12 == _T_464 ? welem[18] : _GEN_4883; // @[Execute.scala 117:10]
  assign _GEN_4885 = 6'h13 == _T_464 ? welem[19] : _GEN_4884; // @[Execute.scala 117:10]
  assign _GEN_4886 = 6'h14 == _T_464 ? welem[20] : _GEN_4885; // @[Execute.scala 117:10]
  assign _GEN_4887 = 6'h15 == _T_464 ? welem[21] : _GEN_4886; // @[Execute.scala 117:10]
  assign _GEN_4888 = 6'h16 == _T_464 ? welem[22] : _GEN_4887; // @[Execute.scala 117:10]
  assign _GEN_4889 = 6'h17 == _T_464 ? welem[23] : _GEN_4888; // @[Execute.scala 117:10]
  assign _GEN_4890 = 6'h18 == _T_464 ? welem[24] : _GEN_4889; // @[Execute.scala 117:10]
  assign _GEN_4891 = 6'h19 == _T_464 ? welem[25] : _GEN_4890; // @[Execute.scala 117:10]
  assign _GEN_4892 = 6'h1a == _T_464 ? welem[26] : _GEN_4891; // @[Execute.scala 117:10]
  assign _GEN_4893 = 6'h1b == _T_464 ? welem[27] : _GEN_4892; // @[Execute.scala 117:10]
  assign _GEN_4894 = 6'h1c == _T_464 ? welem[28] : _GEN_4893; // @[Execute.scala 117:10]
  assign _GEN_4895 = 6'h1d == _T_464 ? welem[29] : _GEN_4894; // @[Execute.scala 117:10]
  assign _GEN_4896 = 6'h1e == _T_464 ? welem[30] : _GEN_4895; // @[Execute.scala 117:10]
  assign _GEN_4897 = 6'h1f == _T_464 ? welem[31] : _GEN_4896; // @[Execute.scala 117:10]
  assign _GEN_4898 = 6'h20 == _T_464 ? welem[32] : _GEN_4897; // @[Execute.scala 117:10]
  assign _GEN_4899 = 6'h21 == _T_464 ? welem[33] : _GEN_4898; // @[Execute.scala 117:10]
  assign _GEN_4900 = 6'h22 == _T_464 ? welem[34] : _GEN_4899; // @[Execute.scala 117:10]
  assign _GEN_4901 = 6'h23 == _T_464 ? welem[35] : _GEN_4900; // @[Execute.scala 117:10]
  assign _GEN_4902 = 6'h24 == _T_464 ? welem[36] : _GEN_4901; // @[Execute.scala 117:10]
  assign _GEN_4903 = 6'h25 == _T_464 ? welem[37] : _GEN_4902; // @[Execute.scala 117:10]
  assign _GEN_4904 = 6'h26 == _T_464 ? welem[38] : _GEN_4903; // @[Execute.scala 117:10]
  assign _GEN_4905 = 6'h27 == _T_464 ? welem[39] : _GEN_4904; // @[Execute.scala 117:10]
  assign _GEN_4906 = 6'h28 == _T_464 ? welem[40] : _GEN_4905; // @[Execute.scala 117:10]
  assign _GEN_4907 = 6'h29 == _T_464 ? welem[41] : _GEN_4906; // @[Execute.scala 117:10]
  assign _GEN_4908 = 6'h2a == _T_464 ? welem[42] : _GEN_4907; // @[Execute.scala 117:10]
  assign _GEN_4909 = 6'h2b == _T_464 ? welem[43] : _GEN_4908; // @[Execute.scala 117:10]
  assign _GEN_4910 = 6'h2c == _T_464 ? welem[44] : _GEN_4909; // @[Execute.scala 117:10]
  assign _GEN_4911 = 6'h2d == _T_464 ? welem[45] : _GEN_4910; // @[Execute.scala 117:10]
  assign _GEN_4912 = 6'h2e == _T_464 ? welem[46] : _GEN_4911; // @[Execute.scala 117:10]
  assign _GEN_4913 = 6'h2f == _T_464 ? welem[47] : _GEN_4912; // @[Execute.scala 117:10]
  assign _GEN_4914 = 6'h30 == _T_464 ? welem[48] : _GEN_4913; // @[Execute.scala 117:10]
  assign _GEN_4915 = 6'h31 == _T_464 ? welem[49] : _GEN_4914; // @[Execute.scala 117:10]
  assign _GEN_4916 = 6'h32 == _T_464 ? welem[50] : _GEN_4915; // @[Execute.scala 117:10]
  assign _GEN_4917 = 6'h33 == _T_464 ? welem[51] : _GEN_4916; // @[Execute.scala 117:10]
  assign _GEN_4918 = 6'h34 == _T_464 ? welem[52] : _GEN_4917; // @[Execute.scala 117:10]
  assign _GEN_4919 = 6'h35 == _T_464 ? welem[53] : _GEN_4918; // @[Execute.scala 117:10]
  assign _GEN_4920 = 6'h36 == _T_464 ? welem[54] : _GEN_4919; // @[Execute.scala 117:10]
  assign _GEN_4921 = 6'h37 == _T_464 ? welem[55] : _GEN_4920; // @[Execute.scala 117:10]
  assign _GEN_4922 = 6'h38 == _T_464 ? welem[56] : _GEN_4921; // @[Execute.scala 117:10]
  assign _GEN_4923 = 6'h39 == _T_464 ? welem[57] : _GEN_4922; // @[Execute.scala 117:10]
  assign _GEN_4924 = 6'h3a == _T_464 ? welem[58] : _GEN_4923; // @[Execute.scala 117:10]
  assign _GEN_4925 = 6'h3b == _T_464 ? welem[59] : _GEN_4924; // @[Execute.scala 117:10]
  assign _GEN_4926 = 6'h3c == _T_464 ? welem[60] : _GEN_4925; // @[Execute.scala 117:10]
  assign _GEN_4927 = 6'h3d == _T_464 ? welem[61] : _GEN_4926; // @[Execute.scala 117:10]
  assign _GEN_4928 = 6'h3e == _T_464 ? welem[62] : _GEN_4927; // @[Execute.scala 117:10]
  assign _GEN_4929 = 6'h3f == _T_464 ? welem[63] : _GEN_4928; // @[Execute.scala 117:10]
  assign _GEN_4931 = 6'h1 == _T_468 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4932 = 6'h2 == _T_468 ? welem[2] : _GEN_4931; // @[Execute.scala 117:10]
  assign _GEN_4933 = 6'h3 == _T_468 ? welem[3] : _GEN_4932; // @[Execute.scala 117:10]
  assign _GEN_4934 = 6'h4 == _T_468 ? welem[4] : _GEN_4933; // @[Execute.scala 117:10]
  assign _GEN_4935 = 6'h5 == _T_468 ? welem[5] : _GEN_4934; // @[Execute.scala 117:10]
  assign _GEN_4936 = 6'h6 == _T_468 ? welem[6] : _GEN_4935; // @[Execute.scala 117:10]
  assign _GEN_4937 = 6'h7 == _T_468 ? welem[7] : _GEN_4936; // @[Execute.scala 117:10]
  assign _GEN_4938 = 6'h8 == _T_468 ? welem[8] : _GEN_4937; // @[Execute.scala 117:10]
  assign _GEN_4939 = 6'h9 == _T_468 ? welem[9] : _GEN_4938; // @[Execute.scala 117:10]
  assign _GEN_4940 = 6'ha == _T_468 ? welem[10] : _GEN_4939; // @[Execute.scala 117:10]
  assign _GEN_4941 = 6'hb == _T_468 ? welem[11] : _GEN_4940; // @[Execute.scala 117:10]
  assign _GEN_4942 = 6'hc == _T_468 ? welem[12] : _GEN_4941; // @[Execute.scala 117:10]
  assign _GEN_4943 = 6'hd == _T_468 ? welem[13] : _GEN_4942; // @[Execute.scala 117:10]
  assign _GEN_4944 = 6'he == _T_468 ? welem[14] : _GEN_4943; // @[Execute.scala 117:10]
  assign _GEN_4945 = 6'hf == _T_468 ? welem[15] : _GEN_4944; // @[Execute.scala 117:10]
  assign _GEN_4946 = 6'h10 == _T_468 ? welem[16] : _GEN_4945; // @[Execute.scala 117:10]
  assign _GEN_4947 = 6'h11 == _T_468 ? welem[17] : _GEN_4946; // @[Execute.scala 117:10]
  assign _GEN_4948 = 6'h12 == _T_468 ? welem[18] : _GEN_4947; // @[Execute.scala 117:10]
  assign _GEN_4949 = 6'h13 == _T_468 ? welem[19] : _GEN_4948; // @[Execute.scala 117:10]
  assign _GEN_4950 = 6'h14 == _T_468 ? welem[20] : _GEN_4949; // @[Execute.scala 117:10]
  assign _GEN_4951 = 6'h15 == _T_468 ? welem[21] : _GEN_4950; // @[Execute.scala 117:10]
  assign _GEN_4952 = 6'h16 == _T_468 ? welem[22] : _GEN_4951; // @[Execute.scala 117:10]
  assign _GEN_4953 = 6'h17 == _T_468 ? welem[23] : _GEN_4952; // @[Execute.scala 117:10]
  assign _GEN_4954 = 6'h18 == _T_468 ? welem[24] : _GEN_4953; // @[Execute.scala 117:10]
  assign _GEN_4955 = 6'h19 == _T_468 ? welem[25] : _GEN_4954; // @[Execute.scala 117:10]
  assign _GEN_4956 = 6'h1a == _T_468 ? welem[26] : _GEN_4955; // @[Execute.scala 117:10]
  assign _GEN_4957 = 6'h1b == _T_468 ? welem[27] : _GEN_4956; // @[Execute.scala 117:10]
  assign _GEN_4958 = 6'h1c == _T_468 ? welem[28] : _GEN_4957; // @[Execute.scala 117:10]
  assign _GEN_4959 = 6'h1d == _T_468 ? welem[29] : _GEN_4958; // @[Execute.scala 117:10]
  assign _GEN_4960 = 6'h1e == _T_468 ? welem[30] : _GEN_4959; // @[Execute.scala 117:10]
  assign _GEN_4961 = 6'h1f == _T_468 ? welem[31] : _GEN_4960; // @[Execute.scala 117:10]
  assign _GEN_4962 = 6'h20 == _T_468 ? welem[32] : _GEN_4961; // @[Execute.scala 117:10]
  assign _GEN_4963 = 6'h21 == _T_468 ? welem[33] : _GEN_4962; // @[Execute.scala 117:10]
  assign _GEN_4964 = 6'h22 == _T_468 ? welem[34] : _GEN_4963; // @[Execute.scala 117:10]
  assign _GEN_4965 = 6'h23 == _T_468 ? welem[35] : _GEN_4964; // @[Execute.scala 117:10]
  assign _GEN_4966 = 6'h24 == _T_468 ? welem[36] : _GEN_4965; // @[Execute.scala 117:10]
  assign _GEN_4967 = 6'h25 == _T_468 ? welem[37] : _GEN_4966; // @[Execute.scala 117:10]
  assign _GEN_4968 = 6'h26 == _T_468 ? welem[38] : _GEN_4967; // @[Execute.scala 117:10]
  assign _GEN_4969 = 6'h27 == _T_468 ? welem[39] : _GEN_4968; // @[Execute.scala 117:10]
  assign _GEN_4970 = 6'h28 == _T_468 ? welem[40] : _GEN_4969; // @[Execute.scala 117:10]
  assign _GEN_4971 = 6'h29 == _T_468 ? welem[41] : _GEN_4970; // @[Execute.scala 117:10]
  assign _GEN_4972 = 6'h2a == _T_468 ? welem[42] : _GEN_4971; // @[Execute.scala 117:10]
  assign _GEN_4973 = 6'h2b == _T_468 ? welem[43] : _GEN_4972; // @[Execute.scala 117:10]
  assign _GEN_4974 = 6'h2c == _T_468 ? welem[44] : _GEN_4973; // @[Execute.scala 117:10]
  assign _GEN_4975 = 6'h2d == _T_468 ? welem[45] : _GEN_4974; // @[Execute.scala 117:10]
  assign _GEN_4976 = 6'h2e == _T_468 ? welem[46] : _GEN_4975; // @[Execute.scala 117:10]
  assign _GEN_4977 = 6'h2f == _T_468 ? welem[47] : _GEN_4976; // @[Execute.scala 117:10]
  assign _GEN_4978 = 6'h30 == _T_468 ? welem[48] : _GEN_4977; // @[Execute.scala 117:10]
  assign _GEN_4979 = 6'h31 == _T_468 ? welem[49] : _GEN_4978; // @[Execute.scala 117:10]
  assign _GEN_4980 = 6'h32 == _T_468 ? welem[50] : _GEN_4979; // @[Execute.scala 117:10]
  assign _GEN_4981 = 6'h33 == _T_468 ? welem[51] : _GEN_4980; // @[Execute.scala 117:10]
  assign _GEN_4982 = 6'h34 == _T_468 ? welem[52] : _GEN_4981; // @[Execute.scala 117:10]
  assign _GEN_4983 = 6'h35 == _T_468 ? welem[53] : _GEN_4982; // @[Execute.scala 117:10]
  assign _GEN_4984 = 6'h36 == _T_468 ? welem[54] : _GEN_4983; // @[Execute.scala 117:10]
  assign _GEN_4985 = 6'h37 == _T_468 ? welem[55] : _GEN_4984; // @[Execute.scala 117:10]
  assign _GEN_4986 = 6'h38 == _T_468 ? welem[56] : _GEN_4985; // @[Execute.scala 117:10]
  assign _GEN_4987 = 6'h39 == _T_468 ? welem[57] : _GEN_4986; // @[Execute.scala 117:10]
  assign _GEN_4988 = 6'h3a == _T_468 ? welem[58] : _GEN_4987; // @[Execute.scala 117:10]
  assign _GEN_4989 = 6'h3b == _T_468 ? welem[59] : _GEN_4988; // @[Execute.scala 117:10]
  assign _GEN_4990 = 6'h3c == _T_468 ? welem[60] : _GEN_4989; // @[Execute.scala 117:10]
  assign _GEN_4991 = 6'h3d == _T_468 ? welem[61] : _GEN_4990; // @[Execute.scala 117:10]
  assign _GEN_4992 = 6'h3e == _T_468 ? welem[62] : _GEN_4991; // @[Execute.scala 117:10]
  assign _GEN_4993 = 6'h3f == _T_468 ? welem[63] : _GEN_4992; // @[Execute.scala 117:10]
  assign _T_471 = _T_462 ? _GEN_4929 : _GEN_4993; // @[Execute.scala 117:10]
  assign _T_472 = r < 6'h1a; // @[Execute.scala 117:15]
  assign _T_474 = r - 6'h1a; // @[Execute.scala 117:37]
  assign _T_478 = 6'h26 + r; // @[Execute.scala 117:60]
  assign _GEN_4995 = 6'h1 == _T_474 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_4996 = 6'h2 == _T_474 ? welem[2] : _GEN_4995; // @[Execute.scala 117:10]
  assign _GEN_4997 = 6'h3 == _T_474 ? welem[3] : _GEN_4996; // @[Execute.scala 117:10]
  assign _GEN_4998 = 6'h4 == _T_474 ? welem[4] : _GEN_4997; // @[Execute.scala 117:10]
  assign _GEN_4999 = 6'h5 == _T_474 ? welem[5] : _GEN_4998; // @[Execute.scala 117:10]
  assign _GEN_5000 = 6'h6 == _T_474 ? welem[6] : _GEN_4999; // @[Execute.scala 117:10]
  assign _GEN_5001 = 6'h7 == _T_474 ? welem[7] : _GEN_5000; // @[Execute.scala 117:10]
  assign _GEN_5002 = 6'h8 == _T_474 ? welem[8] : _GEN_5001; // @[Execute.scala 117:10]
  assign _GEN_5003 = 6'h9 == _T_474 ? welem[9] : _GEN_5002; // @[Execute.scala 117:10]
  assign _GEN_5004 = 6'ha == _T_474 ? welem[10] : _GEN_5003; // @[Execute.scala 117:10]
  assign _GEN_5005 = 6'hb == _T_474 ? welem[11] : _GEN_5004; // @[Execute.scala 117:10]
  assign _GEN_5006 = 6'hc == _T_474 ? welem[12] : _GEN_5005; // @[Execute.scala 117:10]
  assign _GEN_5007 = 6'hd == _T_474 ? welem[13] : _GEN_5006; // @[Execute.scala 117:10]
  assign _GEN_5008 = 6'he == _T_474 ? welem[14] : _GEN_5007; // @[Execute.scala 117:10]
  assign _GEN_5009 = 6'hf == _T_474 ? welem[15] : _GEN_5008; // @[Execute.scala 117:10]
  assign _GEN_5010 = 6'h10 == _T_474 ? welem[16] : _GEN_5009; // @[Execute.scala 117:10]
  assign _GEN_5011 = 6'h11 == _T_474 ? welem[17] : _GEN_5010; // @[Execute.scala 117:10]
  assign _GEN_5012 = 6'h12 == _T_474 ? welem[18] : _GEN_5011; // @[Execute.scala 117:10]
  assign _GEN_5013 = 6'h13 == _T_474 ? welem[19] : _GEN_5012; // @[Execute.scala 117:10]
  assign _GEN_5014 = 6'h14 == _T_474 ? welem[20] : _GEN_5013; // @[Execute.scala 117:10]
  assign _GEN_5015 = 6'h15 == _T_474 ? welem[21] : _GEN_5014; // @[Execute.scala 117:10]
  assign _GEN_5016 = 6'h16 == _T_474 ? welem[22] : _GEN_5015; // @[Execute.scala 117:10]
  assign _GEN_5017 = 6'h17 == _T_474 ? welem[23] : _GEN_5016; // @[Execute.scala 117:10]
  assign _GEN_5018 = 6'h18 == _T_474 ? welem[24] : _GEN_5017; // @[Execute.scala 117:10]
  assign _GEN_5019 = 6'h19 == _T_474 ? welem[25] : _GEN_5018; // @[Execute.scala 117:10]
  assign _GEN_5020 = 6'h1a == _T_474 ? welem[26] : _GEN_5019; // @[Execute.scala 117:10]
  assign _GEN_5021 = 6'h1b == _T_474 ? welem[27] : _GEN_5020; // @[Execute.scala 117:10]
  assign _GEN_5022 = 6'h1c == _T_474 ? welem[28] : _GEN_5021; // @[Execute.scala 117:10]
  assign _GEN_5023 = 6'h1d == _T_474 ? welem[29] : _GEN_5022; // @[Execute.scala 117:10]
  assign _GEN_5024 = 6'h1e == _T_474 ? welem[30] : _GEN_5023; // @[Execute.scala 117:10]
  assign _GEN_5025 = 6'h1f == _T_474 ? welem[31] : _GEN_5024; // @[Execute.scala 117:10]
  assign _GEN_5026 = 6'h20 == _T_474 ? welem[32] : _GEN_5025; // @[Execute.scala 117:10]
  assign _GEN_5027 = 6'h21 == _T_474 ? welem[33] : _GEN_5026; // @[Execute.scala 117:10]
  assign _GEN_5028 = 6'h22 == _T_474 ? welem[34] : _GEN_5027; // @[Execute.scala 117:10]
  assign _GEN_5029 = 6'h23 == _T_474 ? welem[35] : _GEN_5028; // @[Execute.scala 117:10]
  assign _GEN_5030 = 6'h24 == _T_474 ? welem[36] : _GEN_5029; // @[Execute.scala 117:10]
  assign _GEN_5031 = 6'h25 == _T_474 ? welem[37] : _GEN_5030; // @[Execute.scala 117:10]
  assign _GEN_5032 = 6'h26 == _T_474 ? welem[38] : _GEN_5031; // @[Execute.scala 117:10]
  assign _GEN_5033 = 6'h27 == _T_474 ? welem[39] : _GEN_5032; // @[Execute.scala 117:10]
  assign _GEN_5034 = 6'h28 == _T_474 ? welem[40] : _GEN_5033; // @[Execute.scala 117:10]
  assign _GEN_5035 = 6'h29 == _T_474 ? welem[41] : _GEN_5034; // @[Execute.scala 117:10]
  assign _GEN_5036 = 6'h2a == _T_474 ? welem[42] : _GEN_5035; // @[Execute.scala 117:10]
  assign _GEN_5037 = 6'h2b == _T_474 ? welem[43] : _GEN_5036; // @[Execute.scala 117:10]
  assign _GEN_5038 = 6'h2c == _T_474 ? welem[44] : _GEN_5037; // @[Execute.scala 117:10]
  assign _GEN_5039 = 6'h2d == _T_474 ? welem[45] : _GEN_5038; // @[Execute.scala 117:10]
  assign _GEN_5040 = 6'h2e == _T_474 ? welem[46] : _GEN_5039; // @[Execute.scala 117:10]
  assign _GEN_5041 = 6'h2f == _T_474 ? welem[47] : _GEN_5040; // @[Execute.scala 117:10]
  assign _GEN_5042 = 6'h30 == _T_474 ? welem[48] : _GEN_5041; // @[Execute.scala 117:10]
  assign _GEN_5043 = 6'h31 == _T_474 ? welem[49] : _GEN_5042; // @[Execute.scala 117:10]
  assign _GEN_5044 = 6'h32 == _T_474 ? welem[50] : _GEN_5043; // @[Execute.scala 117:10]
  assign _GEN_5045 = 6'h33 == _T_474 ? welem[51] : _GEN_5044; // @[Execute.scala 117:10]
  assign _GEN_5046 = 6'h34 == _T_474 ? welem[52] : _GEN_5045; // @[Execute.scala 117:10]
  assign _GEN_5047 = 6'h35 == _T_474 ? welem[53] : _GEN_5046; // @[Execute.scala 117:10]
  assign _GEN_5048 = 6'h36 == _T_474 ? welem[54] : _GEN_5047; // @[Execute.scala 117:10]
  assign _GEN_5049 = 6'h37 == _T_474 ? welem[55] : _GEN_5048; // @[Execute.scala 117:10]
  assign _GEN_5050 = 6'h38 == _T_474 ? welem[56] : _GEN_5049; // @[Execute.scala 117:10]
  assign _GEN_5051 = 6'h39 == _T_474 ? welem[57] : _GEN_5050; // @[Execute.scala 117:10]
  assign _GEN_5052 = 6'h3a == _T_474 ? welem[58] : _GEN_5051; // @[Execute.scala 117:10]
  assign _GEN_5053 = 6'h3b == _T_474 ? welem[59] : _GEN_5052; // @[Execute.scala 117:10]
  assign _GEN_5054 = 6'h3c == _T_474 ? welem[60] : _GEN_5053; // @[Execute.scala 117:10]
  assign _GEN_5055 = 6'h3d == _T_474 ? welem[61] : _GEN_5054; // @[Execute.scala 117:10]
  assign _GEN_5056 = 6'h3e == _T_474 ? welem[62] : _GEN_5055; // @[Execute.scala 117:10]
  assign _GEN_5057 = 6'h3f == _T_474 ? welem[63] : _GEN_5056; // @[Execute.scala 117:10]
  assign _GEN_5059 = 6'h1 == _T_478 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5060 = 6'h2 == _T_478 ? welem[2] : _GEN_5059; // @[Execute.scala 117:10]
  assign _GEN_5061 = 6'h3 == _T_478 ? welem[3] : _GEN_5060; // @[Execute.scala 117:10]
  assign _GEN_5062 = 6'h4 == _T_478 ? welem[4] : _GEN_5061; // @[Execute.scala 117:10]
  assign _GEN_5063 = 6'h5 == _T_478 ? welem[5] : _GEN_5062; // @[Execute.scala 117:10]
  assign _GEN_5064 = 6'h6 == _T_478 ? welem[6] : _GEN_5063; // @[Execute.scala 117:10]
  assign _GEN_5065 = 6'h7 == _T_478 ? welem[7] : _GEN_5064; // @[Execute.scala 117:10]
  assign _GEN_5066 = 6'h8 == _T_478 ? welem[8] : _GEN_5065; // @[Execute.scala 117:10]
  assign _GEN_5067 = 6'h9 == _T_478 ? welem[9] : _GEN_5066; // @[Execute.scala 117:10]
  assign _GEN_5068 = 6'ha == _T_478 ? welem[10] : _GEN_5067; // @[Execute.scala 117:10]
  assign _GEN_5069 = 6'hb == _T_478 ? welem[11] : _GEN_5068; // @[Execute.scala 117:10]
  assign _GEN_5070 = 6'hc == _T_478 ? welem[12] : _GEN_5069; // @[Execute.scala 117:10]
  assign _GEN_5071 = 6'hd == _T_478 ? welem[13] : _GEN_5070; // @[Execute.scala 117:10]
  assign _GEN_5072 = 6'he == _T_478 ? welem[14] : _GEN_5071; // @[Execute.scala 117:10]
  assign _GEN_5073 = 6'hf == _T_478 ? welem[15] : _GEN_5072; // @[Execute.scala 117:10]
  assign _GEN_5074 = 6'h10 == _T_478 ? welem[16] : _GEN_5073; // @[Execute.scala 117:10]
  assign _GEN_5075 = 6'h11 == _T_478 ? welem[17] : _GEN_5074; // @[Execute.scala 117:10]
  assign _GEN_5076 = 6'h12 == _T_478 ? welem[18] : _GEN_5075; // @[Execute.scala 117:10]
  assign _GEN_5077 = 6'h13 == _T_478 ? welem[19] : _GEN_5076; // @[Execute.scala 117:10]
  assign _GEN_5078 = 6'h14 == _T_478 ? welem[20] : _GEN_5077; // @[Execute.scala 117:10]
  assign _GEN_5079 = 6'h15 == _T_478 ? welem[21] : _GEN_5078; // @[Execute.scala 117:10]
  assign _GEN_5080 = 6'h16 == _T_478 ? welem[22] : _GEN_5079; // @[Execute.scala 117:10]
  assign _GEN_5081 = 6'h17 == _T_478 ? welem[23] : _GEN_5080; // @[Execute.scala 117:10]
  assign _GEN_5082 = 6'h18 == _T_478 ? welem[24] : _GEN_5081; // @[Execute.scala 117:10]
  assign _GEN_5083 = 6'h19 == _T_478 ? welem[25] : _GEN_5082; // @[Execute.scala 117:10]
  assign _GEN_5084 = 6'h1a == _T_478 ? welem[26] : _GEN_5083; // @[Execute.scala 117:10]
  assign _GEN_5085 = 6'h1b == _T_478 ? welem[27] : _GEN_5084; // @[Execute.scala 117:10]
  assign _GEN_5086 = 6'h1c == _T_478 ? welem[28] : _GEN_5085; // @[Execute.scala 117:10]
  assign _GEN_5087 = 6'h1d == _T_478 ? welem[29] : _GEN_5086; // @[Execute.scala 117:10]
  assign _GEN_5088 = 6'h1e == _T_478 ? welem[30] : _GEN_5087; // @[Execute.scala 117:10]
  assign _GEN_5089 = 6'h1f == _T_478 ? welem[31] : _GEN_5088; // @[Execute.scala 117:10]
  assign _GEN_5090 = 6'h20 == _T_478 ? welem[32] : _GEN_5089; // @[Execute.scala 117:10]
  assign _GEN_5091 = 6'h21 == _T_478 ? welem[33] : _GEN_5090; // @[Execute.scala 117:10]
  assign _GEN_5092 = 6'h22 == _T_478 ? welem[34] : _GEN_5091; // @[Execute.scala 117:10]
  assign _GEN_5093 = 6'h23 == _T_478 ? welem[35] : _GEN_5092; // @[Execute.scala 117:10]
  assign _GEN_5094 = 6'h24 == _T_478 ? welem[36] : _GEN_5093; // @[Execute.scala 117:10]
  assign _GEN_5095 = 6'h25 == _T_478 ? welem[37] : _GEN_5094; // @[Execute.scala 117:10]
  assign _GEN_5096 = 6'h26 == _T_478 ? welem[38] : _GEN_5095; // @[Execute.scala 117:10]
  assign _GEN_5097 = 6'h27 == _T_478 ? welem[39] : _GEN_5096; // @[Execute.scala 117:10]
  assign _GEN_5098 = 6'h28 == _T_478 ? welem[40] : _GEN_5097; // @[Execute.scala 117:10]
  assign _GEN_5099 = 6'h29 == _T_478 ? welem[41] : _GEN_5098; // @[Execute.scala 117:10]
  assign _GEN_5100 = 6'h2a == _T_478 ? welem[42] : _GEN_5099; // @[Execute.scala 117:10]
  assign _GEN_5101 = 6'h2b == _T_478 ? welem[43] : _GEN_5100; // @[Execute.scala 117:10]
  assign _GEN_5102 = 6'h2c == _T_478 ? welem[44] : _GEN_5101; // @[Execute.scala 117:10]
  assign _GEN_5103 = 6'h2d == _T_478 ? welem[45] : _GEN_5102; // @[Execute.scala 117:10]
  assign _GEN_5104 = 6'h2e == _T_478 ? welem[46] : _GEN_5103; // @[Execute.scala 117:10]
  assign _GEN_5105 = 6'h2f == _T_478 ? welem[47] : _GEN_5104; // @[Execute.scala 117:10]
  assign _GEN_5106 = 6'h30 == _T_478 ? welem[48] : _GEN_5105; // @[Execute.scala 117:10]
  assign _GEN_5107 = 6'h31 == _T_478 ? welem[49] : _GEN_5106; // @[Execute.scala 117:10]
  assign _GEN_5108 = 6'h32 == _T_478 ? welem[50] : _GEN_5107; // @[Execute.scala 117:10]
  assign _GEN_5109 = 6'h33 == _T_478 ? welem[51] : _GEN_5108; // @[Execute.scala 117:10]
  assign _GEN_5110 = 6'h34 == _T_478 ? welem[52] : _GEN_5109; // @[Execute.scala 117:10]
  assign _GEN_5111 = 6'h35 == _T_478 ? welem[53] : _GEN_5110; // @[Execute.scala 117:10]
  assign _GEN_5112 = 6'h36 == _T_478 ? welem[54] : _GEN_5111; // @[Execute.scala 117:10]
  assign _GEN_5113 = 6'h37 == _T_478 ? welem[55] : _GEN_5112; // @[Execute.scala 117:10]
  assign _GEN_5114 = 6'h38 == _T_478 ? welem[56] : _GEN_5113; // @[Execute.scala 117:10]
  assign _GEN_5115 = 6'h39 == _T_478 ? welem[57] : _GEN_5114; // @[Execute.scala 117:10]
  assign _GEN_5116 = 6'h3a == _T_478 ? welem[58] : _GEN_5115; // @[Execute.scala 117:10]
  assign _GEN_5117 = 6'h3b == _T_478 ? welem[59] : _GEN_5116; // @[Execute.scala 117:10]
  assign _GEN_5118 = 6'h3c == _T_478 ? welem[60] : _GEN_5117; // @[Execute.scala 117:10]
  assign _GEN_5119 = 6'h3d == _T_478 ? welem[61] : _GEN_5118; // @[Execute.scala 117:10]
  assign _GEN_5120 = 6'h3e == _T_478 ? welem[62] : _GEN_5119; // @[Execute.scala 117:10]
  assign _GEN_5121 = 6'h3f == _T_478 ? welem[63] : _GEN_5120; // @[Execute.scala 117:10]
  assign _T_481 = _T_472 ? _GEN_5057 : _GEN_5121; // @[Execute.scala 117:10]
  assign _T_482 = r < 6'h19; // @[Execute.scala 117:15]
  assign _T_484 = r - 6'h19; // @[Execute.scala 117:37]
  assign _T_488 = 6'h27 + r; // @[Execute.scala 117:60]
  assign _GEN_5123 = 6'h1 == _T_484 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5124 = 6'h2 == _T_484 ? welem[2] : _GEN_5123; // @[Execute.scala 117:10]
  assign _GEN_5125 = 6'h3 == _T_484 ? welem[3] : _GEN_5124; // @[Execute.scala 117:10]
  assign _GEN_5126 = 6'h4 == _T_484 ? welem[4] : _GEN_5125; // @[Execute.scala 117:10]
  assign _GEN_5127 = 6'h5 == _T_484 ? welem[5] : _GEN_5126; // @[Execute.scala 117:10]
  assign _GEN_5128 = 6'h6 == _T_484 ? welem[6] : _GEN_5127; // @[Execute.scala 117:10]
  assign _GEN_5129 = 6'h7 == _T_484 ? welem[7] : _GEN_5128; // @[Execute.scala 117:10]
  assign _GEN_5130 = 6'h8 == _T_484 ? welem[8] : _GEN_5129; // @[Execute.scala 117:10]
  assign _GEN_5131 = 6'h9 == _T_484 ? welem[9] : _GEN_5130; // @[Execute.scala 117:10]
  assign _GEN_5132 = 6'ha == _T_484 ? welem[10] : _GEN_5131; // @[Execute.scala 117:10]
  assign _GEN_5133 = 6'hb == _T_484 ? welem[11] : _GEN_5132; // @[Execute.scala 117:10]
  assign _GEN_5134 = 6'hc == _T_484 ? welem[12] : _GEN_5133; // @[Execute.scala 117:10]
  assign _GEN_5135 = 6'hd == _T_484 ? welem[13] : _GEN_5134; // @[Execute.scala 117:10]
  assign _GEN_5136 = 6'he == _T_484 ? welem[14] : _GEN_5135; // @[Execute.scala 117:10]
  assign _GEN_5137 = 6'hf == _T_484 ? welem[15] : _GEN_5136; // @[Execute.scala 117:10]
  assign _GEN_5138 = 6'h10 == _T_484 ? welem[16] : _GEN_5137; // @[Execute.scala 117:10]
  assign _GEN_5139 = 6'h11 == _T_484 ? welem[17] : _GEN_5138; // @[Execute.scala 117:10]
  assign _GEN_5140 = 6'h12 == _T_484 ? welem[18] : _GEN_5139; // @[Execute.scala 117:10]
  assign _GEN_5141 = 6'h13 == _T_484 ? welem[19] : _GEN_5140; // @[Execute.scala 117:10]
  assign _GEN_5142 = 6'h14 == _T_484 ? welem[20] : _GEN_5141; // @[Execute.scala 117:10]
  assign _GEN_5143 = 6'h15 == _T_484 ? welem[21] : _GEN_5142; // @[Execute.scala 117:10]
  assign _GEN_5144 = 6'h16 == _T_484 ? welem[22] : _GEN_5143; // @[Execute.scala 117:10]
  assign _GEN_5145 = 6'h17 == _T_484 ? welem[23] : _GEN_5144; // @[Execute.scala 117:10]
  assign _GEN_5146 = 6'h18 == _T_484 ? welem[24] : _GEN_5145; // @[Execute.scala 117:10]
  assign _GEN_5147 = 6'h19 == _T_484 ? welem[25] : _GEN_5146; // @[Execute.scala 117:10]
  assign _GEN_5148 = 6'h1a == _T_484 ? welem[26] : _GEN_5147; // @[Execute.scala 117:10]
  assign _GEN_5149 = 6'h1b == _T_484 ? welem[27] : _GEN_5148; // @[Execute.scala 117:10]
  assign _GEN_5150 = 6'h1c == _T_484 ? welem[28] : _GEN_5149; // @[Execute.scala 117:10]
  assign _GEN_5151 = 6'h1d == _T_484 ? welem[29] : _GEN_5150; // @[Execute.scala 117:10]
  assign _GEN_5152 = 6'h1e == _T_484 ? welem[30] : _GEN_5151; // @[Execute.scala 117:10]
  assign _GEN_5153 = 6'h1f == _T_484 ? welem[31] : _GEN_5152; // @[Execute.scala 117:10]
  assign _GEN_5154 = 6'h20 == _T_484 ? welem[32] : _GEN_5153; // @[Execute.scala 117:10]
  assign _GEN_5155 = 6'h21 == _T_484 ? welem[33] : _GEN_5154; // @[Execute.scala 117:10]
  assign _GEN_5156 = 6'h22 == _T_484 ? welem[34] : _GEN_5155; // @[Execute.scala 117:10]
  assign _GEN_5157 = 6'h23 == _T_484 ? welem[35] : _GEN_5156; // @[Execute.scala 117:10]
  assign _GEN_5158 = 6'h24 == _T_484 ? welem[36] : _GEN_5157; // @[Execute.scala 117:10]
  assign _GEN_5159 = 6'h25 == _T_484 ? welem[37] : _GEN_5158; // @[Execute.scala 117:10]
  assign _GEN_5160 = 6'h26 == _T_484 ? welem[38] : _GEN_5159; // @[Execute.scala 117:10]
  assign _GEN_5161 = 6'h27 == _T_484 ? welem[39] : _GEN_5160; // @[Execute.scala 117:10]
  assign _GEN_5162 = 6'h28 == _T_484 ? welem[40] : _GEN_5161; // @[Execute.scala 117:10]
  assign _GEN_5163 = 6'h29 == _T_484 ? welem[41] : _GEN_5162; // @[Execute.scala 117:10]
  assign _GEN_5164 = 6'h2a == _T_484 ? welem[42] : _GEN_5163; // @[Execute.scala 117:10]
  assign _GEN_5165 = 6'h2b == _T_484 ? welem[43] : _GEN_5164; // @[Execute.scala 117:10]
  assign _GEN_5166 = 6'h2c == _T_484 ? welem[44] : _GEN_5165; // @[Execute.scala 117:10]
  assign _GEN_5167 = 6'h2d == _T_484 ? welem[45] : _GEN_5166; // @[Execute.scala 117:10]
  assign _GEN_5168 = 6'h2e == _T_484 ? welem[46] : _GEN_5167; // @[Execute.scala 117:10]
  assign _GEN_5169 = 6'h2f == _T_484 ? welem[47] : _GEN_5168; // @[Execute.scala 117:10]
  assign _GEN_5170 = 6'h30 == _T_484 ? welem[48] : _GEN_5169; // @[Execute.scala 117:10]
  assign _GEN_5171 = 6'h31 == _T_484 ? welem[49] : _GEN_5170; // @[Execute.scala 117:10]
  assign _GEN_5172 = 6'h32 == _T_484 ? welem[50] : _GEN_5171; // @[Execute.scala 117:10]
  assign _GEN_5173 = 6'h33 == _T_484 ? welem[51] : _GEN_5172; // @[Execute.scala 117:10]
  assign _GEN_5174 = 6'h34 == _T_484 ? welem[52] : _GEN_5173; // @[Execute.scala 117:10]
  assign _GEN_5175 = 6'h35 == _T_484 ? welem[53] : _GEN_5174; // @[Execute.scala 117:10]
  assign _GEN_5176 = 6'h36 == _T_484 ? welem[54] : _GEN_5175; // @[Execute.scala 117:10]
  assign _GEN_5177 = 6'h37 == _T_484 ? welem[55] : _GEN_5176; // @[Execute.scala 117:10]
  assign _GEN_5178 = 6'h38 == _T_484 ? welem[56] : _GEN_5177; // @[Execute.scala 117:10]
  assign _GEN_5179 = 6'h39 == _T_484 ? welem[57] : _GEN_5178; // @[Execute.scala 117:10]
  assign _GEN_5180 = 6'h3a == _T_484 ? welem[58] : _GEN_5179; // @[Execute.scala 117:10]
  assign _GEN_5181 = 6'h3b == _T_484 ? welem[59] : _GEN_5180; // @[Execute.scala 117:10]
  assign _GEN_5182 = 6'h3c == _T_484 ? welem[60] : _GEN_5181; // @[Execute.scala 117:10]
  assign _GEN_5183 = 6'h3d == _T_484 ? welem[61] : _GEN_5182; // @[Execute.scala 117:10]
  assign _GEN_5184 = 6'h3e == _T_484 ? welem[62] : _GEN_5183; // @[Execute.scala 117:10]
  assign _GEN_5185 = 6'h3f == _T_484 ? welem[63] : _GEN_5184; // @[Execute.scala 117:10]
  assign _GEN_5187 = 6'h1 == _T_488 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5188 = 6'h2 == _T_488 ? welem[2] : _GEN_5187; // @[Execute.scala 117:10]
  assign _GEN_5189 = 6'h3 == _T_488 ? welem[3] : _GEN_5188; // @[Execute.scala 117:10]
  assign _GEN_5190 = 6'h4 == _T_488 ? welem[4] : _GEN_5189; // @[Execute.scala 117:10]
  assign _GEN_5191 = 6'h5 == _T_488 ? welem[5] : _GEN_5190; // @[Execute.scala 117:10]
  assign _GEN_5192 = 6'h6 == _T_488 ? welem[6] : _GEN_5191; // @[Execute.scala 117:10]
  assign _GEN_5193 = 6'h7 == _T_488 ? welem[7] : _GEN_5192; // @[Execute.scala 117:10]
  assign _GEN_5194 = 6'h8 == _T_488 ? welem[8] : _GEN_5193; // @[Execute.scala 117:10]
  assign _GEN_5195 = 6'h9 == _T_488 ? welem[9] : _GEN_5194; // @[Execute.scala 117:10]
  assign _GEN_5196 = 6'ha == _T_488 ? welem[10] : _GEN_5195; // @[Execute.scala 117:10]
  assign _GEN_5197 = 6'hb == _T_488 ? welem[11] : _GEN_5196; // @[Execute.scala 117:10]
  assign _GEN_5198 = 6'hc == _T_488 ? welem[12] : _GEN_5197; // @[Execute.scala 117:10]
  assign _GEN_5199 = 6'hd == _T_488 ? welem[13] : _GEN_5198; // @[Execute.scala 117:10]
  assign _GEN_5200 = 6'he == _T_488 ? welem[14] : _GEN_5199; // @[Execute.scala 117:10]
  assign _GEN_5201 = 6'hf == _T_488 ? welem[15] : _GEN_5200; // @[Execute.scala 117:10]
  assign _GEN_5202 = 6'h10 == _T_488 ? welem[16] : _GEN_5201; // @[Execute.scala 117:10]
  assign _GEN_5203 = 6'h11 == _T_488 ? welem[17] : _GEN_5202; // @[Execute.scala 117:10]
  assign _GEN_5204 = 6'h12 == _T_488 ? welem[18] : _GEN_5203; // @[Execute.scala 117:10]
  assign _GEN_5205 = 6'h13 == _T_488 ? welem[19] : _GEN_5204; // @[Execute.scala 117:10]
  assign _GEN_5206 = 6'h14 == _T_488 ? welem[20] : _GEN_5205; // @[Execute.scala 117:10]
  assign _GEN_5207 = 6'h15 == _T_488 ? welem[21] : _GEN_5206; // @[Execute.scala 117:10]
  assign _GEN_5208 = 6'h16 == _T_488 ? welem[22] : _GEN_5207; // @[Execute.scala 117:10]
  assign _GEN_5209 = 6'h17 == _T_488 ? welem[23] : _GEN_5208; // @[Execute.scala 117:10]
  assign _GEN_5210 = 6'h18 == _T_488 ? welem[24] : _GEN_5209; // @[Execute.scala 117:10]
  assign _GEN_5211 = 6'h19 == _T_488 ? welem[25] : _GEN_5210; // @[Execute.scala 117:10]
  assign _GEN_5212 = 6'h1a == _T_488 ? welem[26] : _GEN_5211; // @[Execute.scala 117:10]
  assign _GEN_5213 = 6'h1b == _T_488 ? welem[27] : _GEN_5212; // @[Execute.scala 117:10]
  assign _GEN_5214 = 6'h1c == _T_488 ? welem[28] : _GEN_5213; // @[Execute.scala 117:10]
  assign _GEN_5215 = 6'h1d == _T_488 ? welem[29] : _GEN_5214; // @[Execute.scala 117:10]
  assign _GEN_5216 = 6'h1e == _T_488 ? welem[30] : _GEN_5215; // @[Execute.scala 117:10]
  assign _GEN_5217 = 6'h1f == _T_488 ? welem[31] : _GEN_5216; // @[Execute.scala 117:10]
  assign _GEN_5218 = 6'h20 == _T_488 ? welem[32] : _GEN_5217; // @[Execute.scala 117:10]
  assign _GEN_5219 = 6'h21 == _T_488 ? welem[33] : _GEN_5218; // @[Execute.scala 117:10]
  assign _GEN_5220 = 6'h22 == _T_488 ? welem[34] : _GEN_5219; // @[Execute.scala 117:10]
  assign _GEN_5221 = 6'h23 == _T_488 ? welem[35] : _GEN_5220; // @[Execute.scala 117:10]
  assign _GEN_5222 = 6'h24 == _T_488 ? welem[36] : _GEN_5221; // @[Execute.scala 117:10]
  assign _GEN_5223 = 6'h25 == _T_488 ? welem[37] : _GEN_5222; // @[Execute.scala 117:10]
  assign _GEN_5224 = 6'h26 == _T_488 ? welem[38] : _GEN_5223; // @[Execute.scala 117:10]
  assign _GEN_5225 = 6'h27 == _T_488 ? welem[39] : _GEN_5224; // @[Execute.scala 117:10]
  assign _GEN_5226 = 6'h28 == _T_488 ? welem[40] : _GEN_5225; // @[Execute.scala 117:10]
  assign _GEN_5227 = 6'h29 == _T_488 ? welem[41] : _GEN_5226; // @[Execute.scala 117:10]
  assign _GEN_5228 = 6'h2a == _T_488 ? welem[42] : _GEN_5227; // @[Execute.scala 117:10]
  assign _GEN_5229 = 6'h2b == _T_488 ? welem[43] : _GEN_5228; // @[Execute.scala 117:10]
  assign _GEN_5230 = 6'h2c == _T_488 ? welem[44] : _GEN_5229; // @[Execute.scala 117:10]
  assign _GEN_5231 = 6'h2d == _T_488 ? welem[45] : _GEN_5230; // @[Execute.scala 117:10]
  assign _GEN_5232 = 6'h2e == _T_488 ? welem[46] : _GEN_5231; // @[Execute.scala 117:10]
  assign _GEN_5233 = 6'h2f == _T_488 ? welem[47] : _GEN_5232; // @[Execute.scala 117:10]
  assign _GEN_5234 = 6'h30 == _T_488 ? welem[48] : _GEN_5233; // @[Execute.scala 117:10]
  assign _GEN_5235 = 6'h31 == _T_488 ? welem[49] : _GEN_5234; // @[Execute.scala 117:10]
  assign _GEN_5236 = 6'h32 == _T_488 ? welem[50] : _GEN_5235; // @[Execute.scala 117:10]
  assign _GEN_5237 = 6'h33 == _T_488 ? welem[51] : _GEN_5236; // @[Execute.scala 117:10]
  assign _GEN_5238 = 6'h34 == _T_488 ? welem[52] : _GEN_5237; // @[Execute.scala 117:10]
  assign _GEN_5239 = 6'h35 == _T_488 ? welem[53] : _GEN_5238; // @[Execute.scala 117:10]
  assign _GEN_5240 = 6'h36 == _T_488 ? welem[54] : _GEN_5239; // @[Execute.scala 117:10]
  assign _GEN_5241 = 6'h37 == _T_488 ? welem[55] : _GEN_5240; // @[Execute.scala 117:10]
  assign _GEN_5242 = 6'h38 == _T_488 ? welem[56] : _GEN_5241; // @[Execute.scala 117:10]
  assign _GEN_5243 = 6'h39 == _T_488 ? welem[57] : _GEN_5242; // @[Execute.scala 117:10]
  assign _GEN_5244 = 6'h3a == _T_488 ? welem[58] : _GEN_5243; // @[Execute.scala 117:10]
  assign _GEN_5245 = 6'h3b == _T_488 ? welem[59] : _GEN_5244; // @[Execute.scala 117:10]
  assign _GEN_5246 = 6'h3c == _T_488 ? welem[60] : _GEN_5245; // @[Execute.scala 117:10]
  assign _GEN_5247 = 6'h3d == _T_488 ? welem[61] : _GEN_5246; // @[Execute.scala 117:10]
  assign _GEN_5248 = 6'h3e == _T_488 ? welem[62] : _GEN_5247; // @[Execute.scala 117:10]
  assign _GEN_5249 = 6'h3f == _T_488 ? welem[63] : _GEN_5248; // @[Execute.scala 117:10]
  assign _T_491 = _T_482 ? _GEN_5185 : _GEN_5249; // @[Execute.scala 117:10]
  assign _T_492 = r < 6'h18; // @[Execute.scala 117:15]
  assign _T_494 = r - 6'h18; // @[Execute.scala 117:37]
  assign _T_498 = 6'h28 + r; // @[Execute.scala 117:60]
  assign _GEN_5251 = 6'h1 == _T_494 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5252 = 6'h2 == _T_494 ? welem[2] : _GEN_5251; // @[Execute.scala 117:10]
  assign _GEN_5253 = 6'h3 == _T_494 ? welem[3] : _GEN_5252; // @[Execute.scala 117:10]
  assign _GEN_5254 = 6'h4 == _T_494 ? welem[4] : _GEN_5253; // @[Execute.scala 117:10]
  assign _GEN_5255 = 6'h5 == _T_494 ? welem[5] : _GEN_5254; // @[Execute.scala 117:10]
  assign _GEN_5256 = 6'h6 == _T_494 ? welem[6] : _GEN_5255; // @[Execute.scala 117:10]
  assign _GEN_5257 = 6'h7 == _T_494 ? welem[7] : _GEN_5256; // @[Execute.scala 117:10]
  assign _GEN_5258 = 6'h8 == _T_494 ? welem[8] : _GEN_5257; // @[Execute.scala 117:10]
  assign _GEN_5259 = 6'h9 == _T_494 ? welem[9] : _GEN_5258; // @[Execute.scala 117:10]
  assign _GEN_5260 = 6'ha == _T_494 ? welem[10] : _GEN_5259; // @[Execute.scala 117:10]
  assign _GEN_5261 = 6'hb == _T_494 ? welem[11] : _GEN_5260; // @[Execute.scala 117:10]
  assign _GEN_5262 = 6'hc == _T_494 ? welem[12] : _GEN_5261; // @[Execute.scala 117:10]
  assign _GEN_5263 = 6'hd == _T_494 ? welem[13] : _GEN_5262; // @[Execute.scala 117:10]
  assign _GEN_5264 = 6'he == _T_494 ? welem[14] : _GEN_5263; // @[Execute.scala 117:10]
  assign _GEN_5265 = 6'hf == _T_494 ? welem[15] : _GEN_5264; // @[Execute.scala 117:10]
  assign _GEN_5266 = 6'h10 == _T_494 ? welem[16] : _GEN_5265; // @[Execute.scala 117:10]
  assign _GEN_5267 = 6'h11 == _T_494 ? welem[17] : _GEN_5266; // @[Execute.scala 117:10]
  assign _GEN_5268 = 6'h12 == _T_494 ? welem[18] : _GEN_5267; // @[Execute.scala 117:10]
  assign _GEN_5269 = 6'h13 == _T_494 ? welem[19] : _GEN_5268; // @[Execute.scala 117:10]
  assign _GEN_5270 = 6'h14 == _T_494 ? welem[20] : _GEN_5269; // @[Execute.scala 117:10]
  assign _GEN_5271 = 6'h15 == _T_494 ? welem[21] : _GEN_5270; // @[Execute.scala 117:10]
  assign _GEN_5272 = 6'h16 == _T_494 ? welem[22] : _GEN_5271; // @[Execute.scala 117:10]
  assign _GEN_5273 = 6'h17 == _T_494 ? welem[23] : _GEN_5272; // @[Execute.scala 117:10]
  assign _GEN_5274 = 6'h18 == _T_494 ? welem[24] : _GEN_5273; // @[Execute.scala 117:10]
  assign _GEN_5275 = 6'h19 == _T_494 ? welem[25] : _GEN_5274; // @[Execute.scala 117:10]
  assign _GEN_5276 = 6'h1a == _T_494 ? welem[26] : _GEN_5275; // @[Execute.scala 117:10]
  assign _GEN_5277 = 6'h1b == _T_494 ? welem[27] : _GEN_5276; // @[Execute.scala 117:10]
  assign _GEN_5278 = 6'h1c == _T_494 ? welem[28] : _GEN_5277; // @[Execute.scala 117:10]
  assign _GEN_5279 = 6'h1d == _T_494 ? welem[29] : _GEN_5278; // @[Execute.scala 117:10]
  assign _GEN_5280 = 6'h1e == _T_494 ? welem[30] : _GEN_5279; // @[Execute.scala 117:10]
  assign _GEN_5281 = 6'h1f == _T_494 ? welem[31] : _GEN_5280; // @[Execute.scala 117:10]
  assign _GEN_5282 = 6'h20 == _T_494 ? welem[32] : _GEN_5281; // @[Execute.scala 117:10]
  assign _GEN_5283 = 6'h21 == _T_494 ? welem[33] : _GEN_5282; // @[Execute.scala 117:10]
  assign _GEN_5284 = 6'h22 == _T_494 ? welem[34] : _GEN_5283; // @[Execute.scala 117:10]
  assign _GEN_5285 = 6'h23 == _T_494 ? welem[35] : _GEN_5284; // @[Execute.scala 117:10]
  assign _GEN_5286 = 6'h24 == _T_494 ? welem[36] : _GEN_5285; // @[Execute.scala 117:10]
  assign _GEN_5287 = 6'h25 == _T_494 ? welem[37] : _GEN_5286; // @[Execute.scala 117:10]
  assign _GEN_5288 = 6'h26 == _T_494 ? welem[38] : _GEN_5287; // @[Execute.scala 117:10]
  assign _GEN_5289 = 6'h27 == _T_494 ? welem[39] : _GEN_5288; // @[Execute.scala 117:10]
  assign _GEN_5290 = 6'h28 == _T_494 ? welem[40] : _GEN_5289; // @[Execute.scala 117:10]
  assign _GEN_5291 = 6'h29 == _T_494 ? welem[41] : _GEN_5290; // @[Execute.scala 117:10]
  assign _GEN_5292 = 6'h2a == _T_494 ? welem[42] : _GEN_5291; // @[Execute.scala 117:10]
  assign _GEN_5293 = 6'h2b == _T_494 ? welem[43] : _GEN_5292; // @[Execute.scala 117:10]
  assign _GEN_5294 = 6'h2c == _T_494 ? welem[44] : _GEN_5293; // @[Execute.scala 117:10]
  assign _GEN_5295 = 6'h2d == _T_494 ? welem[45] : _GEN_5294; // @[Execute.scala 117:10]
  assign _GEN_5296 = 6'h2e == _T_494 ? welem[46] : _GEN_5295; // @[Execute.scala 117:10]
  assign _GEN_5297 = 6'h2f == _T_494 ? welem[47] : _GEN_5296; // @[Execute.scala 117:10]
  assign _GEN_5298 = 6'h30 == _T_494 ? welem[48] : _GEN_5297; // @[Execute.scala 117:10]
  assign _GEN_5299 = 6'h31 == _T_494 ? welem[49] : _GEN_5298; // @[Execute.scala 117:10]
  assign _GEN_5300 = 6'h32 == _T_494 ? welem[50] : _GEN_5299; // @[Execute.scala 117:10]
  assign _GEN_5301 = 6'h33 == _T_494 ? welem[51] : _GEN_5300; // @[Execute.scala 117:10]
  assign _GEN_5302 = 6'h34 == _T_494 ? welem[52] : _GEN_5301; // @[Execute.scala 117:10]
  assign _GEN_5303 = 6'h35 == _T_494 ? welem[53] : _GEN_5302; // @[Execute.scala 117:10]
  assign _GEN_5304 = 6'h36 == _T_494 ? welem[54] : _GEN_5303; // @[Execute.scala 117:10]
  assign _GEN_5305 = 6'h37 == _T_494 ? welem[55] : _GEN_5304; // @[Execute.scala 117:10]
  assign _GEN_5306 = 6'h38 == _T_494 ? welem[56] : _GEN_5305; // @[Execute.scala 117:10]
  assign _GEN_5307 = 6'h39 == _T_494 ? welem[57] : _GEN_5306; // @[Execute.scala 117:10]
  assign _GEN_5308 = 6'h3a == _T_494 ? welem[58] : _GEN_5307; // @[Execute.scala 117:10]
  assign _GEN_5309 = 6'h3b == _T_494 ? welem[59] : _GEN_5308; // @[Execute.scala 117:10]
  assign _GEN_5310 = 6'h3c == _T_494 ? welem[60] : _GEN_5309; // @[Execute.scala 117:10]
  assign _GEN_5311 = 6'h3d == _T_494 ? welem[61] : _GEN_5310; // @[Execute.scala 117:10]
  assign _GEN_5312 = 6'h3e == _T_494 ? welem[62] : _GEN_5311; // @[Execute.scala 117:10]
  assign _GEN_5313 = 6'h3f == _T_494 ? welem[63] : _GEN_5312; // @[Execute.scala 117:10]
  assign _GEN_5315 = 6'h1 == _T_498 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5316 = 6'h2 == _T_498 ? welem[2] : _GEN_5315; // @[Execute.scala 117:10]
  assign _GEN_5317 = 6'h3 == _T_498 ? welem[3] : _GEN_5316; // @[Execute.scala 117:10]
  assign _GEN_5318 = 6'h4 == _T_498 ? welem[4] : _GEN_5317; // @[Execute.scala 117:10]
  assign _GEN_5319 = 6'h5 == _T_498 ? welem[5] : _GEN_5318; // @[Execute.scala 117:10]
  assign _GEN_5320 = 6'h6 == _T_498 ? welem[6] : _GEN_5319; // @[Execute.scala 117:10]
  assign _GEN_5321 = 6'h7 == _T_498 ? welem[7] : _GEN_5320; // @[Execute.scala 117:10]
  assign _GEN_5322 = 6'h8 == _T_498 ? welem[8] : _GEN_5321; // @[Execute.scala 117:10]
  assign _GEN_5323 = 6'h9 == _T_498 ? welem[9] : _GEN_5322; // @[Execute.scala 117:10]
  assign _GEN_5324 = 6'ha == _T_498 ? welem[10] : _GEN_5323; // @[Execute.scala 117:10]
  assign _GEN_5325 = 6'hb == _T_498 ? welem[11] : _GEN_5324; // @[Execute.scala 117:10]
  assign _GEN_5326 = 6'hc == _T_498 ? welem[12] : _GEN_5325; // @[Execute.scala 117:10]
  assign _GEN_5327 = 6'hd == _T_498 ? welem[13] : _GEN_5326; // @[Execute.scala 117:10]
  assign _GEN_5328 = 6'he == _T_498 ? welem[14] : _GEN_5327; // @[Execute.scala 117:10]
  assign _GEN_5329 = 6'hf == _T_498 ? welem[15] : _GEN_5328; // @[Execute.scala 117:10]
  assign _GEN_5330 = 6'h10 == _T_498 ? welem[16] : _GEN_5329; // @[Execute.scala 117:10]
  assign _GEN_5331 = 6'h11 == _T_498 ? welem[17] : _GEN_5330; // @[Execute.scala 117:10]
  assign _GEN_5332 = 6'h12 == _T_498 ? welem[18] : _GEN_5331; // @[Execute.scala 117:10]
  assign _GEN_5333 = 6'h13 == _T_498 ? welem[19] : _GEN_5332; // @[Execute.scala 117:10]
  assign _GEN_5334 = 6'h14 == _T_498 ? welem[20] : _GEN_5333; // @[Execute.scala 117:10]
  assign _GEN_5335 = 6'h15 == _T_498 ? welem[21] : _GEN_5334; // @[Execute.scala 117:10]
  assign _GEN_5336 = 6'h16 == _T_498 ? welem[22] : _GEN_5335; // @[Execute.scala 117:10]
  assign _GEN_5337 = 6'h17 == _T_498 ? welem[23] : _GEN_5336; // @[Execute.scala 117:10]
  assign _GEN_5338 = 6'h18 == _T_498 ? welem[24] : _GEN_5337; // @[Execute.scala 117:10]
  assign _GEN_5339 = 6'h19 == _T_498 ? welem[25] : _GEN_5338; // @[Execute.scala 117:10]
  assign _GEN_5340 = 6'h1a == _T_498 ? welem[26] : _GEN_5339; // @[Execute.scala 117:10]
  assign _GEN_5341 = 6'h1b == _T_498 ? welem[27] : _GEN_5340; // @[Execute.scala 117:10]
  assign _GEN_5342 = 6'h1c == _T_498 ? welem[28] : _GEN_5341; // @[Execute.scala 117:10]
  assign _GEN_5343 = 6'h1d == _T_498 ? welem[29] : _GEN_5342; // @[Execute.scala 117:10]
  assign _GEN_5344 = 6'h1e == _T_498 ? welem[30] : _GEN_5343; // @[Execute.scala 117:10]
  assign _GEN_5345 = 6'h1f == _T_498 ? welem[31] : _GEN_5344; // @[Execute.scala 117:10]
  assign _GEN_5346 = 6'h20 == _T_498 ? welem[32] : _GEN_5345; // @[Execute.scala 117:10]
  assign _GEN_5347 = 6'h21 == _T_498 ? welem[33] : _GEN_5346; // @[Execute.scala 117:10]
  assign _GEN_5348 = 6'h22 == _T_498 ? welem[34] : _GEN_5347; // @[Execute.scala 117:10]
  assign _GEN_5349 = 6'h23 == _T_498 ? welem[35] : _GEN_5348; // @[Execute.scala 117:10]
  assign _GEN_5350 = 6'h24 == _T_498 ? welem[36] : _GEN_5349; // @[Execute.scala 117:10]
  assign _GEN_5351 = 6'h25 == _T_498 ? welem[37] : _GEN_5350; // @[Execute.scala 117:10]
  assign _GEN_5352 = 6'h26 == _T_498 ? welem[38] : _GEN_5351; // @[Execute.scala 117:10]
  assign _GEN_5353 = 6'h27 == _T_498 ? welem[39] : _GEN_5352; // @[Execute.scala 117:10]
  assign _GEN_5354 = 6'h28 == _T_498 ? welem[40] : _GEN_5353; // @[Execute.scala 117:10]
  assign _GEN_5355 = 6'h29 == _T_498 ? welem[41] : _GEN_5354; // @[Execute.scala 117:10]
  assign _GEN_5356 = 6'h2a == _T_498 ? welem[42] : _GEN_5355; // @[Execute.scala 117:10]
  assign _GEN_5357 = 6'h2b == _T_498 ? welem[43] : _GEN_5356; // @[Execute.scala 117:10]
  assign _GEN_5358 = 6'h2c == _T_498 ? welem[44] : _GEN_5357; // @[Execute.scala 117:10]
  assign _GEN_5359 = 6'h2d == _T_498 ? welem[45] : _GEN_5358; // @[Execute.scala 117:10]
  assign _GEN_5360 = 6'h2e == _T_498 ? welem[46] : _GEN_5359; // @[Execute.scala 117:10]
  assign _GEN_5361 = 6'h2f == _T_498 ? welem[47] : _GEN_5360; // @[Execute.scala 117:10]
  assign _GEN_5362 = 6'h30 == _T_498 ? welem[48] : _GEN_5361; // @[Execute.scala 117:10]
  assign _GEN_5363 = 6'h31 == _T_498 ? welem[49] : _GEN_5362; // @[Execute.scala 117:10]
  assign _GEN_5364 = 6'h32 == _T_498 ? welem[50] : _GEN_5363; // @[Execute.scala 117:10]
  assign _GEN_5365 = 6'h33 == _T_498 ? welem[51] : _GEN_5364; // @[Execute.scala 117:10]
  assign _GEN_5366 = 6'h34 == _T_498 ? welem[52] : _GEN_5365; // @[Execute.scala 117:10]
  assign _GEN_5367 = 6'h35 == _T_498 ? welem[53] : _GEN_5366; // @[Execute.scala 117:10]
  assign _GEN_5368 = 6'h36 == _T_498 ? welem[54] : _GEN_5367; // @[Execute.scala 117:10]
  assign _GEN_5369 = 6'h37 == _T_498 ? welem[55] : _GEN_5368; // @[Execute.scala 117:10]
  assign _GEN_5370 = 6'h38 == _T_498 ? welem[56] : _GEN_5369; // @[Execute.scala 117:10]
  assign _GEN_5371 = 6'h39 == _T_498 ? welem[57] : _GEN_5370; // @[Execute.scala 117:10]
  assign _GEN_5372 = 6'h3a == _T_498 ? welem[58] : _GEN_5371; // @[Execute.scala 117:10]
  assign _GEN_5373 = 6'h3b == _T_498 ? welem[59] : _GEN_5372; // @[Execute.scala 117:10]
  assign _GEN_5374 = 6'h3c == _T_498 ? welem[60] : _GEN_5373; // @[Execute.scala 117:10]
  assign _GEN_5375 = 6'h3d == _T_498 ? welem[61] : _GEN_5374; // @[Execute.scala 117:10]
  assign _GEN_5376 = 6'h3e == _T_498 ? welem[62] : _GEN_5375; // @[Execute.scala 117:10]
  assign _GEN_5377 = 6'h3f == _T_498 ? welem[63] : _GEN_5376; // @[Execute.scala 117:10]
  assign _T_501 = _T_492 ? _GEN_5313 : _GEN_5377; // @[Execute.scala 117:10]
  assign _T_502 = r < 6'h17; // @[Execute.scala 117:15]
  assign _T_504 = r - 6'h17; // @[Execute.scala 117:37]
  assign _T_508 = 6'h29 + r; // @[Execute.scala 117:60]
  assign _GEN_5379 = 6'h1 == _T_504 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5380 = 6'h2 == _T_504 ? welem[2] : _GEN_5379; // @[Execute.scala 117:10]
  assign _GEN_5381 = 6'h3 == _T_504 ? welem[3] : _GEN_5380; // @[Execute.scala 117:10]
  assign _GEN_5382 = 6'h4 == _T_504 ? welem[4] : _GEN_5381; // @[Execute.scala 117:10]
  assign _GEN_5383 = 6'h5 == _T_504 ? welem[5] : _GEN_5382; // @[Execute.scala 117:10]
  assign _GEN_5384 = 6'h6 == _T_504 ? welem[6] : _GEN_5383; // @[Execute.scala 117:10]
  assign _GEN_5385 = 6'h7 == _T_504 ? welem[7] : _GEN_5384; // @[Execute.scala 117:10]
  assign _GEN_5386 = 6'h8 == _T_504 ? welem[8] : _GEN_5385; // @[Execute.scala 117:10]
  assign _GEN_5387 = 6'h9 == _T_504 ? welem[9] : _GEN_5386; // @[Execute.scala 117:10]
  assign _GEN_5388 = 6'ha == _T_504 ? welem[10] : _GEN_5387; // @[Execute.scala 117:10]
  assign _GEN_5389 = 6'hb == _T_504 ? welem[11] : _GEN_5388; // @[Execute.scala 117:10]
  assign _GEN_5390 = 6'hc == _T_504 ? welem[12] : _GEN_5389; // @[Execute.scala 117:10]
  assign _GEN_5391 = 6'hd == _T_504 ? welem[13] : _GEN_5390; // @[Execute.scala 117:10]
  assign _GEN_5392 = 6'he == _T_504 ? welem[14] : _GEN_5391; // @[Execute.scala 117:10]
  assign _GEN_5393 = 6'hf == _T_504 ? welem[15] : _GEN_5392; // @[Execute.scala 117:10]
  assign _GEN_5394 = 6'h10 == _T_504 ? welem[16] : _GEN_5393; // @[Execute.scala 117:10]
  assign _GEN_5395 = 6'h11 == _T_504 ? welem[17] : _GEN_5394; // @[Execute.scala 117:10]
  assign _GEN_5396 = 6'h12 == _T_504 ? welem[18] : _GEN_5395; // @[Execute.scala 117:10]
  assign _GEN_5397 = 6'h13 == _T_504 ? welem[19] : _GEN_5396; // @[Execute.scala 117:10]
  assign _GEN_5398 = 6'h14 == _T_504 ? welem[20] : _GEN_5397; // @[Execute.scala 117:10]
  assign _GEN_5399 = 6'h15 == _T_504 ? welem[21] : _GEN_5398; // @[Execute.scala 117:10]
  assign _GEN_5400 = 6'h16 == _T_504 ? welem[22] : _GEN_5399; // @[Execute.scala 117:10]
  assign _GEN_5401 = 6'h17 == _T_504 ? welem[23] : _GEN_5400; // @[Execute.scala 117:10]
  assign _GEN_5402 = 6'h18 == _T_504 ? welem[24] : _GEN_5401; // @[Execute.scala 117:10]
  assign _GEN_5403 = 6'h19 == _T_504 ? welem[25] : _GEN_5402; // @[Execute.scala 117:10]
  assign _GEN_5404 = 6'h1a == _T_504 ? welem[26] : _GEN_5403; // @[Execute.scala 117:10]
  assign _GEN_5405 = 6'h1b == _T_504 ? welem[27] : _GEN_5404; // @[Execute.scala 117:10]
  assign _GEN_5406 = 6'h1c == _T_504 ? welem[28] : _GEN_5405; // @[Execute.scala 117:10]
  assign _GEN_5407 = 6'h1d == _T_504 ? welem[29] : _GEN_5406; // @[Execute.scala 117:10]
  assign _GEN_5408 = 6'h1e == _T_504 ? welem[30] : _GEN_5407; // @[Execute.scala 117:10]
  assign _GEN_5409 = 6'h1f == _T_504 ? welem[31] : _GEN_5408; // @[Execute.scala 117:10]
  assign _GEN_5410 = 6'h20 == _T_504 ? welem[32] : _GEN_5409; // @[Execute.scala 117:10]
  assign _GEN_5411 = 6'h21 == _T_504 ? welem[33] : _GEN_5410; // @[Execute.scala 117:10]
  assign _GEN_5412 = 6'h22 == _T_504 ? welem[34] : _GEN_5411; // @[Execute.scala 117:10]
  assign _GEN_5413 = 6'h23 == _T_504 ? welem[35] : _GEN_5412; // @[Execute.scala 117:10]
  assign _GEN_5414 = 6'h24 == _T_504 ? welem[36] : _GEN_5413; // @[Execute.scala 117:10]
  assign _GEN_5415 = 6'h25 == _T_504 ? welem[37] : _GEN_5414; // @[Execute.scala 117:10]
  assign _GEN_5416 = 6'h26 == _T_504 ? welem[38] : _GEN_5415; // @[Execute.scala 117:10]
  assign _GEN_5417 = 6'h27 == _T_504 ? welem[39] : _GEN_5416; // @[Execute.scala 117:10]
  assign _GEN_5418 = 6'h28 == _T_504 ? welem[40] : _GEN_5417; // @[Execute.scala 117:10]
  assign _GEN_5419 = 6'h29 == _T_504 ? welem[41] : _GEN_5418; // @[Execute.scala 117:10]
  assign _GEN_5420 = 6'h2a == _T_504 ? welem[42] : _GEN_5419; // @[Execute.scala 117:10]
  assign _GEN_5421 = 6'h2b == _T_504 ? welem[43] : _GEN_5420; // @[Execute.scala 117:10]
  assign _GEN_5422 = 6'h2c == _T_504 ? welem[44] : _GEN_5421; // @[Execute.scala 117:10]
  assign _GEN_5423 = 6'h2d == _T_504 ? welem[45] : _GEN_5422; // @[Execute.scala 117:10]
  assign _GEN_5424 = 6'h2e == _T_504 ? welem[46] : _GEN_5423; // @[Execute.scala 117:10]
  assign _GEN_5425 = 6'h2f == _T_504 ? welem[47] : _GEN_5424; // @[Execute.scala 117:10]
  assign _GEN_5426 = 6'h30 == _T_504 ? welem[48] : _GEN_5425; // @[Execute.scala 117:10]
  assign _GEN_5427 = 6'h31 == _T_504 ? welem[49] : _GEN_5426; // @[Execute.scala 117:10]
  assign _GEN_5428 = 6'h32 == _T_504 ? welem[50] : _GEN_5427; // @[Execute.scala 117:10]
  assign _GEN_5429 = 6'h33 == _T_504 ? welem[51] : _GEN_5428; // @[Execute.scala 117:10]
  assign _GEN_5430 = 6'h34 == _T_504 ? welem[52] : _GEN_5429; // @[Execute.scala 117:10]
  assign _GEN_5431 = 6'h35 == _T_504 ? welem[53] : _GEN_5430; // @[Execute.scala 117:10]
  assign _GEN_5432 = 6'h36 == _T_504 ? welem[54] : _GEN_5431; // @[Execute.scala 117:10]
  assign _GEN_5433 = 6'h37 == _T_504 ? welem[55] : _GEN_5432; // @[Execute.scala 117:10]
  assign _GEN_5434 = 6'h38 == _T_504 ? welem[56] : _GEN_5433; // @[Execute.scala 117:10]
  assign _GEN_5435 = 6'h39 == _T_504 ? welem[57] : _GEN_5434; // @[Execute.scala 117:10]
  assign _GEN_5436 = 6'h3a == _T_504 ? welem[58] : _GEN_5435; // @[Execute.scala 117:10]
  assign _GEN_5437 = 6'h3b == _T_504 ? welem[59] : _GEN_5436; // @[Execute.scala 117:10]
  assign _GEN_5438 = 6'h3c == _T_504 ? welem[60] : _GEN_5437; // @[Execute.scala 117:10]
  assign _GEN_5439 = 6'h3d == _T_504 ? welem[61] : _GEN_5438; // @[Execute.scala 117:10]
  assign _GEN_5440 = 6'h3e == _T_504 ? welem[62] : _GEN_5439; // @[Execute.scala 117:10]
  assign _GEN_5441 = 6'h3f == _T_504 ? welem[63] : _GEN_5440; // @[Execute.scala 117:10]
  assign _GEN_5443 = 6'h1 == _T_508 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5444 = 6'h2 == _T_508 ? welem[2] : _GEN_5443; // @[Execute.scala 117:10]
  assign _GEN_5445 = 6'h3 == _T_508 ? welem[3] : _GEN_5444; // @[Execute.scala 117:10]
  assign _GEN_5446 = 6'h4 == _T_508 ? welem[4] : _GEN_5445; // @[Execute.scala 117:10]
  assign _GEN_5447 = 6'h5 == _T_508 ? welem[5] : _GEN_5446; // @[Execute.scala 117:10]
  assign _GEN_5448 = 6'h6 == _T_508 ? welem[6] : _GEN_5447; // @[Execute.scala 117:10]
  assign _GEN_5449 = 6'h7 == _T_508 ? welem[7] : _GEN_5448; // @[Execute.scala 117:10]
  assign _GEN_5450 = 6'h8 == _T_508 ? welem[8] : _GEN_5449; // @[Execute.scala 117:10]
  assign _GEN_5451 = 6'h9 == _T_508 ? welem[9] : _GEN_5450; // @[Execute.scala 117:10]
  assign _GEN_5452 = 6'ha == _T_508 ? welem[10] : _GEN_5451; // @[Execute.scala 117:10]
  assign _GEN_5453 = 6'hb == _T_508 ? welem[11] : _GEN_5452; // @[Execute.scala 117:10]
  assign _GEN_5454 = 6'hc == _T_508 ? welem[12] : _GEN_5453; // @[Execute.scala 117:10]
  assign _GEN_5455 = 6'hd == _T_508 ? welem[13] : _GEN_5454; // @[Execute.scala 117:10]
  assign _GEN_5456 = 6'he == _T_508 ? welem[14] : _GEN_5455; // @[Execute.scala 117:10]
  assign _GEN_5457 = 6'hf == _T_508 ? welem[15] : _GEN_5456; // @[Execute.scala 117:10]
  assign _GEN_5458 = 6'h10 == _T_508 ? welem[16] : _GEN_5457; // @[Execute.scala 117:10]
  assign _GEN_5459 = 6'h11 == _T_508 ? welem[17] : _GEN_5458; // @[Execute.scala 117:10]
  assign _GEN_5460 = 6'h12 == _T_508 ? welem[18] : _GEN_5459; // @[Execute.scala 117:10]
  assign _GEN_5461 = 6'h13 == _T_508 ? welem[19] : _GEN_5460; // @[Execute.scala 117:10]
  assign _GEN_5462 = 6'h14 == _T_508 ? welem[20] : _GEN_5461; // @[Execute.scala 117:10]
  assign _GEN_5463 = 6'h15 == _T_508 ? welem[21] : _GEN_5462; // @[Execute.scala 117:10]
  assign _GEN_5464 = 6'h16 == _T_508 ? welem[22] : _GEN_5463; // @[Execute.scala 117:10]
  assign _GEN_5465 = 6'h17 == _T_508 ? welem[23] : _GEN_5464; // @[Execute.scala 117:10]
  assign _GEN_5466 = 6'h18 == _T_508 ? welem[24] : _GEN_5465; // @[Execute.scala 117:10]
  assign _GEN_5467 = 6'h19 == _T_508 ? welem[25] : _GEN_5466; // @[Execute.scala 117:10]
  assign _GEN_5468 = 6'h1a == _T_508 ? welem[26] : _GEN_5467; // @[Execute.scala 117:10]
  assign _GEN_5469 = 6'h1b == _T_508 ? welem[27] : _GEN_5468; // @[Execute.scala 117:10]
  assign _GEN_5470 = 6'h1c == _T_508 ? welem[28] : _GEN_5469; // @[Execute.scala 117:10]
  assign _GEN_5471 = 6'h1d == _T_508 ? welem[29] : _GEN_5470; // @[Execute.scala 117:10]
  assign _GEN_5472 = 6'h1e == _T_508 ? welem[30] : _GEN_5471; // @[Execute.scala 117:10]
  assign _GEN_5473 = 6'h1f == _T_508 ? welem[31] : _GEN_5472; // @[Execute.scala 117:10]
  assign _GEN_5474 = 6'h20 == _T_508 ? welem[32] : _GEN_5473; // @[Execute.scala 117:10]
  assign _GEN_5475 = 6'h21 == _T_508 ? welem[33] : _GEN_5474; // @[Execute.scala 117:10]
  assign _GEN_5476 = 6'h22 == _T_508 ? welem[34] : _GEN_5475; // @[Execute.scala 117:10]
  assign _GEN_5477 = 6'h23 == _T_508 ? welem[35] : _GEN_5476; // @[Execute.scala 117:10]
  assign _GEN_5478 = 6'h24 == _T_508 ? welem[36] : _GEN_5477; // @[Execute.scala 117:10]
  assign _GEN_5479 = 6'h25 == _T_508 ? welem[37] : _GEN_5478; // @[Execute.scala 117:10]
  assign _GEN_5480 = 6'h26 == _T_508 ? welem[38] : _GEN_5479; // @[Execute.scala 117:10]
  assign _GEN_5481 = 6'h27 == _T_508 ? welem[39] : _GEN_5480; // @[Execute.scala 117:10]
  assign _GEN_5482 = 6'h28 == _T_508 ? welem[40] : _GEN_5481; // @[Execute.scala 117:10]
  assign _GEN_5483 = 6'h29 == _T_508 ? welem[41] : _GEN_5482; // @[Execute.scala 117:10]
  assign _GEN_5484 = 6'h2a == _T_508 ? welem[42] : _GEN_5483; // @[Execute.scala 117:10]
  assign _GEN_5485 = 6'h2b == _T_508 ? welem[43] : _GEN_5484; // @[Execute.scala 117:10]
  assign _GEN_5486 = 6'h2c == _T_508 ? welem[44] : _GEN_5485; // @[Execute.scala 117:10]
  assign _GEN_5487 = 6'h2d == _T_508 ? welem[45] : _GEN_5486; // @[Execute.scala 117:10]
  assign _GEN_5488 = 6'h2e == _T_508 ? welem[46] : _GEN_5487; // @[Execute.scala 117:10]
  assign _GEN_5489 = 6'h2f == _T_508 ? welem[47] : _GEN_5488; // @[Execute.scala 117:10]
  assign _GEN_5490 = 6'h30 == _T_508 ? welem[48] : _GEN_5489; // @[Execute.scala 117:10]
  assign _GEN_5491 = 6'h31 == _T_508 ? welem[49] : _GEN_5490; // @[Execute.scala 117:10]
  assign _GEN_5492 = 6'h32 == _T_508 ? welem[50] : _GEN_5491; // @[Execute.scala 117:10]
  assign _GEN_5493 = 6'h33 == _T_508 ? welem[51] : _GEN_5492; // @[Execute.scala 117:10]
  assign _GEN_5494 = 6'h34 == _T_508 ? welem[52] : _GEN_5493; // @[Execute.scala 117:10]
  assign _GEN_5495 = 6'h35 == _T_508 ? welem[53] : _GEN_5494; // @[Execute.scala 117:10]
  assign _GEN_5496 = 6'h36 == _T_508 ? welem[54] : _GEN_5495; // @[Execute.scala 117:10]
  assign _GEN_5497 = 6'h37 == _T_508 ? welem[55] : _GEN_5496; // @[Execute.scala 117:10]
  assign _GEN_5498 = 6'h38 == _T_508 ? welem[56] : _GEN_5497; // @[Execute.scala 117:10]
  assign _GEN_5499 = 6'h39 == _T_508 ? welem[57] : _GEN_5498; // @[Execute.scala 117:10]
  assign _GEN_5500 = 6'h3a == _T_508 ? welem[58] : _GEN_5499; // @[Execute.scala 117:10]
  assign _GEN_5501 = 6'h3b == _T_508 ? welem[59] : _GEN_5500; // @[Execute.scala 117:10]
  assign _GEN_5502 = 6'h3c == _T_508 ? welem[60] : _GEN_5501; // @[Execute.scala 117:10]
  assign _GEN_5503 = 6'h3d == _T_508 ? welem[61] : _GEN_5502; // @[Execute.scala 117:10]
  assign _GEN_5504 = 6'h3e == _T_508 ? welem[62] : _GEN_5503; // @[Execute.scala 117:10]
  assign _GEN_5505 = 6'h3f == _T_508 ? welem[63] : _GEN_5504; // @[Execute.scala 117:10]
  assign _T_511 = _T_502 ? _GEN_5441 : _GEN_5505; // @[Execute.scala 117:10]
  assign _T_512 = r < 6'h16; // @[Execute.scala 117:15]
  assign _T_514 = r - 6'h16; // @[Execute.scala 117:37]
  assign _T_518 = 6'h2a + r; // @[Execute.scala 117:60]
  assign _GEN_5507 = 6'h1 == _T_514 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5508 = 6'h2 == _T_514 ? welem[2] : _GEN_5507; // @[Execute.scala 117:10]
  assign _GEN_5509 = 6'h3 == _T_514 ? welem[3] : _GEN_5508; // @[Execute.scala 117:10]
  assign _GEN_5510 = 6'h4 == _T_514 ? welem[4] : _GEN_5509; // @[Execute.scala 117:10]
  assign _GEN_5511 = 6'h5 == _T_514 ? welem[5] : _GEN_5510; // @[Execute.scala 117:10]
  assign _GEN_5512 = 6'h6 == _T_514 ? welem[6] : _GEN_5511; // @[Execute.scala 117:10]
  assign _GEN_5513 = 6'h7 == _T_514 ? welem[7] : _GEN_5512; // @[Execute.scala 117:10]
  assign _GEN_5514 = 6'h8 == _T_514 ? welem[8] : _GEN_5513; // @[Execute.scala 117:10]
  assign _GEN_5515 = 6'h9 == _T_514 ? welem[9] : _GEN_5514; // @[Execute.scala 117:10]
  assign _GEN_5516 = 6'ha == _T_514 ? welem[10] : _GEN_5515; // @[Execute.scala 117:10]
  assign _GEN_5517 = 6'hb == _T_514 ? welem[11] : _GEN_5516; // @[Execute.scala 117:10]
  assign _GEN_5518 = 6'hc == _T_514 ? welem[12] : _GEN_5517; // @[Execute.scala 117:10]
  assign _GEN_5519 = 6'hd == _T_514 ? welem[13] : _GEN_5518; // @[Execute.scala 117:10]
  assign _GEN_5520 = 6'he == _T_514 ? welem[14] : _GEN_5519; // @[Execute.scala 117:10]
  assign _GEN_5521 = 6'hf == _T_514 ? welem[15] : _GEN_5520; // @[Execute.scala 117:10]
  assign _GEN_5522 = 6'h10 == _T_514 ? welem[16] : _GEN_5521; // @[Execute.scala 117:10]
  assign _GEN_5523 = 6'h11 == _T_514 ? welem[17] : _GEN_5522; // @[Execute.scala 117:10]
  assign _GEN_5524 = 6'h12 == _T_514 ? welem[18] : _GEN_5523; // @[Execute.scala 117:10]
  assign _GEN_5525 = 6'h13 == _T_514 ? welem[19] : _GEN_5524; // @[Execute.scala 117:10]
  assign _GEN_5526 = 6'h14 == _T_514 ? welem[20] : _GEN_5525; // @[Execute.scala 117:10]
  assign _GEN_5527 = 6'h15 == _T_514 ? welem[21] : _GEN_5526; // @[Execute.scala 117:10]
  assign _GEN_5528 = 6'h16 == _T_514 ? welem[22] : _GEN_5527; // @[Execute.scala 117:10]
  assign _GEN_5529 = 6'h17 == _T_514 ? welem[23] : _GEN_5528; // @[Execute.scala 117:10]
  assign _GEN_5530 = 6'h18 == _T_514 ? welem[24] : _GEN_5529; // @[Execute.scala 117:10]
  assign _GEN_5531 = 6'h19 == _T_514 ? welem[25] : _GEN_5530; // @[Execute.scala 117:10]
  assign _GEN_5532 = 6'h1a == _T_514 ? welem[26] : _GEN_5531; // @[Execute.scala 117:10]
  assign _GEN_5533 = 6'h1b == _T_514 ? welem[27] : _GEN_5532; // @[Execute.scala 117:10]
  assign _GEN_5534 = 6'h1c == _T_514 ? welem[28] : _GEN_5533; // @[Execute.scala 117:10]
  assign _GEN_5535 = 6'h1d == _T_514 ? welem[29] : _GEN_5534; // @[Execute.scala 117:10]
  assign _GEN_5536 = 6'h1e == _T_514 ? welem[30] : _GEN_5535; // @[Execute.scala 117:10]
  assign _GEN_5537 = 6'h1f == _T_514 ? welem[31] : _GEN_5536; // @[Execute.scala 117:10]
  assign _GEN_5538 = 6'h20 == _T_514 ? welem[32] : _GEN_5537; // @[Execute.scala 117:10]
  assign _GEN_5539 = 6'h21 == _T_514 ? welem[33] : _GEN_5538; // @[Execute.scala 117:10]
  assign _GEN_5540 = 6'h22 == _T_514 ? welem[34] : _GEN_5539; // @[Execute.scala 117:10]
  assign _GEN_5541 = 6'h23 == _T_514 ? welem[35] : _GEN_5540; // @[Execute.scala 117:10]
  assign _GEN_5542 = 6'h24 == _T_514 ? welem[36] : _GEN_5541; // @[Execute.scala 117:10]
  assign _GEN_5543 = 6'h25 == _T_514 ? welem[37] : _GEN_5542; // @[Execute.scala 117:10]
  assign _GEN_5544 = 6'h26 == _T_514 ? welem[38] : _GEN_5543; // @[Execute.scala 117:10]
  assign _GEN_5545 = 6'h27 == _T_514 ? welem[39] : _GEN_5544; // @[Execute.scala 117:10]
  assign _GEN_5546 = 6'h28 == _T_514 ? welem[40] : _GEN_5545; // @[Execute.scala 117:10]
  assign _GEN_5547 = 6'h29 == _T_514 ? welem[41] : _GEN_5546; // @[Execute.scala 117:10]
  assign _GEN_5548 = 6'h2a == _T_514 ? welem[42] : _GEN_5547; // @[Execute.scala 117:10]
  assign _GEN_5549 = 6'h2b == _T_514 ? welem[43] : _GEN_5548; // @[Execute.scala 117:10]
  assign _GEN_5550 = 6'h2c == _T_514 ? welem[44] : _GEN_5549; // @[Execute.scala 117:10]
  assign _GEN_5551 = 6'h2d == _T_514 ? welem[45] : _GEN_5550; // @[Execute.scala 117:10]
  assign _GEN_5552 = 6'h2e == _T_514 ? welem[46] : _GEN_5551; // @[Execute.scala 117:10]
  assign _GEN_5553 = 6'h2f == _T_514 ? welem[47] : _GEN_5552; // @[Execute.scala 117:10]
  assign _GEN_5554 = 6'h30 == _T_514 ? welem[48] : _GEN_5553; // @[Execute.scala 117:10]
  assign _GEN_5555 = 6'h31 == _T_514 ? welem[49] : _GEN_5554; // @[Execute.scala 117:10]
  assign _GEN_5556 = 6'h32 == _T_514 ? welem[50] : _GEN_5555; // @[Execute.scala 117:10]
  assign _GEN_5557 = 6'h33 == _T_514 ? welem[51] : _GEN_5556; // @[Execute.scala 117:10]
  assign _GEN_5558 = 6'h34 == _T_514 ? welem[52] : _GEN_5557; // @[Execute.scala 117:10]
  assign _GEN_5559 = 6'h35 == _T_514 ? welem[53] : _GEN_5558; // @[Execute.scala 117:10]
  assign _GEN_5560 = 6'h36 == _T_514 ? welem[54] : _GEN_5559; // @[Execute.scala 117:10]
  assign _GEN_5561 = 6'h37 == _T_514 ? welem[55] : _GEN_5560; // @[Execute.scala 117:10]
  assign _GEN_5562 = 6'h38 == _T_514 ? welem[56] : _GEN_5561; // @[Execute.scala 117:10]
  assign _GEN_5563 = 6'h39 == _T_514 ? welem[57] : _GEN_5562; // @[Execute.scala 117:10]
  assign _GEN_5564 = 6'h3a == _T_514 ? welem[58] : _GEN_5563; // @[Execute.scala 117:10]
  assign _GEN_5565 = 6'h3b == _T_514 ? welem[59] : _GEN_5564; // @[Execute.scala 117:10]
  assign _GEN_5566 = 6'h3c == _T_514 ? welem[60] : _GEN_5565; // @[Execute.scala 117:10]
  assign _GEN_5567 = 6'h3d == _T_514 ? welem[61] : _GEN_5566; // @[Execute.scala 117:10]
  assign _GEN_5568 = 6'h3e == _T_514 ? welem[62] : _GEN_5567; // @[Execute.scala 117:10]
  assign _GEN_5569 = 6'h3f == _T_514 ? welem[63] : _GEN_5568; // @[Execute.scala 117:10]
  assign _GEN_5571 = 6'h1 == _T_518 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5572 = 6'h2 == _T_518 ? welem[2] : _GEN_5571; // @[Execute.scala 117:10]
  assign _GEN_5573 = 6'h3 == _T_518 ? welem[3] : _GEN_5572; // @[Execute.scala 117:10]
  assign _GEN_5574 = 6'h4 == _T_518 ? welem[4] : _GEN_5573; // @[Execute.scala 117:10]
  assign _GEN_5575 = 6'h5 == _T_518 ? welem[5] : _GEN_5574; // @[Execute.scala 117:10]
  assign _GEN_5576 = 6'h6 == _T_518 ? welem[6] : _GEN_5575; // @[Execute.scala 117:10]
  assign _GEN_5577 = 6'h7 == _T_518 ? welem[7] : _GEN_5576; // @[Execute.scala 117:10]
  assign _GEN_5578 = 6'h8 == _T_518 ? welem[8] : _GEN_5577; // @[Execute.scala 117:10]
  assign _GEN_5579 = 6'h9 == _T_518 ? welem[9] : _GEN_5578; // @[Execute.scala 117:10]
  assign _GEN_5580 = 6'ha == _T_518 ? welem[10] : _GEN_5579; // @[Execute.scala 117:10]
  assign _GEN_5581 = 6'hb == _T_518 ? welem[11] : _GEN_5580; // @[Execute.scala 117:10]
  assign _GEN_5582 = 6'hc == _T_518 ? welem[12] : _GEN_5581; // @[Execute.scala 117:10]
  assign _GEN_5583 = 6'hd == _T_518 ? welem[13] : _GEN_5582; // @[Execute.scala 117:10]
  assign _GEN_5584 = 6'he == _T_518 ? welem[14] : _GEN_5583; // @[Execute.scala 117:10]
  assign _GEN_5585 = 6'hf == _T_518 ? welem[15] : _GEN_5584; // @[Execute.scala 117:10]
  assign _GEN_5586 = 6'h10 == _T_518 ? welem[16] : _GEN_5585; // @[Execute.scala 117:10]
  assign _GEN_5587 = 6'h11 == _T_518 ? welem[17] : _GEN_5586; // @[Execute.scala 117:10]
  assign _GEN_5588 = 6'h12 == _T_518 ? welem[18] : _GEN_5587; // @[Execute.scala 117:10]
  assign _GEN_5589 = 6'h13 == _T_518 ? welem[19] : _GEN_5588; // @[Execute.scala 117:10]
  assign _GEN_5590 = 6'h14 == _T_518 ? welem[20] : _GEN_5589; // @[Execute.scala 117:10]
  assign _GEN_5591 = 6'h15 == _T_518 ? welem[21] : _GEN_5590; // @[Execute.scala 117:10]
  assign _GEN_5592 = 6'h16 == _T_518 ? welem[22] : _GEN_5591; // @[Execute.scala 117:10]
  assign _GEN_5593 = 6'h17 == _T_518 ? welem[23] : _GEN_5592; // @[Execute.scala 117:10]
  assign _GEN_5594 = 6'h18 == _T_518 ? welem[24] : _GEN_5593; // @[Execute.scala 117:10]
  assign _GEN_5595 = 6'h19 == _T_518 ? welem[25] : _GEN_5594; // @[Execute.scala 117:10]
  assign _GEN_5596 = 6'h1a == _T_518 ? welem[26] : _GEN_5595; // @[Execute.scala 117:10]
  assign _GEN_5597 = 6'h1b == _T_518 ? welem[27] : _GEN_5596; // @[Execute.scala 117:10]
  assign _GEN_5598 = 6'h1c == _T_518 ? welem[28] : _GEN_5597; // @[Execute.scala 117:10]
  assign _GEN_5599 = 6'h1d == _T_518 ? welem[29] : _GEN_5598; // @[Execute.scala 117:10]
  assign _GEN_5600 = 6'h1e == _T_518 ? welem[30] : _GEN_5599; // @[Execute.scala 117:10]
  assign _GEN_5601 = 6'h1f == _T_518 ? welem[31] : _GEN_5600; // @[Execute.scala 117:10]
  assign _GEN_5602 = 6'h20 == _T_518 ? welem[32] : _GEN_5601; // @[Execute.scala 117:10]
  assign _GEN_5603 = 6'h21 == _T_518 ? welem[33] : _GEN_5602; // @[Execute.scala 117:10]
  assign _GEN_5604 = 6'h22 == _T_518 ? welem[34] : _GEN_5603; // @[Execute.scala 117:10]
  assign _GEN_5605 = 6'h23 == _T_518 ? welem[35] : _GEN_5604; // @[Execute.scala 117:10]
  assign _GEN_5606 = 6'h24 == _T_518 ? welem[36] : _GEN_5605; // @[Execute.scala 117:10]
  assign _GEN_5607 = 6'h25 == _T_518 ? welem[37] : _GEN_5606; // @[Execute.scala 117:10]
  assign _GEN_5608 = 6'h26 == _T_518 ? welem[38] : _GEN_5607; // @[Execute.scala 117:10]
  assign _GEN_5609 = 6'h27 == _T_518 ? welem[39] : _GEN_5608; // @[Execute.scala 117:10]
  assign _GEN_5610 = 6'h28 == _T_518 ? welem[40] : _GEN_5609; // @[Execute.scala 117:10]
  assign _GEN_5611 = 6'h29 == _T_518 ? welem[41] : _GEN_5610; // @[Execute.scala 117:10]
  assign _GEN_5612 = 6'h2a == _T_518 ? welem[42] : _GEN_5611; // @[Execute.scala 117:10]
  assign _GEN_5613 = 6'h2b == _T_518 ? welem[43] : _GEN_5612; // @[Execute.scala 117:10]
  assign _GEN_5614 = 6'h2c == _T_518 ? welem[44] : _GEN_5613; // @[Execute.scala 117:10]
  assign _GEN_5615 = 6'h2d == _T_518 ? welem[45] : _GEN_5614; // @[Execute.scala 117:10]
  assign _GEN_5616 = 6'h2e == _T_518 ? welem[46] : _GEN_5615; // @[Execute.scala 117:10]
  assign _GEN_5617 = 6'h2f == _T_518 ? welem[47] : _GEN_5616; // @[Execute.scala 117:10]
  assign _GEN_5618 = 6'h30 == _T_518 ? welem[48] : _GEN_5617; // @[Execute.scala 117:10]
  assign _GEN_5619 = 6'h31 == _T_518 ? welem[49] : _GEN_5618; // @[Execute.scala 117:10]
  assign _GEN_5620 = 6'h32 == _T_518 ? welem[50] : _GEN_5619; // @[Execute.scala 117:10]
  assign _GEN_5621 = 6'h33 == _T_518 ? welem[51] : _GEN_5620; // @[Execute.scala 117:10]
  assign _GEN_5622 = 6'h34 == _T_518 ? welem[52] : _GEN_5621; // @[Execute.scala 117:10]
  assign _GEN_5623 = 6'h35 == _T_518 ? welem[53] : _GEN_5622; // @[Execute.scala 117:10]
  assign _GEN_5624 = 6'h36 == _T_518 ? welem[54] : _GEN_5623; // @[Execute.scala 117:10]
  assign _GEN_5625 = 6'h37 == _T_518 ? welem[55] : _GEN_5624; // @[Execute.scala 117:10]
  assign _GEN_5626 = 6'h38 == _T_518 ? welem[56] : _GEN_5625; // @[Execute.scala 117:10]
  assign _GEN_5627 = 6'h39 == _T_518 ? welem[57] : _GEN_5626; // @[Execute.scala 117:10]
  assign _GEN_5628 = 6'h3a == _T_518 ? welem[58] : _GEN_5627; // @[Execute.scala 117:10]
  assign _GEN_5629 = 6'h3b == _T_518 ? welem[59] : _GEN_5628; // @[Execute.scala 117:10]
  assign _GEN_5630 = 6'h3c == _T_518 ? welem[60] : _GEN_5629; // @[Execute.scala 117:10]
  assign _GEN_5631 = 6'h3d == _T_518 ? welem[61] : _GEN_5630; // @[Execute.scala 117:10]
  assign _GEN_5632 = 6'h3e == _T_518 ? welem[62] : _GEN_5631; // @[Execute.scala 117:10]
  assign _GEN_5633 = 6'h3f == _T_518 ? welem[63] : _GEN_5632; // @[Execute.scala 117:10]
  assign _T_521 = _T_512 ? _GEN_5569 : _GEN_5633; // @[Execute.scala 117:10]
  assign _T_522 = r < 6'h15; // @[Execute.scala 117:15]
  assign _T_524 = r - 6'h15; // @[Execute.scala 117:37]
  assign _T_528 = 6'h2b + r; // @[Execute.scala 117:60]
  assign _GEN_5635 = 6'h1 == _T_524 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5636 = 6'h2 == _T_524 ? welem[2] : _GEN_5635; // @[Execute.scala 117:10]
  assign _GEN_5637 = 6'h3 == _T_524 ? welem[3] : _GEN_5636; // @[Execute.scala 117:10]
  assign _GEN_5638 = 6'h4 == _T_524 ? welem[4] : _GEN_5637; // @[Execute.scala 117:10]
  assign _GEN_5639 = 6'h5 == _T_524 ? welem[5] : _GEN_5638; // @[Execute.scala 117:10]
  assign _GEN_5640 = 6'h6 == _T_524 ? welem[6] : _GEN_5639; // @[Execute.scala 117:10]
  assign _GEN_5641 = 6'h7 == _T_524 ? welem[7] : _GEN_5640; // @[Execute.scala 117:10]
  assign _GEN_5642 = 6'h8 == _T_524 ? welem[8] : _GEN_5641; // @[Execute.scala 117:10]
  assign _GEN_5643 = 6'h9 == _T_524 ? welem[9] : _GEN_5642; // @[Execute.scala 117:10]
  assign _GEN_5644 = 6'ha == _T_524 ? welem[10] : _GEN_5643; // @[Execute.scala 117:10]
  assign _GEN_5645 = 6'hb == _T_524 ? welem[11] : _GEN_5644; // @[Execute.scala 117:10]
  assign _GEN_5646 = 6'hc == _T_524 ? welem[12] : _GEN_5645; // @[Execute.scala 117:10]
  assign _GEN_5647 = 6'hd == _T_524 ? welem[13] : _GEN_5646; // @[Execute.scala 117:10]
  assign _GEN_5648 = 6'he == _T_524 ? welem[14] : _GEN_5647; // @[Execute.scala 117:10]
  assign _GEN_5649 = 6'hf == _T_524 ? welem[15] : _GEN_5648; // @[Execute.scala 117:10]
  assign _GEN_5650 = 6'h10 == _T_524 ? welem[16] : _GEN_5649; // @[Execute.scala 117:10]
  assign _GEN_5651 = 6'h11 == _T_524 ? welem[17] : _GEN_5650; // @[Execute.scala 117:10]
  assign _GEN_5652 = 6'h12 == _T_524 ? welem[18] : _GEN_5651; // @[Execute.scala 117:10]
  assign _GEN_5653 = 6'h13 == _T_524 ? welem[19] : _GEN_5652; // @[Execute.scala 117:10]
  assign _GEN_5654 = 6'h14 == _T_524 ? welem[20] : _GEN_5653; // @[Execute.scala 117:10]
  assign _GEN_5655 = 6'h15 == _T_524 ? welem[21] : _GEN_5654; // @[Execute.scala 117:10]
  assign _GEN_5656 = 6'h16 == _T_524 ? welem[22] : _GEN_5655; // @[Execute.scala 117:10]
  assign _GEN_5657 = 6'h17 == _T_524 ? welem[23] : _GEN_5656; // @[Execute.scala 117:10]
  assign _GEN_5658 = 6'h18 == _T_524 ? welem[24] : _GEN_5657; // @[Execute.scala 117:10]
  assign _GEN_5659 = 6'h19 == _T_524 ? welem[25] : _GEN_5658; // @[Execute.scala 117:10]
  assign _GEN_5660 = 6'h1a == _T_524 ? welem[26] : _GEN_5659; // @[Execute.scala 117:10]
  assign _GEN_5661 = 6'h1b == _T_524 ? welem[27] : _GEN_5660; // @[Execute.scala 117:10]
  assign _GEN_5662 = 6'h1c == _T_524 ? welem[28] : _GEN_5661; // @[Execute.scala 117:10]
  assign _GEN_5663 = 6'h1d == _T_524 ? welem[29] : _GEN_5662; // @[Execute.scala 117:10]
  assign _GEN_5664 = 6'h1e == _T_524 ? welem[30] : _GEN_5663; // @[Execute.scala 117:10]
  assign _GEN_5665 = 6'h1f == _T_524 ? welem[31] : _GEN_5664; // @[Execute.scala 117:10]
  assign _GEN_5666 = 6'h20 == _T_524 ? welem[32] : _GEN_5665; // @[Execute.scala 117:10]
  assign _GEN_5667 = 6'h21 == _T_524 ? welem[33] : _GEN_5666; // @[Execute.scala 117:10]
  assign _GEN_5668 = 6'h22 == _T_524 ? welem[34] : _GEN_5667; // @[Execute.scala 117:10]
  assign _GEN_5669 = 6'h23 == _T_524 ? welem[35] : _GEN_5668; // @[Execute.scala 117:10]
  assign _GEN_5670 = 6'h24 == _T_524 ? welem[36] : _GEN_5669; // @[Execute.scala 117:10]
  assign _GEN_5671 = 6'h25 == _T_524 ? welem[37] : _GEN_5670; // @[Execute.scala 117:10]
  assign _GEN_5672 = 6'h26 == _T_524 ? welem[38] : _GEN_5671; // @[Execute.scala 117:10]
  assign _GEN_5673 = 6'h27 == _T_524 ? welem[39] : _GEN_5672; // @[Execute.scala 117:10]
  assign _GEN_5674 = 6'h28 == _T_524 ? welem[40] : _GEN_5673; // @[Execute.scala 117:10]
  assign _GEN_5675 = 6'h29 == _T_524 ? welem[41] : _GEN_5674; // @[Execute.scala 117:10]
  assign _GEN_5676 = 6'h2a == _T_524 ? welem[42] : _GEN_5675; // @[Execute.scala 117:10]
  assign _GEN_5677 = 6'h2b == _T_524 ? welem[43] : _GEN_5676; // @[Execute.scala 117:10]
  assign _GEN_5678 = 6'h2c == _T_524 ? welem[44] : _GEN_5677; // @[Execute.scala 117:10]
  assign _GEN_5679 = 6'h2d == _T_524 ? welem[45] : _GEN_5678; // @[Execute.scala 117:10]
  assign _GEN_5680 = 6'h2e == _T_524 ? welem[46] : _GEN_5679; // @[Execute.scala 117:10]
  assign _GEN_5681 = 6'h2f == _T_524 ? welem[47] : _GEN_5680; // @[Execute.scala 117:10]
  assign _GEN_5682 = 6'h30 == _T_524 ? welem[48] : _GEN_5681; // @[Execute.scala 117:10]
  assign _GEN_5683 = 6'h31 == _T_524 ? welem[49] : _GEN_5682; // @[Execute.scala 117:10]
  assign _GEN_5684 = 6'h32 == _T_524 ? welem[50] : _GEN_5683; // @[Execute.scala 117:10]
  assign _GEN_5685 = 6'h33 == _T_524 ? welem[51] : _GEN_5684; // @[Execute.scala 117:10]
  assign _GEN_5686 = 6'h34 == _T_524 ? welem[52] : _GEN_5685; // @[Execute.scala 117:10]
  assign _GEN_5687 = 6'h35 == _T_524 ? welem[53] : _GEN_5686; // @[Execute.scala 117:10]
  assign _GEN_5688 = 6'h36 == _T_524 ? welem[54] : _GEN_5687; // @[Execute.scala 117:10]
  assign _GEN_5689 = 6'h37 == _T_524 ? welem[55] : _GEN_5688; // @[Execute.scala 117:10]
  assign _GEN_5690 = 6'h38 == _T_524 ? welem[56] : _GEN_5689; // @[Execute.scala 117:10]
  assign _GEN_5691 = 6'h39 == _T_524 ? welem[57] : _GEN_5690; // @[Execute.scala 117:10]
  assign _GEN_5692 = 6'h3a == _T_524 ? welem[58] : _GEN_5691; // @[Execute.scala 117:10]
  assign _GEN_5693 = 6'h3b == _T_524 ? welem[59] : _GEN_5692; // @[Execute.scala 117:10]
  assign _GEN_5694 = 6'h3c == _T_524 ? welem[60] : _GEN_5693; // @[Execute.scala 117:10]
  assign _GEN_5695 = 6'h3d == _T_524 ? welem[61] : _GEN_5694; // @[Execute.scala 117:10]
  assign _GEN_5696 = 6'h3e == _T_524 ? welem[62] : _GEN_5695; // @[Execute.scala 117:10]
  assign _GEN_5697 = 6'h3f == _T_524 ? welem[63] : _GEN_5696; // @[Execute.scala 117:10]
  assign _GEN_5699 = 6'h1 == _T_528 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5700 = 6'h2 == _T_528 ? welem[2] : _GEN_5699; // @[Execute.scala 117:10]
  assign _GEN_5701 = 6'h3 == _T_528 ? welem[3] : _GEN_5700; // @[Execute.scala 117:10]
  assign _GEN_5702 = 6'h4 == _T_528 ? welem[4] : _GEN_5701; // @[Execute.scala 117:10]
  assign _GEN_5703 = 6'h5 == _T_528 ? welem[5] : _GEN_5702; // @[Execute.scala 117:10]
  assign _GEN_5704 = 6'h6 == _T_528 ? welem[6] : _GEN_5703; // @[Execute.scala 117:10]
  assign _GEN_5705 = 6'h7 == _T_528 ? welem[7] : _GEN_5704; // @[Execute.scala 117:10]
  assign _GEN_5706 = 6'h8 == _T_528 ? welem[8] : _GEN_5705; // @[Execute.scala 117:10]
  assign _GEN_5707 = 6'h9 == _T_528 ? welem[9] : _GEN_5706; // @[Execute.scala 117:10]
  assign _GEN_5708 = 6'ha == _T_528 ? welem[10] : _GEN_5707; // @[Execute.scala 117:10]
  assign _GEN_5709 = 6'hb == _T_528 ? welem[11] : _GEN_5708; // @[Execute.scala 117:10]
  assign _GEN_5710 = 6'hc == _T_528 ? welem[12] : _GEN_5709; // @[Execute.scala 117:10]
  assign _GEN_5711 = 6'hd == _T_528 ? welem[13] : _GEN_5710; // @[Execute.scala 117:10]
  assign _GEN_5712 = 6'he == _T_528 ? welem[14] : _GEN_5711; // @[Execute.scala 117:10]
  assign _GEN_5713 = 6'hf == _T_528 ? welem[15] : _GEN_5712; // @[Execute.scala 117:10]
  assign _GEN_5714 = 6'h10 == _T_528 ? welem[16] : _GEN_5713; // @[Execute.scala 117:10]
  assign _GEN_5715 = 6'h11 == _T_528 ? welem[17] : _GEN_5714; // @[Execute.scala 117:10]
  assign _GEN_5716 = 6'h12 == _T_528 ? welem[18] : _GEN_5715; // @[Execute.scala 117:10]
  assign _GEN_5717 = 6'h13 == _T_528 ? welem[19] : _GEN_5716; // @[Execute.scala 117:10]
  assign _GEN_5718 = 6'h14 == _T_528 ? welem[20] : _GEN_5717; // @[Execute.scala 117:10]
  assign _GEN_5719 = 6'h15 == _T_528 ? welem[21] : _GEN_5718; // @[Execute.scala 117:10]
  assign _GEN_5720 = 6'h16 == _T_528 ? welem[22] : _GEN_5719; // @[Execute.scala 117:10]
  assign _GEN_5721 = 6'h17 == _T_528 ? welem[23] : _GEN_5720; // @[Execute.scala 117:10]
  assign _GEN_5722 = 6'h18 == _T_528 ? welem[24] : _GEN_5721; // @[Execute.scala 117:10]
  assign _GEN_5723 = 6'h19 == _T_528 ? welem[25] : _GEN_5722; // @[Execute.scala 117:10]
  assign _GEN_5724 = 6'h1a == _T_528 ? welem[26] : _GEN_5723; // @[Execute.scala 117:10]
  assign _GEN_5725 = 6'h1b == _T_528 ? welem[27] : _GEN_5724; // @[Execute.scala 117:10]
  assign _GEN_5726 = 6'h1c == _T_528 ? welem[28] : _GEN_5725; // @[Execute.scala 117:10]
  assign _GEN_5727 = 6'h1d == _T_528 ? welem[29] : _GEN_5726; // @[Execute.scala 117:10]
  assign _GEN_5728 = 6'h1e == _T_528 ? welem[30] : _GEN_5727; // @[Execute.scala 117:10]
  assign _GEN_5729 = 6'h1f == _T_528 ? welem[31] : _GEN_5728; // @[Execute.scala 117:10]
  assign _GEN_5730 = 6'h20 == _T_528 ? welem[32] : _GEN_5729; // @[Execute.scala 117:10]
  assign _GEN_5731 = 6'h21 == _T_528 ? welem[33] : _GEN_5730; // @[Execute.scala 117:10]
  assign _GEN_5732 = 6'h22 == _T_528 ? welem[34] : _GEN_5731; // @[Execute.scala 117:10]
  assign _GEN_5733 = 6'h23 == _T_528 ? welem[35] : _GEN_5732; // @[Execute.scala 117:10]
  assign _GEN_5734 = 6'h24 == _T_528 ? welem[36] : _GEN_5733; // @[Execute.scala 117:10]
  assign _GEN_5735 = 6'h25 == _T_528 ? welem[37] : _GEN_5734; // @[Execute.scala 117:10]
  assign _GEN_5736 = 6'h26 == _T_528 ? welem[38] : _GEN_5735; // @[Execute.scala 117:10]
  assign _GEN_5737 = 6'h27 == _T_528 ? welem[39] : _GEN_5736; // @[Execute.scala 117:10]
  assign _GEN_5738 = 6'h28 == _T_528 ? welem[40] : _GEN_5737; // @[Execute.scala 117:10]
  assign _GEN_5739 = 6'h29 == _T_528 ? welem[41] : _GEN_5738; // @[Execute.scala 117:10]
  assign _GEN_5740 = 6'h2a == _T_528 ? welem[42] : _GEN_5739; // @[Execute.scala 117:10]
  assign _GEN_5741 = 6'h2b == _T_528 ? welem[43] : _GEN_5740; // @[Execute.scala 117:10]
  assign _GEN_5742 = 6'h2c == _T_528 ? welem[44] : _GEN_5741; // @[Execute.scala 117:10]
  assign _GEN_5743 = 6'h2d == _T_528 ? welem[45] : _GEN_5742; // @[Execute.scala 117:10]
  assign _GEN_5744 = 6'h2e == _T_528 ? welem[46] : _GEN_5743; // @[Execute.scala 117:10]
  assign _GEN_5745 = 6'h2f == _T_528 ? welem[47] : _GEN_5744; // @[Execute.scala 117:10]
  assign _GEN_5746 = 6'h30 == _T_528 ? welem[48] : _GEN_5745; // @[Execute.scala 117:10]
  assign _GEN_5747 = 6'h31 == _T_528 ? welem[49] : _GEN_5746; // @[Execute.scala 117:10]
  assign _GEN_5748 = 6'h32 == _T_528 ? welem[50] : _GEN_5747; // @[Execute.scala 117:10]
  assign _GEN_5749 = 6'h33 == _T_528 ? welem[51] : _GEN_5748; // @[Execute.scala 117:10]
  assign _GEN_5750 = 6'h34 == _T_528 ? welem[52] : _GEN_5749; // @[Execute.scala 117:10]
  assign _GEN_5751 = 6'h35 == _T_528 ? welem[53] : _GEN_5750; // @[Execute.scala 117:10]
  assign _GEN_5752 = 6'h36 == _T_528 ? welem[54] : _GEN_5751; // @[Execute.scala 117:10]
  assign _GEN_5753 = 6'h37 == _T_528 ? welem[55] : _GEN_5752; // @[Execute.scala 117:10]
  assign _GEN_5754 = 6'h38 == _T_528 ? welem[56] : _GEN_5753; // @[Execute.scala 117:10]
  assign _GEN_5755 = 6'h39 == _T_528 ? welem[57] : _GEN_5754; // @[Execute.scala 117:10]
  assign _GEN_5756 = 6'h3a == _T_528 ? welem[58] : _GEN_5755; // @[Execute.scala 117:10]
  assign _GEN_5757 = 6'h3b == _T_528 ? welem[59] : _GEN_5756; // @[Execute.scala 117:10]
  assign _GEN_5758 = 6'h3c == _T_528 ? welem[60] : _GEN_5757; // @[Execute.scala 117:10]
  assign _GEN_5759 = 6'h3d == _T_528 ? welem[61] : _GEN_5758; // @[Execute.scala 117:10]
  assign _GEN_5760 = 6'h3e == _T_528 ? welem[62] : _GEN_5759; // @[Execute.scala 117:10]
  assign _GEN_5761 = 6'h3f == _T_528 ? welem[63] : _GEN_5760; // @[Execute.scala 117:10]
  assign _T_531 = _T_522 ? _GEN_5697 : _GEN_5761; // @[Execute.scala 117:10]
  assign _T_532 = r < 6'h14; // @[Execute.scala 117:15]
  assign _T_534 = r - 6'h14; // @[Execute.scala 117:37]
  assign _T_538 = 6'h2c + r; // @[Execute.scala 117:60]
  assign _GEN_5763 = 6'h1 == _T_534 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5764 = 6'h2 == _T_534 ? welem[2] : _GEN_5763; // @[Execute.scala 117:10]
  assign _GEN_5765 = 6'h3 == _T_534 ? welem[3] : _GEN_5764; // @[Execute.scala 117:10]
  assign _GEN_5766 = 6'h4 == _T_534 ? welem[4] : _GEN_5765; // @[Execute.scala 117:10]
  assign _GEN_5767 = 6'h5 == _T_534 ? welem[5] : _GEN_5766; // @[Execute.scala 117:10]
  assign _GEN_5768 = 6'h6 == _T_534 ? welem[6] : _GEN_5767; // @[Execute.scala 117:10]
  assign _GEN_5769 = 6'h7 == _T_534 ? welem[7] : _GEN_5768; // @[Execute.scala 117:10]
  assign _GEN_5770 = 6'h8 == _T_534 ? welem[8] : _GEN_5769; // @[Execute.scala 117:10]
  assign _GEN_5771 = 6'h9 == _T_534 ? welem[9] : _GEN_5770; // @[Execute.scala 117:10]
  assign _GEN_5772 = 6'ha == _T_534 ? welem[10] : _GEN_5771; // @[Execute.scala 117:10]
  assign _GEN_5773 = 6'hb == _T_534 ? welem[11] : _GEN_5772; // @[Execute.scala 117:10]
  assign _GEN_5774 = 6'hc == _T_534 ? welem[12] : _GEN_5773; // @[Execute.scala 117:10]
  assign _GEN_5775 = 6'hd == _T_534 ? welem[13] : _GEN_5774; // @[Execute.scala 117:10]
  assign _GEN_5776 = 6'he == _T_534 ? welem[14] : _GEN_5775; // @[Execute.scala 117:10]
  assign _GEN_5777 = 6'hf == _T_534 ? welem[15] : _GEN_5776; // @[Execute.scala 117:10]
  assign _GEN_5778 = 6'h10 == _T_534 ? welem[16] : _GEN_5777; // @[Execute.scala 117:10]
  assign _GEN_5779 = 6'h11 == _T_534 ? welem[17] : _GEN_5778; // @[Execute.scala 117:10]
  assign _GEN_5780 = 6'h12 == _T_534 ? welem[18] : _GEN_5779; // @[Execute.scala 117:10]
  assign _GEN_5781 = 6'h13 == _T_534 ? welem[19] : _GEN_5780; // @[Execute.scala 117:10]
  assign _GEN_5782 = 6'h14 == _T_534 ? welem[20] : _GEN_5781; // @[Execute.scala 117:10]
  assign _GEN_5783 = 6'h15 == _T_534 ? welem[21] : _GEN_5782; // @[Execute.scala 117:10]
  assign _GEN_5784 = 6'h16 == _T_534 ? welem[22] : _GEN_5783; // @[Execute.scala 117:10]
  assign _GEN_5785 = 6'h17 == _T_534 ? welem[23] : _GEN_5784; // @[Execute.scala 117:10]
  assign _GEN_5786 = 6'h18 == _T_534 ? welem[24] : _GEN_5785; // @[Execute.scala 117:10]
  assign _GEN_5787 = 6'h19 == _T_534 ? welem[25] : _GEN_5786; // @[Execute.scala 117:10]
  assign _GEN_5788 = 6'h1a == _T_534 ? welem[26] : _GEN_5787; // @[Execute.scala 117:10]
  assign _GEN_5789 = 6'h1b == _T_534 ? welem[27] : _GEN_5788; // @[Execute.scala 117:10]
  assign _GEN_5790 = 6'h1c == _T_534 ? welem[28] : _GEN_5789; // @[Execute.scala 117:10]
  assign _GEN_5791 = 6'h1d == _T_534 ? welem[29] : _GEN_5790; // @[Execute.scala 117:10]
  assign _GEN_5792 = 6'h1e == _T_534 ? welem[30] : _GEN_5791; // @[Execute.scala 117:10]
  assign _GEN_5793 = 6'h1f == _T_534 ? welem[31] : _GEN_5792; // @[Execute.scala 117:10]
  assign _GEN_5794 = 6'h20 == _T_534 ? welem[32] : _GEN_5793; // @[Execute.scala 117:10]
  assign _GEN_5795 = 6'h21 == _T_534 ? welem[33] : _GEN_5794; // @[Execute.scala 117:10]
  assign _GEN_5796 = 6'h22 == _T_534 ? welem[34] : _GEN_5795; // @[Execute.scala 117:10]
  assign _GEN_5797 = 6'h23 == _T_534 ? welem[35] : _GEN_5796; // @[Execute.scala 117:10]
  assign _GEN_5798 = 6'h24 == _T_534 ? welem[36] : _GEN_5797; // @[Execute.scala 117:10]
  assign _GEN_5799 = 6'h25 == _T_534 ? welem[37] : _GEN_5798; // @[Execute.scala 117:10]
  assign _GEN_5800 = 6'h26 == _T_534 ? welem[38] : _GEN_5799; // @[Execute.scala 117:10]
  assign _GEN_5801 = 6'h27 == _T_534 ? welem[39] : _GEN_5800; // @[Execute.scala 117:10]
  assign _GEN_5802 = 6'h28 == _T_534 ? welem[40] : _GEN_5801; // @[Execute.scala 117:10]
  assign _GEN_5803 = 6'h29 == _T_534 ? welem[41] : _GEN_5802; // @[Execute.scala 117:10]
  assign _GEN_5804 = 6'h2a == _T_534 ? welem[42] : _GEN_5803; // @[Execute.scala 117:10]
  assign _GEN_5805 = 6'h2b == _T_534 ? welem[43] : _GEN_5804; // @[Execute.scala 117:10]
  assign _GEN_5806 = 6'h2c == _T_534 ? welem[44] : _GEN_5805; // @[Execute.scala 117:10]
  assign _GEN_5807 = 6'h2d == _T_534 ? welem[45] : _GEN_5806; // @[Execute.scala 117:10]
  assign _GEN_5808 = 6'h2e == _T_534 ? welem[46] : _GEN_5807; // @[Execute.scala 117:10]
  assign _GEN_5809 = 6'h2f == _T_534 ? welem[47] : _GEN_5808; // @[Execute.scala 117:10]
  assign _GEN_5810 = 6'h30 == _T_534 ? welem[48] : _GEN_5809; // @[Execute.scala 117:10]
  assign _GEN_5811 = 6'h31 == _T_534 ? welem[49] : _GEN_5810; // @[Execute.scala 117:10]
  assign _GEN_5812 = 6'h32 == _T_534 ? welem[50] : _GEN_5811; // @[Execute.scala 117:10]
  assign _GEN_5813 = 6'h33 == _T_534 ? welem[51] : _GEN_5812; // @[Execute.scala 117:10]
  assign _GEN_5814 = 6'h34 == _T_534 ? welem[52] : _GEN_5813; // @[Execute.scala 117:10]
  assign _GEN_5815 = 6'h35 == _T_534 ? welem[53] : _GEN_5814; // @[Execute.scala 117:10]
  assign _GEN_5816 = 6'h36 == _T_534 ? welem[54] : _GEN_5815; // @[Execute.scala 117:10]
  assign _GEN_5817 = 6'h37 == _T_534 ? welem[55] : _GEN_5816; // @[Execute.scala 117:10]
  assign _GEN_5818 = 6'h38 == _T_534 ? welem[56] : _GEN_5817; // @[Execute.scala 117:10]
  assign _GEN_5819 = 6'h39 == _T_534 ? welem[57] : _GEN_5818; // @[Execute.scala 117:10]
  assign _GEN_5820 = 6'h3a == _T_534 ? welem[58] : _GEN_5819; // @[Execute.scala 117:10]
  assign _GEN_5821 = 6'h3b == _T_534 ? welem[59] : _GEN_5820; // @[Execute.scala 117:10]
  assign _GEN_5822 = 6'h3c == _T_534 ? welem[60] : _GEN_5821; // @[Execute.scala 117:10]
  assign _GEN_5823 = 6'h3d == _T_534 ? welem[61] : _GEN_5822; // @[Execute.scala 117:10]
  assign _GEN_5824 = 6'h3e == _T_534 ? welem[62] : _GEN_5823; // @[Execute.scala 117:10]
  assign _GEN_5825 = 6'h3f == _T_534 ? welem[63] : _GEN_5824; // @[Execute.scala 117:10]
  assign _GEN_5827 = 6'h1 == _T_538 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5828 = 6'h2 == _T_538 ? welem[2] : _GEN_5827; // @[Execute.scala 117:10]
  assign _GEN_5829 = 6'h3 == _T_538 ? welem[3] : _GEN_5828; // @[Execute.scala 117:10]
  assign _GEN_5830 = 6'h4 == _T_538 ? welem[4] : _GEN_5829; // @[Execute.scala 117:10]
  assign _GEN_5831 = 6'h5 == _T_538 ? welem[5] : _GEN_5830; // @[Execute.scala 117:10]
  assign _GEN_5832 = 6'h6 == _T_538 ? welem[6] : _GEN_5831; // @[Execute.scala 117:10]
  assign _GEN_5833 = 6'h7 == _T_538 ? welem[7] : _GEN_5832; // @[Execute.scala 117:10]
  assign _GEN_5834 = 6'h8 == _T_538 ? welem[8] : _GEN_5833; // @[Execute.scala 117:10]
  assign _GEN_5835 = 6'h9 == _T_538 ? welem[9] : _GEN_5834; // @[Execute.scala 117:10]
  assign _GEN_5836 = 6'ha == _T_538 ? welem[10] : _GEN_5835; // @[Execute.scala 117:10]
  assign _GEN_5837 = 6'hb == _T_538 ? welem[11] : _GEN_5836; // @[Execute.scala 117:10]
  assign _GEN_5838 = 6'hc == _T_538 ? welem[12] : _GEN_5837; // @[Execute.scala 117:10]
  assign _GEN_5839 = 6'hd == _T_538 ? welem[13] : _GEN_5838; // @[Execute.scala 117:10]
  assign _GEN_5840 = 6'he == _T_538 ? welem[14] : _GEN_5839; // @[Execute.scala 117:10]
  assign _GEN_5841 = 6'hf == _T_538 ? welem[15] : _GEN_5840; // @[Execute.scala 117:10]
  assign _GEN_5842 = 6'h10 == _T_538 ? welem[16] : _GEN_5841; // @[Execute.scala 117:10]
  assign _GEN_5843 = 6'h11 == _T_538 ? welem[17] : _GEN_5842; // @[Execute.scala 117:10]
  assign _GEN_5844 = 6'h12 == _T_538 ? welem[18] : _GEN_5843; // @[Execute.scala 117:10]
  assign _GEN_5845 = 6'h13 == _T_538 ? welem[19] : _GEN_5844; // @[Execute.scala 117:10]
  assign _GEN_5846 = 6'h14 == _T_538 ? welem[20] : _GEN_5845; // @[Execute.scala 117:10]
  assign _GEN_5847 = 6'h15 == _T_538 ? welem[21] : _GEN_5846; // @[Execute.scala 117:10]
  assign _GEN_5848 = 6'h16 == _T_538 ? welem[22] : _GEN_5847; // @[Execute.scala 117:10]
  assign _GEN_5849 = 6'h17 == _T_538 ? welem[23] : _GEN_5848; // @[Execute.scala 117:10]
  assign _GEN_5850 = 6'h18 == _T_538 ? welem[24] : _GEN_5849; // @[Execute.scala 117:10]
  assign _GEN_5851 = 6'h19 == _T_538 ? welem[25] : _GEN_5850; // @[Execute.scala 117:10]
  assign _GEN_5852 = 6'h1a == _T_538 ? welem[26] : _GEN_5851; // @[Execute.scala 117:10]
  assign _GEN_5853 = 6'h1b == _T_538 ? welem[27] : _GEN_5852; // @[Execute.scala 117:10]
  assign _GEN_5854 = 6'h1c == _T_538 ? welem[28] : _GEN_5853; // @[Execute.scala 117:10]
  assign _GEN_5855 = 6'h1d == _T_538 ? welem[29] : _GEN_5854; // @[Execute.scala 117:10]
  assign _GEN_5856 = 6'h1e == _T_538 ? welem[30] : _GEN_5855; // @[Execute.scala 117:10]
  assign _GEN_5857 = 6'h1f == _T_538 ? welem[31] : _GEN_5856; // @[Execute.scala 117:10]
  assign _GEN_5858 = 6'h20 == _T_538 ? welem[32] : _GEN_5857; // @[Execute.scala 117:10]
  assign _GEN_5859 = 6'h21 == _T_538 ? welem[33] : _GEN_5858; // @[Execute.scala 117:10]
  assign _GEN_5860 = 6'h22 == _T_538 ? welem[34] : _GEN_5859; // @[Execute.scala 117:10]
  assign _GEN_5861 = 6'h23 == _T_538 ? welem[35] : _GEN_5860; // @[Execute.scala 117:10]
  assign _GEN_5862 = 6'h24 == _T_538 ? welem[36] : _GEN_5861; // @[Execute.scala 117:10]
  assign _GEN_5863 = 6'h25 == _T_538 ? welem[37] : _GEN_5862; // @[Execute.scala 117:10]
  assign _GEN_5864 = 6'h26 == _T_538 ? welem[38] : _GEN_5863; // @[Execute.scala 117:10]
  assign _GEN_5865 = 6'h27 == _T_538 ? welem[39] : _GEN_5864; // @[Execute.scala 117:10]
  assign _GEN_5866 = 6'h28 == _T_538 ? welem[40] : _GEN_5865; // @[Execute.scala 117:10]
  assign _GEN_5867 = 6'h29 == _T_538 ? welem[41] : _GEN_5866; // @[Execute.scala 117:10]
  assign _GEN_5868 = 6'h2a == _T_538 ? welem[42] : _GEN_5867; // @[Execute.scala 117:10]
  assign _GEN_5869 = 6'h2b == _T_538 ? welem[43] : _GEN_5868; // @[Execute.scala 117:10]
  assign _GEN_5870 = 6'h2c == _T_538 ? welem[44] : _GEN_5869; // @[Execute.scala 117:10]
  assign _GEN_5871 = 6'h2d == _T_538 ? welem[45] : _GEN_5870; // @[Execute.scala 117:10]
  assign _GEN_5872 = 6'h2e == _T_538 ? welem[46] : _GEN_5871; // @[Execute.scala 117:10]
  assign _GEN_5873 = 6'h2f == _T_538 ? welem[47] : _GEN_5872; // @[Execute.scala 117:10]
  assign _GEN_5874 = 6'h30 == _T_538 ? welem[48] : _GEN_5873; // @[Execute.scala 117:10]
  assign _GEN_5875 = 6'h31 == _T_538 ? welem[49] : _GEN_5874; // @[Execute.scala 117:10]
  assign _GEN_5876 = 6'h32 == _T_538 ? welem[50] : _GEN_5875; // @[Execute.scala 117:10]
  assign _GEN_5877 = 6'h33 == _T_538 ? welem[51] : _GEN_5876; // @[Execute.scala 117:10]
  assign _GEN_5878 = 6'h34 == _T_538 ? welem[52] : _GEN_5877; // @[Execute.scala 117:10]
  assign _GEN_5879 = 6'h35 == _T_538 ? welem[53] : _GEN_5878; // @[Execute.scala 117:10]
  assign _GEN_5880 = 6'h36 == _T_538 ? welem[54] : _GEN_5879; // @[Execute.scala 117:10]
  assign _GEN_5881 = 6'h37 == _T_538 ? welem[55] : _GEN_5880; // @[Execute.scala 117:10]
  assign _GEN_5882 = 6'h38 == _T_538 ? welem[56] : _GEN_5881; // @[Execute.scala 117:10]
  assign _GEN_5883 = 6'h39 == _T_538 ? welem[57] : _GEN_5882; // @[Execute.scala 117:10]
  assign _GEN_5884 = 6'h3a == _T_538 ? welem[58] : _GEN_5883; // @[Execute.scala 117:10]
  assign _GEN_5885 = 6'h3b == _T_538 ? welem[59] : _GEN_5884; // @[Execute.scala 117:10]
  assign _GEN_5886 = 6'h3c == _T_538 ? welem[60] : _GEN_5885; // @[Execute.scala 117:10]
  assign _GEN_5887 = 6'h3d == _T_538 ? welem[61] : _GEN_5886; // @[Execute.scala 117:10]
  assign _GEN_5888 = 6'h3e == _T_538 ? welem[62] : _GEN_5887; // @[Execute.scala 117:10]
  assign _GEN_5889 = 6'h3f == _T_538 ? welem[63] : _GEN_5888; // @[Execute.scala 117:10]
  assign _T_541 = _T_532 ? _GEN_5825 : _GEN_5889; // @[Execute.scala 117:10]
  assign _T_542 = r < 6'h13; // @[Execute.scala 117:15]
  assign _T_544 = r - 6'h13; // @[Execute.scala 117:37]
  assign _T_548 = 6'h2d + r; // @[Execute.scala 117:60]
  assign _GEN_5891 = 6'h1 == _T_544 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5892 = 6'h2 == _T_544 ? welem[2] : _GEN_5891; // @[Execute.scala 117:10]
  assign _GEN_5893 = 6'h3 == _T_544 ? welem[3] : _GEN_5892; // @[Execute.scala 117:10]
  assign _GEN_5894 = 6'h4 == _T_544 ? welem[4] : _GEN_5893; // @[Execute.scala 117:10]
  assign _GEN_5895 = 6'h5 == _T_544 ? welem[5] : _GEN_5894; // @[Execute.scala 117:10]
  assign _GEN_5896 = 6'h6 == _T_544 ? welem[6] : _GEN_5895; // @[Execute.scala 117:10]
  assign _GEN_5897 = 6'h7 == _T_544 ? welem[7] : _GEN_5896; // @[Execute.scala 117:10]
  assign _GEN_5898 = 6'h8 == _T_544 ? welem[8] : _GEN_5897; // @[Execute.scala 117:10]
  assign _GEN_5899 = 6'h9 == _T_544 ? welem[9] : _GEN_5898; // @[Execute.scala 117:10]
  assign _GEN_5900 = 6'ha == _T_544 ? welem[10] : _GEN_5899; // @[Execute.scala 117:10]
  assign _GEN_5901 = 6'hb == _T_544 ? welem[11] : _GEN_5900; // @[Execute.scala 117:10]
  assign _GEN_5902 = 6'hc == _T_544 ? welem[12] : _GEN_5901; // @[Execute.scala 117:10]
  assign _GEN_5903 = 6'hd == _T_544 ? welem[13] : _GEN_5902; // @[Execute.scala 117:10]
  assign _GEN_5904 = 6'he == _T_544 ? welem[14] : _GEN_5903; // @[Execute.scala 117:10]
  assign _GEN_5905 = 6'hf == _T_544 ? welem[15] : _GEN_5904; // @[Execute.scala 117:10]
  assign _GEN_5906 = 6'h10 == _T_544 ? welem[16] : _GEN_5905; // @[Execute.scala 117:10]
  assign _GEN_5907 = 6'h11 == _T_544 ? welem[17] : _GEN_5906; // @[Execute.scala 117:10]
  assign _GEN_5908 = 6'h12 == _T_544 ? welem[18] : _GEN_5907; // @[Execute.scala 117:10]
  assign _GEN_5909 = 6'h13 == _T_544 ? welem[19] : _GEN_5908; // @[Execute.scala 117:10]
  assign _GEN_5910 = 6'h14 == _T_544 ? welem[20] : _GEN_5909; // @[Execute.scala 117:10]
  assign _GEN_5911 = 6'h15 == _T_544 ? welem[21] : _GEN_5910; // @[Execute.scala 117:10]
  assign _GEN_5912 = 6'h16 == _T_544 ? welem[22] : _GEN_5911; // @[Execute.scala 117:10]
  assign _GEN_5913 = 6'h17 == _T_544 ? welem[23] : _GEN_5912; // @[Execute.scala 117:10]
  assign _GEN_5914 = 6'h18 == _T_544 ? welem[24] : _GEN_5913; // @[Execute.scala 117:10]
  assign _GEN_5915 = 6'h19 == _T_544 ? welem[25] : _GEN_5914; // @[Execute.scala 117:10]
  assign _GEN_5916 = 6'h1a == _T_544 ? welem[26] : _GEN_5915; // @[Execute.scala 117:10]
  assign _GEN_5917 = 6'h1b == _T_544 ? welem[27] : _GEN_5916; // @[Execute.scala 117:10]
  assign _GEN_5918 = 6'h1c == _T_544 ? welem[28] : _GEN_5917; // @[Execute.scala 117:10]
  assign _GEN_5919 = 6'h1d == _T_544 ? welem[29] : _GEN_5918; // @[Execute.scala 117:10]
  assign _GEN_5920 = 6'h1e == _T_544 ? welem[30] : _GEN_5919; // @[Execute.scala 117:10]
  assign _GEN_5921 = 6'h1f == _T_544 ? welem[31] : _GEN_5920; // @[Execute.scala 117:10]
  assign _GEN_5922 = 6'h20 == _T_544 ? welem[32] : _GEN_5921; // @[Execute.scala 117:10]
  assign _GEN_5923 = 6'h21 == _T_544 ? welem[33] : _GEN_5922; // @[Execute.scala 117:10]
  assign _GEN_5924 = 6'h22 == _T_544 ? welem[34] : _GEN_5923; // @[Execute.scala 117:10]
  assign _GEN_5925 = 6'h23 == _T_544 ? welem[35] : _GEN_5924; // @[Execute.scala 117:10]
  assign _GEN_5926 = 6'h24 == _T_544 ? welem[36] : _GEN_5925; // @[Execute.scala 117:10]
  assign _GEN_5927 = 6'h25 == _T_544 ? welem[37] : _GEN_5926; // @[Execute.scala 117:10]
  assign _GEN_5928 = 6'h26 == _T_544 ? welem[38] : _GEN_5927; // @[Execute.scala 117:10]
  assign _GEN_5929 = 6'h27 == _T_544 ? welem[39] : _GEN_5928; // @[Execute.scala 117:10]
  assign _GEN_5930 = 6'h28 == _T_544 ? welem[40] : _GEN_5929; // @[Execute.scala 117:10]
  assign _GEN_5931 = 6'h29 == _T_544 ? welem[41] : _GEN_5930; // @[Execute.scala 117:10]
  assign _GEN_5932 = 6'h2a == _T_544 ? welem[42] : _GEN_5931; // @[Execute.scala 117:10]
  assign _GEN_5933 = 6'h2b == _T_544 ? welem[43] : _GEN_5932; // @[Execute.scala 117:10]
  assign _GEN_5934 = 6'h2c == _T_544 ? welem[44] : _GEN_5933; // @[Execute.scala 117:10]
  assign _GEN_5935 = 6'h2d == _T_544 ? welem[45] : _GEN_5934; // @[Execute.scala 117:10]
  assign _GEN_5936 = 6'h2e == _T_544 ? welem[46] : _GEN_5935; // @[Execute.scala 117:10]
  assign _GEN_5937 = 6'h2f == _T_544 ? welem[47] : _GEN_5936; // @[Execute.scala 117:10]
  assign _GEN_5938 = 6'h30 == _T_544 ? welem[48] : _GEN_5937; // @[Execute.scala 117:10]
  assign _GEN_5939 = 6'h31 == _T_544 ? welem[49] : _GEN_5938; // @[Execute.scala 117:10]
  assign _GEN_5940 = 6'h32 == _T_544 ? welem[50] : _GEN_5939; // @[Execute.scala 117:10]
  assign _GEN_5941 = 6'h33 == _T_544 ? welem[51] : _GEN_5940; // @[Execute.scala 117:10]
  assign _GEN_5942 = 6'h34 == _T_544 ? welem[52] : _GEN_5941; // @[Execute.scala 117:10]
  assign _GEN_5943 = 6'h35 == _T_544 ? welem[53] : _GEN_5942; // @[Execute.scala 117:10]
  assign _GEN_5944 = 6'h36 == _T_544 ? welem[54] : _GEN_5943; // @[Execute.scala 117:10]
  assign _GEN_5945 = 6'h37 == _T_544 ? welem[55] : _GEN_5944; // @[Execute.scala 117:10]
  assign _GEN_5946 = 6'h38 == _T_544 ? welem[56] : _GEN_5945; // @[Execute.scala 117:10]
  assign _GEN_5947 = 6'h39 == _T_544 ? welem[57] : _GEN_5946; // @[Execute.scala 117:10]
  assign _GEN_5948 = 6'h3a == _T_544 ? welem[58] : _GEN_5947; // @[Execute.scala 117:10]
  assign _GEN_5949 = 6'h3b == _T_544 ? welem[59] : _GEN_5948; // @[Execute.scala 117:10]
  assign _GEN_5950 = 6'h3c == _T_544 ? welem[60] : _GEN_5949; // @[Execute.scala 117:10]
  assign _GEN_5951 = 6'h3d == _T_544 ? welem[61] : _GEN_5950; // @[Execute.scala 117:10]
  assign _GEN_5952 = 6'h3e == _T_544 ? welem[62] : _GEN_5951; // @[Execute.scala 117:10]
  assign _GEN_5953 = 6'h3f == _T_544 ? welem[63] : _GEN_5952; // @[Execute.scala 117:10]
  assign _GEN_5955 = 6'h1 == _T_548 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_5956 = 6'h2 == _T_548 ? welem[2] : _GEN_5955; // @[Execute.scala 117:10]
  assign _GEN_5957 = 6'h3 == _T_548 ? welem[3] : _GEN_5956; // @[Execute.scala 117:10]
  assign _GEN_5958 = 6'h4 == _T_548 ? welem[4] : _GEN_5957; // @[Execute.scala 117:10]
  assign _GEN_5959 = 6'h5 == _T_548 ? welem[5] : _GEN_5958; // @[Execute.scala 117:10]
  assign _GEN_5960 = 6'h6 == _T_548 ? welem[6] : _GEN_5959; // @[Execute.scala 117:10]
  assign _GEN_5961 = 6'h7 == _T_548 ? welem[7] : _GEN_5960; // @[Execute.scala 117:10]
  assign _GEN_5962 = 6'h8 == _T_548 ? welem[8] : _GEN_5961; // @[Execute.scala 117:10]
  assign _GEN_5963 = 6'h9 == _T_548 ? welem[9] : _GEN_5962; // @[Execute.scala 117:10]
  assign _GEN_5964 = 6'ha == _T_548 ? welem[10] : _GEN_5963; // @[Execute.scala 117:10]
  assign _GEN_5965 = 6'hb == _T_548 ? welem[11] : _GEN_5964; // @[Execute.scala 117:10]
  assign _GEN_5966 = 6'hc == _T_548 ? welem[12] : _GEN_5965; // @[Execute.scala 117:10]
  assign _GEN_5967 = 6'hd == _T_548 ? welem[13] : _GEN_5966; // @[Execute.scala 117:10]
  assign _GEN_5968 = 6'he == _T_548 ? welem[14] : _GEN_5967; // @[Execute.scala 117:10]
  assign _GEN_5969 = 6'hf == _T_548 ? welem[15] : _GEN_5968; // @[Execute.scala 117:10]
  assign _GEN_5970 = 6'h10 == _T_548 ? welem[16] : _GEN_5969; // @[Execute.scala 117:10]
  assign _GEN_5971 = 6'h11 == _T_548 ? welem[17] : _GEN_5970; // @[Execute.scala 117:10]
  assign _GEN_5972 = 6'h12 == _T_548 ? welem[18] : _GEN_5971; // @[Execute.scala 117:10]
  assign _GEN_5973 = 6'h13 == _T_548 ? welem[19] : _GEN_5972; // @[Execute.scala 117:10]
  assign _GEN_5974 = 6'h14 == _T_548 ? welem[20] : _GEN_5973; // @[Execute.scala 117:10]
  assign _GEN_5975 = 6'h15 == _T_548 ? welem[21] : _GEN_5974; // @[Execute.scala 117:10]
  assign _GEN_5976 = 6'h16 == _T_548 ? welem[22] : _GEN_5975; // @[Execute.scala 117:10]
  assign _GEN_5977 = 6'h17 == _T_548 ? welem[23] : _GEN_5976; // @[Execute.scala 117:10]
  assign _GEN_5978 = 6'h18 == _T_548 ? welem[24] : _GEN_5977; // @[Execute.scala 117:10]
  assign _GEN_5979 = 6'h19 == _T_548 ? welem[25] : _GEN_5978; // @[Execute.scala 117:10]
  assign _GEN_5980 = 6'h1a == _T_548 ? welem[26] : _GEN_5979; // @[Execute.scala 117:10]
  assign _GEN_5981 = 6'h1b == _T_548 ? welem[27] : _GEN_5980; // @[Execute.scala 117:10]
  assign _GEN_5982 = 6'h1c == _T_548 ? welem[28] : _GEN_5981; // @[Execute.scala 117:10]
  assign _GEN_5983 = 6'h1d == _T_548 ? welem[29] : _GEN_5982; // @[Execute.scala 117:10]
  assign _GEN_5984 = 6'h1e == _T_548 ? welem[30] : _GEN_5983; // @[Execute.scala 117:10]
  assign _GEN_5985 = 6'h1f == _T_548 ? welem[31] : _GEN_5984; // @[Execute.scala 117:10]
  assign _GEN_5986 = 6'h20 == _T_548 ? welem[32] : _GEN_5985; // @[Execute.scala 117:10]
  assign _GEN_5987 = 6'h21 == _T_548 ? welem[33] : _GEN_5986; // @[Execute.scala 117:10]
  assign _GEN_5988 = 6'h22 == _T_548 ? welem[34] : _GEN_5987; // @[Execute.scala 117:10]
  assign _GEN_5989 = 6'h23 == _T_548 ? welem[35] : _GEN_5988; // @[Execute.scala 117:10]
  assign _GEN_5990 = 6'h24 == _T_548 ? welem[36] : _GEN_5989; // @[Execute.scala 117:10]
  assign _GEN_5991 = 6'h25 == _T_548 ? welem[37] : _GEN_5990; // @[Execute.scala 117:10]
  assign _GEN_5992 = 6'h26 == _T_548 ? welem[38] : _GEN_5991; // @[Execute.scala 117:10]
  assign _GEN_5993 = 6'h27 == _T_548 ? welem[39] : _GEN_5992; // @[Execute.scala 117:10]
  assign _GEN_5994 = 6'h28 == _T_548 ? welem[40] : _GEN_5993; // @[Execute.scala 117:10]
  assign _GEN_5995 = 6'h29 == _T_548 ? welem[41] : _GEN_5994; // @[Execute.scala 117:10]
  assign _GEN_5996 = 6'h2a == _T_548 ? welem[42] : _GEN_5995; // @[Execute.scala 117:10]
  assign _GEN_5997 = 6'h2b == _T_548 ? welem[43] : _GEN_5996; // @[Execute.scala 117:10]
  assign _GEN_5998 = 6'h2c == _T_548 ? welem[44] : _GEN_5997; // @[Execute.scala 117:10]
  assign _GEN_5999 = 6'h2d == _T_548 ? welem[45] : _GEN_5998; // @[Execute.scala 117:10]
  assign _GEN_6000 = 6'h2e == _T_548 ? welem[46] : _GEN_5999; // @[Execute.scala 117:10]
  assign _GEN_6001 = 6'h2f == _T_548 ? welem[47] : _GEN_6000; // @[Execute.scala 117:10]
  assign _GEN_6002 = 6'h30 == _T_548 ? welem[48] : _GEN_6001; // @[Execute.scala 117:10]
  assign _GEN_6003 = 6'h31 == _T_548 ? welem[49] : _GEN_6002; // @[Execute.scala 117:10]
  assign _GEN_6004 = 6'h32 == _T_548 ? welem[50] : _GEN_6003; // @[Execute.scala 117:10]
  assign _GEN_6005 = 6'h33 == _T_548 ? welem[51] : _GEN_6004; // @[Execute.scala 117:10]
  assign _GEN_6006 = 6'h34 == _T_548 ? welem[52] : _GEN_6005; // @[Execute.scala 117:10]
  assign _GEN_6007 = 6'h35 == _T_548 ? welem[53] : _GEN_6006; // @[Execute.scala 117:10]
  assign _GEN_6008 = 6'h36 == _T_548 ? welem[54] : _GEN_6007; // @[Execute.scala 117:10]
  assign _GEN_6009 = 6'h37 == _T_548 ? welem[55] : _GEN_6008; // @[Execute.scala 117:10]
  assign _GEN_6010 = 6'h38 == _T_548 ? welem[56] : _GEN_6009; // @[Execute.scala 117:10]
  assign _GEN_6011 = 6'h39 == _T_548 ? welem[57] : _GEN_6010; // @[Execute.scala 117:10]
  assign _GEN_6012 = 6'h3a == _T_548 ? welem[58] : _GEN_6011; // @[Execute.scala 117:10]
  assign _GEN_6013 = 6'h3b == _T_548 ? welem[59] : _GEN_6012; // @[Execute.scala 117:10]
  assign _GEN_6014 = 6'h3c == _T_548 ? welem[60] : _GEN_6013; // @[Execute.scala 117:10]
  assign _GEN_6015 = 6'h3d == _T_548 ? welem[61] : _GEN_6014; // @[Execute.scala 117:10]
  assign _GEN_6016 = 6'h3e == _T_548 ? welem[62] : _GEN_6015; // @[Execute.scala 117:10]
  assign _GEN_6017 = 6'h3f == _T_548 ? welem[63] : _GEN_6016; // @[Execute.scala 117:10]
  assign _T_551 = _T_542 ? _GEN_5953 : _GEN_6017; // @[Execute.scala 117:10]
  assign _T_552 = r < 6'h12; // @[Execute.scala 117:15]
  assign _T_554 = r - 6'h12; // @[Execute.scala 117:37]
  assign _T_558 = 6'h2e + r; // @[Execute.scala 117:60]
  assign _GEN_6019 = 6'h1 == _T_554 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6020 = 6'h2 == _T_554 ? welem[2] : _GEN_6019; // @[Execute.scala 117:10]
  assign _GEN_6021 = 6'h3 == _T_554 ? welem[3] : _GEN_6020; // @[Execute.scala 117:10]
  assign _GEN_6022 = 6'h4 == _T_554 ? welem[4] : _GEN_6021; // @[Execute.scala 117:10]
  assign _GEN_6023 = 6'h5 == _T_554 ? welem[5] : _GEN_6022; // @[Execute.scala 117:10]
  assign _GEN_6024 = 6'h6 == _T_554 ? welem[6] : _GEN_6023; // @[Execute.scala 117:10]
  assign _GEN_6025 = 6'h7 == _T_554 ? welem[7] : _GEN_6024; // @[Execute.scala 117:10]
  assign _GEN_6026 = 6'h8 == _T_554 ? welem[8] : _GEN_6025; // @[Execute.scala 117:10]
  assign _GEN_6027 = 6'h9 == _T_554 ? welem[9] : _GEN_6026; // @[Execute.scala 117:10]
  assign _GEN_6028 = 6'ha == _T_554 ? welem[10] : _GEN_6027; // @[Execute.scala 117:10]
  assign _GEN_6029 = 6'hb == _T_554 ? welem[11] : _GEN_6028; // @[Execute.scala 117:10]
  assign _GEN_6030 = 6'hc == _T_554 ? welem[12] : _GEN_6029; // @[Execute.scala 117:10]
  assign _GEN_6031 = 6'hd == _T_554 ? welem[13] : _GEN_6030; // @[Execute.scala 117:10]
  assign _GEN_6032 = 6'he == _T_554 ? welem[14] : _GEN_6031; // @[Execute.scala 117:10]
  assign _GEN_6033 = 6'hf == _T_554 ? welem[15] : _GEN_6032; // @[Execute.scala 117:10]
  assign _GEN_6034 = 6'h10 == _T_554 ? welem[16] : _GEN_6033; // @[Execute.scala 117:10]
  assign _GEN_6035 = 6'h11 == _T_554 ? welem[17] : _GEN_6034; // @[Execute.scala 117:10]
  assign _GEN_6036 = 6'h12 == _T_554 ? welem[18] : _GEN_6035; // @[Execute.scala 117:10]
  assign _GEN_6037 = 6'h13 == _T_554 ? welem[19] : _GEN_6036; // @[Execute.scala 117:10]
  assign _GEN_6038 = 6'h14 == _T_554 ? welem[20] : _GEN_6037; // @[Execute.scala 117:10]
  assign _GEN_6039 = 6'h15 == _T_554 ? welem[21] : _GEN_6038; // @[Execute.scala 117:10]
  assign _GEN_6040 = 6'h16 == _T_554 ? welem[22] : _GEN_6039; // @[Execute.scala 117:10]
  assign _GEN_6041 = 6'h17 == _T_554 ? welem[23] : _GEN_6040; // @[Execute.scala 117:10]
  assign _GEN_6042 = 6'h18 == _T_554 ? welem[24] : _GEN_6041; // @[Execute.scala 117:10]
  assign _GEN_6043 = 6'h19 == _T_554 ? welem[25] : _GEN_6042; // @[Execute.scala 117:10]
  assign _GEN_6044 = 6'h1a == _T_554 ? welem[26] : _GEN_6043; // @[Execute.scala 117:10]
  assign _GEN_6045 = 6'h1b == _T_554 ? welem[27] : _GEN_6044; // @[Execute.scala 117:10]
  assign _GEN_6046 = 6'h1c == _T_554 ? welem[28] : _GEN_6045; // @[Execute.scala 117:10]
  assign _GEN_6047 = 6'h1d == _T_554 ? welem[29] : _GEN_6046; // @[Execute.scala 117:10]
  assign _GEN_6048 = 6'h1e == _T_554 ? welem[30] : _GEN_6047; // @[Execute.scala 117:10]
  assign _GEN_6049 = 6'h1f == _T_554 ? welem[31] : _GEN_6048; // @[Execute.scala 117:10]
  assign _GEN_6050 = 6'h20 == _T_554 ? welem[32] : _GEN_6049; // @[Execute.scala 117:10]
  assign _GEN_6051 = 6'h21 == _T_554 ? welem[33] : _GEN_6050; // @[Execute.scala 117:10]
  assign _GEN_6052 = 6'h22 == _T_554 ? welem[34] : _GEN_6051; // @[Execute.scala 117:10]
  assign _GEN_6053 = 6'h23 == _T_554 ? welem[35] : _GEN_6052; // @[Execute.scala 117:10]
  assign _GEN_6054 = 6'h24 == _T_554 ? welem[36] : _GEN_6053; // @[Execute.scala 117:10]
  assign _GEN_6055 = 6'h25 == _T_554 ? welem[37] : _GEN_6054; // @[Execute.scala 117:10]
  assign _GEN_6056 = 6'h26 == _T_554 ? welem[38] : _GEN_6055; // @[Execute.scala 117:10]
  assign _GEN_6057 = 6'h27 == _T_554 ? welem[39] : _GEN_6056; // @[Execute.scala 117:10]
  assign _GEN_6058 = 6'h28 == _T_554 ? welem[40] : _GEN_6057; // @[Execute.scala 117:10]
  assign _GEN_6059 = 6'h29 == _T_554 ? welem[41] : _GEN_6058; // @[Execute.scala 117:10]
  assign _GEN_6060 = 6'h2a == _T_554 ? welem[42] : _GEN_6059; // @[Execute.scala 117:10]
  assign _GEN_6061 = 6'h2b == _T_554 ? welem[43] : _GEN_6060; // @[Execute.scala 117:10]
  assign _GEN_6062 = 6'h2c == _T_554 ? welem[44] : _GEN_6061; // @[Execute.scala 117:10]
  assign _GEN_6063 = 6'h2d == _T_554 ? welem[45] : _GEN_6062; // @[Execute.scala 117:10]
  assign _GEN_6064 = 6'h2e == _T_554 ? welem[46] : _GEN_6063; // @[Execute.scala 117:10]
  assign _GEN_6065 = 6'h2f == _T_554 ? welem[47] : _GEN_6064; // @[Execute.scala 117:10]
  assign _GEN_6066 = 6'h30 == _T_554 ? welem[48] : _GEN_6065; // @[Execute.scala 117:10]
  assign _GEN_6067 = 6'h31 == _T_554 ? welem[49] : _GEN_6066; // @[Execute.scala 117:10]
  assign _GEN_6068 = 6'h32 == _T_554 ? welem[50] : _GEN_6067; // @[Execute.scala 117:10]
  assign _GEN_6069 = 6'h33 == _T_554 ? welem[51] : _GEN_6068; // @[Execute.scala 117:10]
  assign _GEN_6070 = 6'h34 == _T_554 ? welem[52] : _GEN_6069; // @[Execute.scala 117:10]
  assign _GEN_6071 = 6'h35 == _T_554 ? welem[53] : _GEN_6070; // @[Execute.scala 117:10]
  assign _GEN_6072 = 6'h36 == _T_554 ? welem[54] : _GEN_6071; // @[Execute.scala 117:10]
  assign _GEN_6073 = 6'h37 == _T_554 ? welem[55] : _GEN_6072; // @[Execute.scala 117:10]
  assign _GEN_6074 = 6'h38 == _T_554 ? welem[56] : _GEN_6073; // @[Execute.scala 117:10]
  assign _GEN_6075 = 6'h39 == _T_554 ? welem[57] : _GEN_6074; // @[Execute.scala 117:10]
  assign _GEN_6076 = 6'h3a == _T_554 ? welem[58] : _GEN_6075; // @[Execute.scala 117:10]
  assign _GEN_6077 = 6'h3b == _T_554 ? welem[59] : _GEN_6076; // @[Execute.scala 117:10]
  assign _GEN_6078 = 6'h3c == _T_554 ? welem[60] : _GEN_6077; // @[Execute.scala 117:10]
  assign _GEN_6079 = 6'h3d == _T_554 ? welem[61] : _GEN_6078; // @[Execute.scala 117:10]
  assign _GEN_6080 = 6'h3e == _T_554 ? welem[62] : _GEN_6079; // @[Execute.scala 117:10]
  assign _GEN_6081 = 6'h3f == _T_554 ? welem[63] : _GEN_6080; // @[Execute.scala 117:10]
  assign _GEN_6083 = 6'h1 == _T_558 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6084 = 6'h2 == _T_558 ? welem[2] : _GEN_6083; // @[Execute.scala 117:10]
  assign _GEN_6085 = 6'h3 == _T_558 ? welem[3] : _GEN_6084; // @[Execute.scala 117:10]
  assign _GEN_6086 = 6'h4 == _T_558 ? welem[4] : _GEN_6085; // @[Execute.scala 117:10]
  assign _GEN_6087 = 6'h5 == _T_558 ? welem[5] : _GEN_6086; // @[Execute.scala 117:10]
  assign _GEN_6088 = 6'h6 == _T_558 ? welem[6] : _GEN_6087; // @[Execute.scala 117:10]
  assign _GEN_6089 = 6'h7 == _T_558 ? welem[7] : _GEN_6088; // @[Execute.scala 117:10]
  assign _GEN_6090 = 6'h8 == _T_558 ? welem[8] : _GEN_6089; // @[Execute.scala 117:10]
  assign _GEN_6091 = 6'h9 == _T_558 ? welem[9] : _GEN_6090; // @[Execute.scala 117:10]
  assign _GEN_6092 = 6'ha == _T_558 ? welem[10] : _GEN_6091; // @[Execute.scala 117:10]
  assign _GEN_6093 = 6'hb == _T_558 ? welem[11] : _GEN_6092; // @[Execute.scala 117:10]
  assign _GEN_6094 = 6'hc == _T_558 ? welem[12] : _GEN_6093; // @[Execute.scala 117:10]
  assign _GEN_6095 = 6'hd == _T_558 ? welem[13] : _GEN_6094; // @[Execute.scala 117:10]
  assign _GEN_6096 = 6'he == _T_558 ? welem[14] : _GEN_6095; // @[Execute.scala 117:10]
  assign _GEN_6097 = 6'hf == _T_558 ? welem[15] : _GEN_6096; // @[Execute.scala 117:10]
  assign _GEN_6098 = 6'h10 == _T_558 ? welem[16] : _GEN_6097; // @[Execute.scala 117:10]
  assign _GEN_6099 = 6'h11 == _T_558 ? welem[17] : _GEN_6098; // @[Execute.scala 117:10]
  assign _GEN_6100 = 6'h12 == _T_558 ? welem[18] : _GEN_6099; // @[Execute.scala 117:10]
  assign _GEN_6101 = 6'h13 == _T_558 ? welem[19] : _GEN_6100; // @[Execute.scala 117:10]
  assign _GEN_6102 = 6'h14 == _T_558 ? welem[20] : _GEN_6101; // @[Execute.scala 117:10]
  assign _GEN_6103 = 6'h15 == _T_558 ? welem[21] : _GEN_6102; // @[Execute.scala 117:10]
  assign _GEN_6104 = 6'h16 == _T_558 ? welem[22] : _GEN_6103; // @[Execute.scala 117:10]
  assign _GEN_6105 = 6'h17 == _T_558 ? welem[23] : _GEN_6104; // @[Execute.scala 117:10]
  assign _GEN_6106 = 6'h18 == _T_558 ? welem[24] : _GEN_6105; // @[Execute.scala 117:10]
  assign _GEN_6107 = 6'h19 == _T_558 ? welem[25] : _GEN_6106; // @[Execute.scala 117:10]
  assign _GEN_6108 = 6'h1a == _T_558 ? welem[26] : _GEN_6107; // @[Execute.scala 117:10]
  assign _GEN_6109 = 6'h1b == _T_558 ? welem[27] : _GEN_6108; // @[Execute.scala 117:10]
  assign _GEN_6110 = 6'h1c == _T_558 ? welem[28] : _GEN_6109; // @[Execute.scala 117:10]
  assign _GEN_6111 = 6'h1d == _T_558 ? welem[29] : _GEN_6110; // @[Execute.scala 117:10]
  assign _GEN_6112 = 6'h1e == _T_558 ? welem[30] : _GEN_6111; // @[Execute.scala 117:10]
  assign _GEN_6113 = 6'h1f == _T_558 ? welem[31] : _GEN_6112; // @[Execute.scala 117:10]
  assign _GEN_6114 = 6'h20 == _T_558 ? welem[32] : _GEN_6113; // @[Execute.scala 117:10]
  assign _GEN_6115 = 6'h21 == _T_558 ? welem[33] : _GEN_6114; // @[Execute.scala 117:10]
  assign _GEN_6116 = 6'h22 == _T_558 ? welem[34] : _GEN_6115; // @[Execute.scala 117:10]
  assign _GEN_6117 = 6'h23 == _T_558 ? welem[35] : _GEN_6116; // @[Execute.scala 117:10]
  assign _GEN_6118 = 6'h24 == _T_558 ? welem[36] : _GEN_6117; // @[Execute.scala 117:10]
  assign _GEN_6119 = 6'h25 == _T_558 ? welem[37] : _GEN_6118; // @[Execute.scala 117:10]
  assign _GEN_6120 = 6'h26 == _T_558 ? welem[38] : _GEN_6119; // @[Execute.scala 117:10]
  assign _GEN_6121 = 6'h27 == _T_558 ? welem[39] : _GEN_6120; // @[Execute.scala 117:10]
  assign _GEN_6122 = 6'h28 == _T_558 ? welem[40] : _GEN_6121; // @[Execute.scala 117:10]
  assign _GEN_6123 = 6'h29 == _T_558 ? welem[41] : _GEN_6122; // @[Execute.scala 117:10]
  assign _GEN_6124 = 6'h2a == _T_558 ? welem[42] : _GEN_6123; // @[Execute.scala 117:10]
  assign _GEN_6125 = 6'h2b == _T_558 ? welem[43] : _GEN_6124; // @[Execute.scala 117:10]
  assign _GEN_6126 = 6'h2c == _T_558 ? welem[44] : _GEN_6125; // @[Execute.scala 117:10]
  assign _GEN_6127 = 6'h2d == _T_558 ? welem[45] : _GEN_6126; // @[Execute.scala 117:10]
  assign _GEN_6128 = 6'h2e == _T_558 ? welem[46] : _GEN_6127; // @[Execute.scala 117:10]
  assign _GEN_6129 = 6'h2f == _T_558 ? welem[47] : _GEN_6128; // @[Execute.scala 117:10]
  assign _GEN_6130 = 6'h30 == _T_558 ? welem[48] : _GEN_6129; // @[Execute.scala 117:10]
  assign _GEN_6131 = 6'h31 == _T_558 ? welem[49] : _GEN_6130; // @[Execute.scala 117:10]
  assign _GEN_6132 = 6'h32 == _T_558 ? welem[50] : _GEN_6131; // @[Execute.scala 117:10]
  assign _GEN_6133 = 6'h33 == _T_558 ? welem[51] : _GEN_6132; // @[Execute.scala 117:10]
  assign _GEN_6134 = 6'h34 == _T_558 ? welem[52] : _GEN_6133; // @[Execute.scala 117:10]
  assign _GEN_6135 = 6'h35 == _T_558 ? welem[53] : _GEN_6134; // @[Execute.scala 117:10]
  assign _GEN_6136 = 6'h36 == _T_558 ? welem[54] : _GEN_6135; // @[Execute.scala 117:10]
  assign _GEN_6137 = 6'h37 == _T_558 ? welem[55] : _GEN_6136; // @[Execute.scala 117:10]
  assign _GEN_6138 = 6'h38 == _T_558 ? welem[56] : _GEN_6137; // @[Execute.scala 117:10]
  assign _GEN_6139 = 6'h39 == _T_558 ? welem[57] : _GEN_6138; // @[Execute.scala 117:10]
  assign _GEN_6140 = 6'h3a == _T_558 ? welem[58] : _GEN_6139; // @[Execute.scala 117:10]
  assign _GEN_6141 = 6'h3b == _T_558 ? welem[59] : _GEN_6140; // @[Execute.scala 117:10]
  assign _GEN_6142 = 6'h3c == _T_558 ? welem[60] : _GEN_6141; // @[Execute.scala 117:10]
  assign _GEN_6143 = 6'h3d == _T_558 ? welem[61] : _GEN_6142; // @[Execute.scala 117:10]
  assign _GEN_6144 = 6'h3e == _T_558 ? welem[62] : _GEN_6143; // @[Execute.scala 117:10]
  assign _GEN_6145 = 6'h3f == _T_558 ? welem[63] : _GEN_6144; // @[Execute.scala 117:10]
  assign _T_561 = _T_552 ? _GEN_6081 : _GEN_6145; // @[Execute.scala 117:10]
  assign _T_562 = r < 6'h11; // @[Execute.scala 117:15]
  assign _T_564 = r - 6'h11; // @[Execute.scala 117:37]
  assign _T_568 = 6'h2f + r; // @[Execute.scala 117:60]
  assign _GEN_6147 = 6'h1 == _T_564 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6148 = 6'h2 == _T_564 ? welem[2] : _GEN_6147; // @[Execute.scala 117:10]
  assign _GEN_6149 = 6'h3 == _T_564 ? welem[3] : _GEN_6148; // @[Execute.scala 117:10]
  assign _GEN_6150 = 6'h4 == _T_564 ? welem[4] : _GEN_6149; // @[Execute.scala 117:10]
  assign _GEN_6151 = 6'h5 == _T_564 ? welem[5] : _GEN_6150; // @[Execute.scala 117:10]
  assign _GEN_6152 = 6'h6 == _T_564 ? welem[6] : _GEN_6151; // @[Execute.scala 117:10]
  assign _GEN_6153 = 6'h7 == _T_564 ? welem[7] : _GEN_6152; // @[Execute.scala 117:10]
  assign _GEN_6154 = 6'h8 == _T_564 ? welem[8] : _GEN_6153; // @[Execute.scala 117:10]
  assign _GEN_6155 = 6'h9 == _T_564 ? welem[9] : _GEN_6154; // @[Execute.scala 117:10]
  assign _GEN_6156 = 6'ha == _T_564 ? welem[10] : _GEN_6155; // @[Execute.scala 117:10]
  assign _GEN_6157 = 6'hb == _T_564 ? welem[11] : _GEN_6156; // @[Execute.scala 117:10]
  assign _GEN_6158 = 6'hc == _T_564 ? welem[12] : _GEN_6157; // @[Execute.scala 117:10]
  assign _GEN_6159 = 6'hd == _T_564 ? welem[13] : _GEN_6158; // @[Execute.scala 117:10]
  assign _GEN_6160 = 6'he == _T_564 ? welem[14] : _GEN_6159; // @[Execute.scala 117:10]
  assign _GEN_6161 = 6'hf == _T_564 ? welem[15] : _GEN_6160; // @[Execute.scala 117:10]
  assign _GEN_6162 = 6'h10 == _T_564 ? welem[16] : _GEN_6161; // @[Execute.scala 117:10]
  assign _GEN_6163 = 6'h11 == _T_564 ? welem[17] : _GEN_6162; // @[Execute.scala 117:10]
  assign _GEN_6164 = 6'h12 == _T_564 ? welem[18] : _GEN_6163; // @[Execute.scala 117:10]
  assign _GEN_6165 = 6'h13 == _T_564 ? welem[19] : _GEN_6164; // @[Execute.scala 117:10]
  assign _GEN_6166 = 6'h14 == _T_564 ? welem[20] : _GEN_6165; // @[Execute.scala 117:10]
  assign _GEN_6167 = 6'h15 == _T_564 ? welem[21] : _GEN_6166; // @[Execute.scala 117:10]
  assign _GEN_6168 = 6'h16 == _T_564 ? welem[22] : _GEN_6167; // @[Execute.scala 117:10]
  assign _GEN_6169 = 6'h17 == _T_564 ? welem[23] : _GEN_6168; // @[Execute.scala 117:10]
  assign _GEN_6170 = 6'h18 == _T_564 ? welem[24] : _GEN_6169; // @[Execute.scala 117:10]
  assign _GEN_6171 = 6'h19 == _T_564 ? welem[25] : _GEN_6170; // @[Execute.scala 117:10]
  assign _GEN_6172 = 6'h1a == _T_564 ? welem[26] : _GEN_6171; // @[Execute.scala 117:10]
  assign _GEN_6173 = 6'h1b == _T_564 ? welem[27] : _GEN_6172; // @[Execute.scala 117:10]
  assign _GEN_6174 = 6'h1c == _T_564 ? welem[28] : _GEN_6173; // @[Execute.scala 117:10]
  assign _GEN_6175 = 6'h1d == _T_564 ? welem[29] : _GEN_6174; // @[Execute.scala 117:10]
  assign _GEN_6176 = 6'h1e == _T_564 ? welem[30] : _GEN_6175; // @[Execute.scala 117:10]
  assign _GEN_6177 = 6'h1f == _T_564 ? welem[31] : _GEN_6176; // @[Execute.scala 117:10]
  assign _GEN_6178 = 6'h20 == _T_564 ? welem[32] : _GEN_6177; // @[Execute.scala 117:10]
  assign _GEN_6179 = 6'h21 == _T_564 ? welem[33] : _GEN_6178; // @[Execute.scala 117:10]
  assign _GEN_6180 = 6'h22 == _T_564 ? welem[34] : _GEN_6179; // @[Execute.scala 117:10]
  assign _GEN_6181 = 6'h23 == _T_564 ? welem[35] : _GEN_6180; // @[Execute.scala 117:10]
  assign _GEN_6182 = 6'h24 == _T_564 ? welem[36] : _GEN_6181; // @[Execute.scala 117:10]
  assign _GEN_6183 = 6'h25 == _T_564 ? welem[37] : _GEN_6182; // @[Execute.scala 117:10]
  assign _GEN_6184 = 6'h26 == _T_564 ? welem[38] : _GEN_6183; // @[Execute.scala 117:10]
  assign _GEN_6185 = 6'h27 == _T_564 ? welem[39] : _GEN_6184; // @[Execute.scala 117:10]
  assign _GEN_6186 = 6'h28 == _T_564 ? welem[40] : _GEN_6185; // @[Execute.scala 117:10]
  assign _GEN_6187 = 6'h29 == _T_564 ? welem[41] : _GEN_6186; // @[Execute.scala 117:10]
  assign _GEN_6188 = 6'h2a == _T_564 ? welem[42] : _GEN_6187; // @[Execute.scala 117:10]
  assign _GEN_6189 = 6'h2b == _T_564 ? welem[43] : _GEN_6188; // @[Execute.scala 117:10]
  assign _GEN_6190 = 6'h2c == _T_564 ? welem[44] : _GEN_6189; // @[Execute.scala 117:10]
  assign _GEN_6191 = 6'h2d == _T_564 ? welem[45] : _GEN_6190; // @[Execute.scala 117:10]
  assign _GEN_6192 = 6'h2e == _T_564 ? welem[46] : _GEN_6191; // @[Execute.scala 117:10]
  assign _GEN_6193 = 6'h2f == _T_564 ? welem[47] : _GEN_6192; // @[Execute.scala 117:10]
  assign _GEN_6194 = 6'h30 == _T_564 ? welem[48] : _GEN_6193; // @[Execute.scala 117:10]
  assign _GEN_6195 = 6'h31 == _T_564 ? welem[49] : _GEN_6194; // @[Execute.scala 117:10]
  assign _GEN_6196 = 6'h32 == _T_564 ? welem[50] : _GEN_6195; // @[Execute.scala 117:10]
  assign _GEN_6197 = 6'h33 == _T_564 ? welem[51] : _GEN_6196; // @[Execute.scala 117:10]
  assign _GEN_6198 = 6'h34 == _T_564 ? welem[52] : _GEN_6197; // @[Execute.scala 117:10]
  assign _GEN_6199 = 6'h35 == _T_564 ? welem[53] : _GEN_6198; // @[Execute.scala 117:10]
  assign _GEN_6200 = 6'h36 == _T_564 ? welem[54] : _GEN_6199; // @[Execute.scala 117:10]
  assign _GEN_6201 = 6'h37 == _T_564 ? welem[55] : _GEN_6200; // @[Execute.scala 117:10]
  assign _GEN_6202 = 6'h38 == _T_564 ? welem[56] : _GEN_6201; // @[Execute.scala 117:10]
  assign _GEN_6203 = 6'h39 == _T_564 ? welem[57] : _GEN_6202; // @[Execute.scala 117:10]
  assign _GEN_6204 = 6'h3a == _T_564 ? welem[58] : _GEN_6203; // @[Execute.scala 117:10]
  assign _GEN_6205 = 6'h3b == _T_564 ? welem[59] : _GEN_6204; // @[Execute.scala 117:10]
  assign _GEN_6206 = 6'h3c == _T_564 ? welem[60] : _GEN_6205; // @[Execute.scala 117:10]
  assign _GEN_6207 = 6'h3d == _T_564 ? welem[61] : _GEN_6206; // @[Execute.scala 117:10]
  assign _GEN_6208 = 6'h3e == _T_564 ? welem[62] : _GEN_6207; // @[Execute.scala 117:10]
  assign _GEN_6209 = 6'h3f == _T_564 ? welem[63] : _GEN_6208; // @[Execute.scala 117:10]
  assign _GEN_6211 = 6'h1 == _T_568 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6212 = 6'h2 == _T_568 ? welem[2] : _GEN_6211; // @[Execute.scala 117:10]
  assign _GEN_6213 = 6'h3 == _T_568 ? welem[3] : _GEN_6212; // @[Execute.scala 117:10]
  assign _GEN_6214 = 6'h4 == _T_568 ? welem[4] : _GEN_6213; // @[Execute.scala 117:10]
  assign _GEN_6215 = 6'h5 == _T_568 ? welem[5] : _GEN_6214; // @[Execute.scala 117:10]
  assign _GEN_6216 = 6'h6 == _T_568 ? welem[6] : _GEN_6215; // @[Execute.scala 117:10]
  assign _GEN_6217 = 6'h7 == _T_568 ? welem[7] : _GEN_6216; // @[Execute.scala 117:10]
  assign _GEN_6218 = 6'h8 == _T_568 ? welem[8] : _GEN_6217; // @[Execute.scala 117:10]
  assign _GEN_6219 = 6'h9 == _T_568 ? welem[9] : _GEN_6218; // @[Execute.scala 117:10]
  assign _GEN_6220 = 6'ha == _T_568 ? welem[10] : _GEN_6219; // @[Execute.scala 117:10]
  assign _GEN_6221 = 6'hb == _T_568 ? welem[11] : _GEN_6220; // @[Execute.scala 117:10]
  assign _GEN_6222 = 6'hc == _T_568 ? welem[12] : _GEN_6221; // @[Execute.scala 117:10]
  assign _GEN_6223 = 6'hd == _T_568 ? welem[13] : _GEN_6222; // @[Execute.scala 117:10]
  assign _GEN_6224 = 6'he == _T_568 ? welem[14] : _GEN_6223; // @[Execute.scala 117:10]
  assign _GEN_6225 = 6'hf == _T_568 ? welem[15] : _GEN_6224; // @[Execute.scala 117:10]
  assign _GEN_6226 = 6'h10 == _T_568 ? welem[16] : _GEN_6225; // @[Execute.scala 117:10]
  assign _GEN_6227 = 6'h11 == _T_568 ? welem[17] : _GEN_6226; // @[Execute.scala 117:10]
  assign _GEN_6228 = 6'h12 == _T_568 ? welem[18] : _GEN_6227; // @[Execute.scala 117:10]
  assign _GEN_6229 = 6'h13 == _T_568 ? welem[19] : _GEN_6228; // @[Execute.scala 117:10]
  assign _GEN_6230 = 6'h14 == _T_568 ? welem[20] : _GEN_6229; // @[Execute.scala 117:10]
  assign _GEN_6231 = 6'h15 == _T_568 ? welem[21] : _GEN_6230; // @[Execute.scala 117:10]
  assign _GEN_6232 = 6'h16 == _T_568 ? welem[22] : _GEN_6231; // @[Execute.scala 117:10]
  assign _GEN_6233 = 6'h17 == _T_568 ? welem[23] : _GEN_6232; // @[Execute.scala 117:10]
  assign _GEN_6234 = 6'h18 == _T_568 ? welem[24] : _GEN_6233; // @[Execute.scala 117:10]
  assign _GEN_6235 = 6'h19 == _T_568 ? welem[25] : _GEN_6234; // @[Execute.scala 117:10]
  assign _GEN_6236 = 6'h1a == _T_568 ? welem[26] : _GEN_6235; // @[Execute.scala 117:10]
  assign _GEN_6237 = 6'h1b == _T_568 ? welem[27] : _GEN_6236; // @[Execute.scala 117:10]
  assign _GEN_6238 = 6'h1c == _T_568 ? welem[28] : _GEN_6237; // @[Execute.scala 117:10]
  assign _GEN_6239 = 6'h1d == _T_568 ? welem[29] : _GEN_6238; // @[Execute.scala 117:10]
  assign _GEN_6240 = 6'h1e == _T_568 ? welem[30] : _GEN_6239; // @[Execute.scala 117:10]
  assign _GEN_6241 = 6'h1f == _T_568 ? welem[31] : _GEN_6240; // @[Execute.scala 117:10]
  assign _GEN_6242 = 6'h20 == _T_568 ? welem[32] : _GEN_6241; // @[Execute.scala 117:10]
  assign _GEN_6243 = 6'h21 == _T_568 ? welem[33] : _GEN_6242; // @[Execute.scala 117:10]
  assign _GEN_6244 = 6'h22 == _T_568 ? welem[34] : _GEN_6243; // @[Execute.scala 117:10]
  assign _GEN_6245 = 6'h23 == _T_568 ? welem[35] : _GEN_6244; // @[Execute.scala 117:10]
  assign _GEN_6246 = 6'h24 == _T_568 ? welem[36] : _GEN_6245; // @[Execute.scala 117:10]
  assign _GEN_6247 = 6'h25 == _T_568 ? welem[37] : _GEN_6246; // @[Execute.scala 117:10]
  assign _GEN_6248 = 6'h26 == _T_568 ? welem[38] : _GEN_6247; // @[Execute.scala 117:10]
  assign _GEN_6249 = 6'h27 == _T_568 ? welem[39] : _GEN_6248; // @[Execute.scala 117:10]
  assign _GEN_6250 = 6'h28 == _T_568 ? welem[40] : _GEN_6249; // @[Execute.scala 117:10]
  assign _GEN_6251 = 6'h29 == _T_568 ? welem[41] : _GEN_6250; // @[Execute.scala 117:10]
  assign _GEN_6252 = 6'h2a == _T_568 ? welem[42] : _GEN_6251; // @[Execute.scala 117:10]
  assign _GEN_6253 = 6'h2b == _T_568 ? welem[43] : _GEN_6252; // @[Execute.scala 117:10]
  assign _GEN_6254 = 6'h2c == _T_568 ? welem[44] : _GEN_6253; // @[Execute.scala 117:10]
  assign _GEN_6255 = 6'h2d == _T_568 ? welem[45] : _GEN_6254; // @[Execute.scala 117:10]
  assign _GEN_6256 = 6'h2e == _T_568 ? welem[46] : _GEN_6255; // @[Execute.scala 117:10]
  assign _GEN_6257 = 6'h2f == _T_568 ? welem[47] : _GEN_6256; // @[Execute.scala 117:10]
  assign _GEN_6258 = 6'h30 == _T_568 ? welem[48] : _GEN_6257; // @[Execute.scala 117:10]
  assign _GEN_6259 = 6'h31 == _T_568 ? welem[49] : _GEN_6258; // @[Execute.scala 117:10]
  assign _GEN_6260 = 6'h32 == _T_568 ? welem[50] : _GEN_6259; // @[Execute.scala 117:10]
  assign _GEN_6261 = 6'h33 == _T_568 ? welem[51] : _GEN_6260; // @[Execute.scala 117:10]
  assign _GEN_6262 = 6'h34 == _T_568 ? welem[52] : _GEN_6261; // @[Execute.scala 117:10]
  assign _GEN_6263 = 6'h35 == _T_568 ? welem[53] : _GEN_6262; // @[Execute.scala 117:10]
  assign _GEN_6264 = 6'h36 == _T_568 ? welem[54] : _GEN_6263; // @[Execute.scala 117:10]
  assign _GEN_6265 = 6'h37 == _T_568 ? welem[55] : _GEN_6264; // @[Execute.scala 117:10]
  assign _GEN_6266 = 6'h38 == _T_568 ? welem[56] : _GEN_6265; // @[Execute.scala 117:10]
  assign _GEN_6267 = 6'h39 == _T_568 ? welem[57] : _GEN_6266; // @[Execute.scala 117:10]
  assign _GEN_6268 = 6'h3a == _T_568 ? welem[58] : _GEN_6267; // @[Execute.scala 117:10]
  assign _GEN_6269 = 6'h3b == _T_568 ? welem[59] : _GEN_6268; // @[Execute.scala 117:10]
  assign _GEN_6270 = 6'h3c == _T_568 ? welem[60] : _GEN_6269; // @[Execute.scala 117:10]
  assign _GEN_6271 = 6'h3d == _T_568 ? welem[61] : _GEN_6270; // @[Execute.scala 117:10]
  assign _GEN_6272 = 6'h3e == _T_568 ? welem[62] : _GEN_6271; // @[Execute.scala 117:10]
  assign _GEN_6273 = 6'h3f == _T_568 ? welem[63] : _GEN_6272; // @[Execute.scala 117:10]
  assign _T_571 = _T_562 ? _GEN_6209 : _GEN_6273; // @[Execute.scala 117:10]
  assign _T_572 = r < 6'h10; // @[Execute.scala 117:15]
  assign _T_574 = r - 6'h10; // @[Execute.scala 117:37]
  assign _T_578 = 6'h30 + r; // @[Execute.scala 117:60]
  assign _GEN_6275 = 6'h1 == _T_574 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6276 = 6'h2 == _T_574 ? welem[2] : _GEN_6275; // @[Execute.scala 117:10]
  assign _GEN_6277 = 6'h3 == _T_574 ? welem[3] : _GEN_6276; // @[Execute.scala 117:10]
  assign _GEN_6278 = 6'h4 == _T_574 ? welem[4] : _GEN_6277; // @[Execute.scala 117:10]
  assign _GEN_6279 = 6'h5 == _T_574 ? welem[5] : _GEN_6278; // @[Execute.scala 117:10]
  assign _GEN_6280 = 6'h6 == _T_574 ? welem[6] : _GEN_6279; // @[Execute.scala 117:10]
  assign _GEN_6281 = 6'h7 == _T_574 ? welem[7] : _GEN_6280; // @[Execute.scala 117:10]
  assign _GEN_6282 = 6'h8 == _T_574 ? welem[8] : _GEN_6281; // @[Execute.scala 117:10]
  assign _GEN_6283 = 6'h9 == _T_574 ? welem[9] : _GEN_6282; // @[Execute.scala 117:10]
  assign _GEN_6284 = 6'ha == _T_574 ? welem[10] : _GEN_6283; // @[Execute.scala 117:10]
  assign _GEN_6285 = 6'hb == _T_574 ? welem[11] : _GEN_6284; // @[Execute.scala 117:10]
  assign _GEN_6286 = 6'hc == _T_574 ? welem[12] : _GEN_6285; // @[Execute.scala 117:10]
  assign _GEN_6287 = 6'hd == _T_574 ? welem[13] : _GEN_6286; // @[Execute.scala 117:10]
  assign _GEN_6288 = 6'he == _T_574 ? welem[14] : _GEN_6287; // @[Execute.scala 117:10]
  assign _GEN_6289 = 6'hf == _T_574 ? welem[15] : _GEN_6288; // @[Execute.scala 117:10]
  assign _GEN_6290 = 6'h10 == _T_574 ? welem[16] : _GEN_6289; // @[Execute.scala 117:10]
  assign _GEN_6291 = 6'h11 == _T_574 ? welem[17] : _GEN_6290; // @[Execute.scala 117:10]
  assign _GEN_6292 = 6'h12 == _T_574 ? welem[18] : _GEN_6291; // @[Execute.scala 117:10]
  assign _GEN_6293 = 6'h13 == _T_574 ? welem[19] : _GEN_6292; // @[Execute.scala 117:10]
  assign _GEN_6294 = 6'h14 == _T_574 ? welem[20] : _GEN_6293; // @[Execute.scala 117:10]
  assign _GEN_6295 = 6'h15 == _T_574 ? welem[21] : _GEN_6294; // @[Execute.scala 117:10]
  assign _GEN_6296 = 6'h16 == _T_574 ? welem[22] : _GEN_6295; // @[Execute.scala 117:10]
  assign _GEN_6297 = 6'h17 == _T_574 ? welem[23] : _GEN_6296; // @[Execute.scala 117:10]
  assign _GEN_6298 = 6'h18 == _T_574 ? welem[24] : _GEN_6297; // @[Execute.scala 117:10]
  assign _GEN_6299 = 6'h19 == _T_574 ? welem[25] : _GEN_6298; // @[Execute.scala 117:10]
  assign _GEN_6300 = 6'h1a == _T_574 ? welem[26] : _GEN_6299; // @[Execute.scala 117:10]
  assign _GEN_6301 = 6'h1b == _T_574 ? welem[27] : _GEN_6300; // @[Execute.scala 117:10]
  assign _GEN_6302 = 6'h1c == _T_574 ? welem[28] : _GEN_6301; // @[Execute.scala 117:10]
  assign _GEN_6303 = 6'h1d == _T_574 ? welem[29] : _GEN_6302; // @[Execute.scala 117:10]
  assign _GEN_6304 = 6'h1e == _T_574 ? welem[30] : _GEN_6303; // @[Execute.scala 117:10]
  assign _GEN_6305 = 6'h1f == _T_574 ? welem[31] : _GEN_6304; // @[Execute.scala 117:10]
  assign _GEN_6306 = 6'h20 == _T_574 ? welem[32] : _GEN_6305; // @[Execute.scala 117:10]
  assign _GEN_6307 = 6'h21 == _T_574 ? welem[33] : _GEN_6306; // @[Execute.scala 117:10]
  assign _GEN_6308 = 6'h22 == _T_574 ? welem[34] : _GEN_6307; // @[Execute.scala 117:10]
  assign _GEN_6309 = 6'h23 == _T_574 ? welem[35] : _GEN_6308; // @[Execute.scala 117:10]
  assign _GEN_6310 = 6'h24 == _T_574 ? welem[36] : _GEN_6309; // @[Execute.scala 117:10]
  assign _GEN_6311 = 6'h25 == _T_574 ? welem[37] : _GEN_6310; // @[Execute.scala 117:10]
  assign _GEN_6312 = 6'h26 == _T_574 ? welem[38] : _GEN_6311; // @[Execute.scala 117:10]
  assign _GEN_6313 = 6'h27 == _T_574 ? welem[39] : _GEN_6312; // @[Execute.scala 117:10]
  assign _GEN_6314 = 6'h28 == _T_574 ? welem[40] : _GEN_6313; // @[Execute.scala 117:10]
  assign _GEN_6315 = 6'h29 == _T_574 ? welem[41] : _GEN_6314; // @[Execute.scala 117:10]
  assign _GEN_6316 = 6'h2a == _T_574 ? welem[42] : _GEN_6315; // @[Execute.scala 117:10]
  assign _GEN_6317 = 6'h2b == _T_574 ? welem[43] : _GEN_6316; // @[Execute.scala 117:10]
  assign _GEN_6318 = 6'h2c == _T_574 ? welem[44] : _GEN_6317; // @[Execute.scala 117:10]
  assign _GEN_6319 = 6'h2d == _T_574 ? welem[45] : _GEN_6318; // @[Execute.scala 117:10]
  assign _GEN_6320 = 6'h2e == _T_574 ? welem[46] : _GEN_6319; // @[Execute.scala 117:10]
  assign _GEN_6321 = 6'h2f == _T_574 ? welem[47] : _GEN_6320; // @[Execute.scala 117:10]
  assign _GEN_6322 = 6'h30 == _T_574 ? welem[48] : _GEN_6321; // @[Execute.scala 117:10]
  assign _GEN_6323 = 6'h31 == _T_574 ? welem[49] : _GEN_6322; // @[Execute.scala 117:10]
  assign _GEN_6324 = 6'h32 == _T_574 ? welem[50] : _GEN_6323; // @[Execute.scala 117:10]
  assign _GEN_6325 = 6'h33 == _T_574 ? welem[51] : _GEN_6324; // @[Execute.scala 117:10]
  assign _GEN_6326 = 6'h34 == _T_574 ? welem[52] : _GEN_6325; // @[Execute.scala 117:10]
  assign _GEN_6327 = 6'h35 == _T_574 ? welem[53] : _GEN_6326; // @[Execute.scala 117:10]
  assign _GEN_6328 = 6'h36 == _T_574 ? welem[54] : _GEN_6327; // @[Execute.scala 117:10]
  assign _GEN_6329 = 6'h37 == _T_574 ? welem[55] : _GEN_6328; // @[Execute.scala 117:10]
  assign _GEN_6330 = 6'h38 == _T_574 ? welem[56] : _GEN_6329; // @[Execute.scala 117:10]
  assign _GEN_6331 = 6'h39 == _T_574 ? welem[57] : _GEN_6330; // @[Execute.scala 117:10]
  assign _GEN_6332 = 6'h3a == _T_574 ? welem[58] : _GEN_6331; // @[Execute.scala 117:10]
  assign _GEN_6333 = 6'h3b == _T_574 ? welem[59] : _GEN_6332; // @[Execute.scala 117:10]
  assign _GEN_6334 = 6'h3c == _T_574 ? welem[60] : _GEN_6333; // @[Execute.scala 117:10]
  assign _GEN_6335 = 6'h3d == _T_574 ? welem[61] : _GEN_6334; // @[Execute.scala 117:10]
  assign _GEN_6336 = 6'h3e == _T_574 ? welem[62] : _GEN_6335; // @[Execute.scala 117:10]
  assign _GEN_6337 = 6'h3f == _T_574 ? welem[63] : _GEN_6336; // @[Execute.scala 117:10]
  assign _GEN_6339 = 6'h1 == _T_578 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6340 = 6'h2 == _T_578 ? welem[2] : _GEN_6339; // @[Execute.scala 117:10]
  assign _GEN_6341 = 6'h3 == _T_578 ? welem[3] : _GEN_6340; // @[Execute.scala 117:10]
  assign _GEN_6342 = 6'h4 == _T_578 ? welem[4] : _GEN_6341; // @[Execute.scala 117:10]
  assign _GEN_6343 = 6'h5 == _T_578 ? welem[5] : _GEN_6342; // @[Execute.scala 117:10]
  assign _GEN_6344 = 6'h6 == _T_578 ? welem[6] : _GEN_6343; // @[Execute.scala 117:10]
  assign _GEN_6345 = 6'h7 == _T_578 ? welem[7] : _GEN_6344; // @[Execute.scala 117:10]
  assign _GEN_6346 = 6'h8 == _T_578 ? welem[8] : _GEN_6345; // @[Execute.scala 117:10]
  assign _GEN_6347 = 6'h9 == _T_578 ? welem[9] : _GEN_6346; // @[Execute.scala 117:10]
  assign _GEN_6348 = 6'ha == _T_578 ? welem[10] : _GEN_6347; // @[Execute.scala 117:10]
  assign _GEN_6349 = 6'hb == _T_578 ? welem[11] : _GEN_6348; // @[Execute.scala 117:10]
  assign _GEN_6350 = 6'hc == _T_578 ? welem[12] : _GEN_6349; // @[Execute.scala 117:10]
  assign _GEN_6351 = 6'hd == _T_578 ? welem[13] : _GEN_6350; // @[Execute.scala 117:10]
  assign _GEN_6352 = 6'he == _T_578 ? welem[14] : _GEN_6351; // @[Execute.scala 117:10]
  assign _GEN_6353 = 6'hf == _T_578 ? welem[15] : _GEN_6352; // @[Execute.scala 117:10]
  assign _GEN_6354 = 6'h10 == _T_578 ? welem[16] : _GEN_6353; // @[Execute.scala 117:10]
  assign _GEN_6355 = 6'h11 == _T_578 ? welem[17] : _GEN_6354; // @[Execute.scala 117:10]
  assign _GEN_6356 = 6'h12 == _T_578 ? welem[18] : _GEN_6355; // @[Execute.scala 117:10]
  assign _GEN_6357 = 6'h13 == _T_578 ? welem[19] : _GEN_6356; // @[Execute.scala 117:10]
  assign _GEN_6358 = 6'h14 == _T_578 ? welem[20] : _GEN_6357; // @[Execute.scala 117:10]
  assign _GEN_6359 = 6'h15 == _T_578 ? welem[21] : _GEN_6358; // @[Execute.scala 117:10]
  assign _GEN_6360 = 6'h16 == _T_578 ? welem[22] : _GEN_6359; // @[Execute.scala 117:10]
  assign _GEN_6361 = 6'h17 == _T_578 ? welem[23] : _GEN_6360; // @[Execute.scala 117:10]
  assign _GEN_6362 = 6'h18 == _T_578 ? welem[24] : _GEN_6361; // @[Execute.scala 117:10]
  assign _GEN_6363 = 6'h19 == _T_578 ? welem[25] : _GEN_6362; // @[Execute.scala 117:10]
  assign _GEN_6364 = 6'h1a == _T_578 ? welem[26] : _GEN_6363; // @[Execute.scala 117:10]
  assign _GEN_6365 = 6'h1b == _T_578 ? welem[27] : _GEN_6364; // @[Execute.scala 117:10]
  assign _GEN_6366 = 6'h1c == _T_578 ? welem[28] : _GEN_6365; // @[Execute.scala 117:10]
  assign _GEN_6367 = 6'h1d == _T_578 ? welem[29] : _GEN_6366; // @[Execute.scala 117:10]
  assign _GEN_6368 = 6'h1e == _T_578 ? welem[30] : _GEN_6367; // @[Execute.scala 117:10]
  assign _GEN_6369 = 6'h1f == _T_578 ? welem[31] : _GEN_6368; // @[Execute.scala 117:10]
  assign _GEN_6370 = 6'h20 == _T_578 ? welem[32] : _GEN_6369; // @[Execute.scala 117:10]
  assign _GEN_6371 = 6'h21 == _T_578 ? welem[33] : _GEN_6370; // @[Execute.scala 117:10]
  assign _GEN_6372 = 6'h22 == _T_578 ? welem[34] : _GEN_6371; // @[Execute.scala 117:10]
  assign _GEN_6373 = 6'h23 == _T_578 ? welem[35] : _GEN_6372; // @[Execute.scala 117:10]
  assign _GEN_6374 = 6'h24 == _T_578 ? welem[36] : _GEN_6373; // @[Execute.scala 117:10]
  assign _GEN_6375 = 6'h25 == _T_578 ? welem[37] : _GEN_6374; // @[Execute.scala 117:10]
  assign _GEN_6376 = 6'h26 == _T_578 ? welem[38] : _GEN_6375; // @[Execute.scala 117:10]
  assign _GEN_6377 = 6'h27 == _T_578 ? welem[39] : _GEN_6376; // @[Execute.scala 117:10]
  assign _GEN_6378 = 6'h28 == _T_578 ? welem[40] : _GEN_6377; // @[Execute.scala 117:10]
  assign _GEN_6379 = 6'h29 == _T_578 ? welem[41] : _GEN_6378; // @[Execute.scala 117:10]
  assign _GEN_6380 = 6'h2a == _T_578 ? welem[42] : _GEN_6379; // @[Execute.scala 117:10]
  assign _GEN_6381 = 6'h2b == _T_578 ? welem[43] : _GEN_6380; // @[Execute.scala 117:10]
  assign _GEN_6382 = 6'h2c == _T_578 ? welem[44] : _GEN_6381; // @[Execute.scala 117:10]
  assign _GEN_6383 = 6'h2d == _T_578 ? welem[45] : _GEN_6382; // @[Execute.scala 117:10]
  assign _GEN_6384 = 6'h2e == _T_578 ? welem[46] : _GEN_6383; // @[Execute.scala 117:10]
  assign _GEN_6385 = 6'h2f == _T_578 ? welem[47] : _GEN_6384; // @[Execute.scala 117:10]
  assign _GEN_6386 = 6'h30 == _T_578 ? welem[48] : _GEN_6385; // @[Execute.scala 117:10]
  assign _GEN_6387 = 6'h31 == _T_578 ? welem[49] : _GEN_6386; // @[Execute.scala 117:10]
  assign _GEN_6388 = 6'h32 == _T_578 ? welem[50] : _GEN_6387; // @[Execute.scala 117:10]
  assign _GEN_6389 = 6'h33 == _T_578 ? welem[51] : _GEN_6388; // @[Execute.scala 117:10]
  assign _GEN_6390 = 6'h34 == _T_578 ? welem[52] : _GEN_6389; // @[Execute.scala 117:10]
  assign _GEN_6391 = 6'h35 == _T_578 ? welem[53] : _GEN_6390; // @[Execute.scala 117:10]
  assign _GEN_6392 = 6'h36 == _T_578 ? welem[54] : _GEN_6391; // @[Execute.scala 117:10]
  assign _GEN_6393 = 6'h37 == _T_578 ? welem[55] : _GEN_6392; // @[Execute.scala 117:10]
  assign _GEN_6394 = 6'h38 == _T_578 ? welem[56] : _GEN_6393; // @[Execute.scala 117:10]
  assign _GEN_6395 = 6'h39 == _T_578 ? welem[57] : _GEN_6394; // @[Execute.scala 117:10]
  assign _GEN_6396 = 6'h3a == _T_578 ? welem[58] : _GEN_6395; // @[Execute.scala 117:10]
  assign _GEN_6397 = 6'h3b == _T_578 ? welem[59] : _GEN_6396; // @[Execute.scala 117:10]
  assign _GEN_6398 = 6'h3c == _T_578 ? welem[60] : _GEN_6397; // @[Execute.scala 117:10]
  assign _GEN_6399 = 6'h3d == _T_578 ? welem[61] : _GEN_6398; // @[Execute.scala 117:10]
  assign _GEN_6400 = 6'h3e == _T_578 ? welem[62] : _GEN_6399; // @[Execute.scala 117:10]
  assign _GEN_6401 = 6'h3f == _T_578 ? welem[63] : _GEN_6400; // @[Execute.scala 117:10]
  assign _T_581 = _T_572 ? _GEN_6337 : _GEN_6401; // @[Execute.scala 117:10]
  assign _T_582 = r < 6'hf; // @[Execute.scala 117:15]
  assign _T_584 = r - 6'hf; // @[Execute.scala 117:37]
  assign _T_588 = 6'h31 + r; // @[Execute.scala 117:60]
  assign _GEN_6403 = 6'h1 == _T_584 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6404 = 6'h2 == _T_584 ? welem[2] : _GEN_6403; // @[Execute.scala 117:10]
  assign _GEN_6405 = 6'h3 == _T_584 ? welem[3] : _GEN_6404; // @[Execute.scala 117:10]
  assign _GEN_6406 = 6'h4 == _T_584 ? welem[4] : _GEN_6405; // @[Execute.scala 117:10]
  assign _GEN_6407 = 6'h5 == _T_584 ? welem[5] : _GEN_6406; // @[Execute.scala 117:10]
  assign _GEN_6408 = 6'h6 == _T_584 ? welem[6] : _GEN_6407; // @[Execute.scala 117:10]
  assign _GEN_6409 = 6'h7 == _T_584 ? welem[7] : _GEN_6408; // @[Execute.scala 117:10]
  assign _GEN_6410 = 6'h8 == _T_584 ? welem[8] : _GEN_6409; // @[Execute.scala 117:10]
  assign _GEN_6411 = 6'h9 == _T_584 ? welem[9] : _GEN_6410; // @[Execute.scala 117:10]
  assign _GEN_6412 = 6'ha == _T_584 ? welem[10] : _GEN_6411; // @[Execute.scala 117:10]
  assign _GEN_6413 = 6'hb == _T_584 ? welem[11] : _GEN_6412; // @[Execute.scala 117:10]
  assign _GEN_6414 = 6'hc == _T_584 ? welem[12] : _GEN_6413; // @[Execute.scala 117:10]
  assign _GEN_6415 = 6'hd == _T_584 ? welem[13] : _GEN_6414; // @[Execute.scala 117:10]
  assign _GEN_6416 = 6'he == _T_584 ? welem[14] : _GEN_6415; // @[Execute.scala 117:10]
  assign _GEN_6417 = 6'hf == _T_584 ? welem[15] : _GEN_6416; // @[Execute.scala 117:10]
  assign _GEN_6418 = 6'h10 == _T_584 ? welem[16] : _GEN_6417; // @[Execute.scala 117:10]
  assign _GEN_6419 = 6'h11 == _T_584 ? welem[17] : _GEN_6418; // @[Execute.scala 117:10]
  assign _GEN_6420 = 6'h12 == _T_584 ? welem[18] : _GEN_6419; // @[Execute.scala 117:10]
  assign _GEN_6421 = 6'h13 == _T_584 ? welem[19] : _GEN_6420; // @[Execute.scala 117:10]
  assign _GEN_6422 = 6'h14 == _T_584 ? welem[20] : _GEN_6421; // @[Execute.scala 117:10]
  assign _GEN_6423 = 6'h15 == _T_584 ? welem[21] : _GEN_6422; // @[Execute.scala 117:10]
  assign _GEN_6424 = 6'h16 == _T_584 ? welem[22] : _GEN_6423; // @[Execute.scala 117:10]
  assign _GEN_6425 = 6'h17 == _T_584 ? welem[23] : _GEN_6424; // @[Execute.scala 117:10]
  assign _GEN_6426 = 6'h18 == _T_584 ? welem[24] : _GEN_6425; // @[Execute.scala 117:10]
  assign _GEN_6427 = 6'h19 == _T_584 ? welem[25] : _GEN_6426; // @[Execute.scala 117:10]
  assign _GEN_6428 = 6'h1a == _T_584 ? welem[26] : _GEN_6427; // @[Execute.scala 117:10]
  assign _GEN_6429 = 6'h1b == _T_584 ? welem[27] : _GEN_6428; // @[Execute.scala 117:10]
  assign _GEN_6430 = 6'h1c == _T_584 ? welem[28] : _GEN_6429; // @[Execute.scala 117:10]
  assign _GEN_6431 = 6'h1d == _T_584 ? welem[29] : _GEN_6430; // @[Execute.scala 117:10]
  assign _GEN_6432 = 6'h1e == _T_584 ? welem[30] : _GEN_6431; // @[Execute.scala 117:10]
  assign _GEN_6433 = 6'h1f == _T_584 ? welem[31] : _GEN_6432; // @[Execute.scala 117:10]
  assign _GEN_6434 = 6'h20 == _T_584 ? welem[32] : _GEN_6433; // @[Execute.scala 117:10]
  assign _GEN_6435 = 6'h21 == _T_584 ? welem[33] : _GEN_6434; // @[Execute.scala 117:10]
  assign _GEN_6436 = 6'h22 == _T_584 ? welem[34] : _GEN_6435; // @[Execute.scala 117:10]
  assign _GEN_6437 = 6'h23 == _T_584 ? welem[35] : _GEN_6436; // @[Execute.scala 117:10]
  assign _GEN_6438 = 6'h24 == _T_584 ? welem[36] : _GEN_6437; // @[Execute.scala 117:10]
  assign _GEN_6439 = 6'h25 == _T_584 ? welem[37] : _GEN_6438; // @[Execute.scala 117:10]
  assign _GEN_6440 = 6'h26 == _T_584 ? welem[38] : _GEN_6439; // @[Execute.scala 117:10]
  assign _GEN_6441 = 6'h27 == _T_584 ? welem[39] : _GEN_6440; // @[Execute.scala 117:10]
  assign _GEN_6442 = 6'h28 == _T_584 ? welem[40] : _GEN_6441; // @[Execute.scala 117:10]
  assign _GEN_6443 = 6'h29 == _T_584 ? welem[41] : _GEN_6442; // @[Execute.scala 117:10]
  assign _GEN_6444 = 6'h2a == _T_584 ? welem[42] : _GEN_6443; // @[Execute.scala 117:10]
  assign _GEN_6445 = 6'h2b == _T_584 ? welem[43] : _GEN_6444; // @[Execute.scala 117:10]
  assign _GEN_6446 = 6'h2c == _T_584 ? welem[44] : _GEN_6445; // @[Execute.scala 117:10]
  assign _GEN_6447 = 6'h2d == _T_584 ? welem[45] : _GEN_6446; // @[Execute.scala 117:10]
  assign _GEN_6448 = 6'h2e == _T_584 ? welem[46] : _GEN_6447; // @[Execute.scala 117:10]
  assign _GEN_6449 = 6'h2f == _T_584 ? welem[47] : _GEN_6448; // @[Execute.scala 117:10]
  assign _GEN_6450 = 6'h30 == _T_584 ? welem[48] : _GEN_6449; // @[Execute.scala 117:10]
  assign _GEN_6451 = 6'h31 == _T_584 ? welem[49] : _GEN_6450; // @[Execute.scala 117:10]
  assign _GEN_6452 = 6'h32 == _T_584 ? welem[50] : _GEN_6451; // @[Execute.scala 117:10]
  assign _GEN_6453 = 6'h33 == _T_584 ? welem[51] : _GEN_6452; // @[Execute.scala 117:10]
  assign _GEN_6454 = 6'h34 == _T_584 ? welem[52] : _GEN_6453; // @[Execute.scala 117:10]
  assign _GEN_6455 = 6'h35 == _T_584 ? welem[53] : _GEN_6454; // @[Execute.scala 117:10]
  assign _GEN_6456 = 6'h36 == _T_584 ? welem[54] : _GEN_6455; // @[Execute.scala 117:10]
  assign _GEN_6457 = 6'h37 == _T_584 ? welem[55] : _GEN_6456; // @[Execute.scala 117:10]
  assign _GEN_6458 = 6'h38 == _T_584 ? welem[56] : _GEN_6457; // @[Execute.scala 117:10]
  assign _GEN_6459 = 6'h39 == _T_584 ? welem[57] : _GEN_6458; // @[Execute.scala 117:10]
  assign _GEN_6460 = 6'h3a == _T_584 ? welem[58] : _GEN_6459; // @[Execute.scala 117:10]
  assign _GEN_6461 = 6'h3b == _T_584 ? welem[59] : _GEN_6460; // @[Execute.scala 117:10]
  assign _GEN_6462 = 6'h3c == _T_584 ? welem[60] : _GEN_6461; // @[Execute.scala 117:10]
  assign _GEN_6463 = 6'h3d == _T_584 ? welem[61] : _GEN_6462; // @[Execute.scala 117:10]
  assign _GEN_6464 = 6'h3e == _T_584 ? welem[62] : _GEN_6463; // @[Execute.scala 117:10]
  assign _GEN_6465 = 6'h3f == _T_584 ? welem[63] : _GEN_6464; // @[Execute.scala 117:10]
  assign _GEN_6467 = 6'h1 == _T_588 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6468 = 6'h2 == _T_588 ? welem[2] : _GEN_6467; // @[Execute.scala 117:10]
  assign _GEN_6469 = 6'h3 == _T_588 ? welem[3] : _GEN_6468; // @[Execute.scala 117:10]
  assign _GEN_6470 = 6'h4 == _T_588 ? welem[4] : _GEN_6469; // @[Execute.scala 117:10]
  assign _GEN_6471 = 6'h5 == _T_588 ? welem[5] : _GEN_6470; // @[Execute.scala 117:10]
  assign _GEN_6472 = 6'h6 == _T_588 ? welem[6] : _GEN_6471; // @[Execute.scala 117:10]
  assign _GEN_6473 = 6'h7 == _T_588 ? welem[7] : _GEN_6472; // @[Execute.scala 117:10]
  assign _GEN_6474 = 6'h8 == _T_588 ? welem[8] : _GEN_6473; // @[Execute.scala 117:10]
  assign _GEN_6475 = 6'h9 == _T_588 ? welem[9] : _GEN_6474; // @[Execute.scala 117:10]
  assign _GEN_6476 = 6'ha == _T_588 ? welem[10] : _GEN_6475; // @[Execute.scala 117:10]
  assign _GEN_6477 = 6'hb == _T_588 ? welem[11] : _GEN_6476; // @[Execute.scala 117:10]
  assign _GEN_6478 = 6'hc == _T_588 ? welem[12] : _GEN_6477; // @[Execute.scala 117:10]
  assign _GEN_6479 = 6'hd == _T_588 ? welem[13] : _GEN_6478; // @[Execute.scala 117:10]
  assign _GEN_6480 = 6'he == _T_588 ? welem[14] : _GEN_6479; // @[Execute.scala 117:10]
  assign _GEN_6481 = 6'hf == _T_588 ? welem[15] : _GEN_6480; // @[Execute.scala 117:10]
  assign _GEN_6482 = 6'h10 == _T_588 ? welem[16] : _GEN_6481; // @[Execute.scala 117:10]
  assign _GEN_6483 = 6'h11 == _T_588 ? welem[17] : _GEN_6482; // @[Execute.scala 117:10]
  assign _GEN_6484 = 6'h12 == _T_588 ? welem[18] : _GEN_6483; // @[Execute.scala 117:10]
  assign _GEN_6485 = 6'h13 == _T_588 ? welem[19] : _GEN_6484; // @[Execute.scala 117:10]
  assign _GEN_6486 = 6'h14 == _T_588 ? welem[20] : _GEN_6485; // @[Execute.scala 117:10]
  assign _GEN_6487 = 6'h15 == _T_588 ? welem[21] : _GEN_6486; // @[Execute.scala 117:10]
  assign _GEN_6488 = 6'h16 == _T_588 ? welem[22] : _GEN_6487; // @[Execute.scala 117:10]
  assign _GEN_6489 = 6'h17 == _T_588 ? welem[23] : _GEN_6488; // @[Execute.scala 117:10]
  assign _GEN_6490 = 6'h18 == _T_588 ? welem[24] : _GEN_6489; // @[Execute.scala 117:10]
  assign _GEN_6491 = 6'h19 == _T_588 ? welem[25] : _GEN_6490; // @[Execute.scala 117:10]
  assign _GEN_6492 = 6'h1a == _T_588 ? welem[26] : _GEN_6491; // @[Execute.scala 117:10]
  assign _GEN_6493 = 6'h1b == _T_588 ? welem[27] : _GEN_6492; // @[Execute.scala 117:10]
  assign _GEN_6494 = 6'h1c == _T_588 ? welem[28] : _GEN_6493; // @[Execute.scala 117:10]
  assign _GEN_6495 = 6'h1d == _T_588 ? welem[29] : _GEN_6494; // @[Execute.scala 117:10]
  assign _GEN_6496 = 6'h1e == _T_588 ? welem[30] : _GEN_6495; // @[Execute.scala 117:10]
  assign _GEN_6497 = 6'h1f == _T_588 ? welem[31] : _GEN_6496; // @[Execute.scala 117:10]
  assign _GEN_6498 = 6'h20 == _T_588 ? welem[32] : _GEN_6497; // @[Execute.scala 117:10]
  assign _GEN_6499 = 6'h21 == _T_588 ? welem[33] : _GEN_6498; // @[Execute.scala 117:10]
  assign _GEN_6500 = 6'h22 == _T_588 ? welem[34] : _GEN_6499; // @[Execute.scala 117:10]
  assign _GEN_6501 = 6'h23 == _T_588 ? welem[35] : _GEN_6500; // @[Execute.scala 117:10]
  assign _GEN_6502 = 6'h24 == _T_588 ? welem[36] : _GEN_6501; // @[Execute.scala 117:10]
  assign _GEN_6503 = 6'h25 == _T_588 ? welem[37] : _GEN_6502; // @[Execute.scala 117:10]
  assign _GEN_6504 = 6'h26 == _T_588 ? welem[38] : _GEN_6503; // @[Execute.scala 117:10]
  assign _GEN_6505 = 6'h27 == _T_588 ? welem[39] : _GEN_6504; // @[Execute.scala 117:10]
  assign _GEN_6506 = 6'h28 == _T_588 ? welem[40] : _GEN_6505; // @[Execute.scala 117:10]
  assign _GEN_6507 = 6'h29 == _T_588 ? welem[41] : _GEN_6506; // @[Execute.scala 117:10]
  assign _GEN_6508 = 6'h2a == _T_588 ? welem[42] : _GEN_6507; // @[Execute.scala 117:10]
  assign _GEN_6509 = 6'h2b == _T_588 ? welem[43] : _GEN_6508; // @[Execute.scala 117:10]
  assign _GEN_6510 = 6'h2c == _T_588 ? welem[44] : _GEN_6509; // @[Execute.scala 117:10]
  assign _GEN_6511 = 6'h2d == _T_588 ? welem[45] : _GEN_6510; // @[Execute.scala 117:10]
  assign _GEN_6512 = 6'h2e == _T_588 ? welem[46] : _GEN_6511; // @[Execute.scala 117:10]
  assign _GEN_6513 = 6'h2f == _T_588 ? welem[47] : _GEN_6512; // @[Execute.scala 117:10]
  assign _GEN_6514 = 6'h30 == _T_588 ? welem[48] : _GEN_6513; // @[Execute.scala 117:10]
  assign _GEN_6515 = 6'h31 == _T_588 ? welem[49] : _GEN_6514; // @[Execute.scala 117:10]
  assign _GEN_6516 = 6'h32 == _T_588 ? welem[50] : _GEN_6515; // @[Execute.scala 117:10]
  assign _GEN_6517 = 6'h33 == _T_588 ? welem[51] : _GEN_6516; // @[Execute.scala 117:10]
  assign _GEN_6518 = 6'h34 == _T_588 ? welem[52] : _GEN_6517; // @[Execute.scala 117:10]
  assign _GEN_6519 = 6'h35 == _T_588 ? welem[53] : _GEN_6518; // @[Execute.scala 117:10]
  assign _GEN_6520 = 6'h36 == _T_588 ? welem[54] : _GEN_6519; // @[Execute.scala 117:10]
  assign _GEN_6521 = 6'h37 == _T_588 ? welem[55] : _GEN_6520; // @[Execute.scala 117:10]
  assign _GEN_6522 = 6'h38 == _T_588 ? welem[56] : _GEN_6521; // @[Execute.scala 117:10]
  assign _GEN_6523 = 6'h39 == _T_588 ? welem[57] : _GEN_6522; // @[Execute.scala 117:10]
  assign _GEN_6524 = 6'h3a == _T_588 ? welem[58] : _GEN_6523; // @[Execute.scala 117:10]
  assign _GEN_6525 = 6'h3b == _T_588 ? welem[59] : _GEN_6524; // @[Execute.scala 117:10]
  assign _GEN_6526 = 6'h3c == _T_588 ? welem[60] : _GEN_6525; // @[Execute.scala 117:10]
  assign _GEN_6527 = 6'h3d == _T_588 ? welem[61] : _GEN_6526; // @[Execute.scala 117:10]
  assign _GEN_6528 = 6'h3e == _T_588 ? welem[62] : _GEN_6527; // @[Execute.scala 117:10]
  assign _GEN_6529 = 6'h3f == _T_588 ? welem[63] : _GEN_6528; // @[Execute.scala 117:10]
  assign _T_591 = _T_582 ? _GEN_6465 : _GEN_6529; // @[Execute.scala 117:10]
  assign _T_592 = r < 6'he; // @[Execute.scala 117:15]
  assign _T_594 = r - 6'he; // @[Execute.scala 117:37]
  assign _T_598 = 6'h32 + r; // @[Execute.scala 117:60]
  assign _GEN_6531 = 6'h1 == _T_594 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6532 = 6'h2 == _T_594 ? welem[2] : _GEN_6531; // @[Execute.scala 117:10]
  assign _GEN_6533 = 6'h3 == _T_594 ? welem[3] : _GEN_6532; // @[Execute.scala 117:10]
  assign _GEN_6534 = 6'h4 == _T_594 ? welem[4] : _GEN_6533; // @[Execute.scala 117:10]
  assign _GEN_6535 = 6'h5 == _T_594 ? welem[5] : _GEN_6534; // @[Execute.scala 117:10]
  assign _GEN_6536 = 6'h6 == _T_594 ? welem[6] : _GEN_6535; // @[Execute.scala 117:10]
  assign _GEN_6537 = 6'h7 == _T_594 ? welem[7] : _GEN_6536; // @[Execute.scala 117:10]
  assign _GEN_6538 = 6'h8 == _T_594 ? welem[8] : _GEN_6537; // @[Execute.scala 117:10]
  assign _GEN_6539 = 6'h9 == _T_594 ? welem[9] : _GEN_6538; // @[Execute.scala 117:10]
  assign _GEN_6540 = 6'ha == _T_594 ? welem[10] : _GEN_6539; // @[Execute.scala 117:10]
  assign _GEN_6541 = 6'hb == _T_594 ? welem[11] : _GEN_6540; // @[Execute.scala 117:10]
  assign _GEN_6542 = 6'hc == _T_594 ? welem[12] : _GEN_6541; // @[Execute.scala 117:10]
  assign _GEN_6543 = 6'hd == _T_594 ? welem[13] : _GEN_6542; // @[Execute.scala 117:10]
  assign _GEN_6544 = 6'he == _T_594 ? welem[14] : _GEN_6543; // @[Execute.scala 117:10]
  assign _GEN_6545 = 6'hf == _T_594 ? welem[15] : _GEN_6544; // @[Execute.scala 117:10]
  assign _GEN_6546 = 6'h10 == _T_594 ? welem[16] : _GEN_6545; // @[Execute.scala 117:10]
  assign _GEN_6547 = 6'h11 == _T_594 ? welem[17] : _GEN_6546; // @[Execute.scala 117:10]
  assign _GEN_6548 = 6'h12 == _T_594 ? welem[18] : _GEN_6547; // @[Execute.scala 117:10]
  assign _GEN_6549 = 6'h13 == _T_594 ? welem[19] : _GEN_6548; // @[Execute.scala 117:10]
  assign _GEN_6550 = 6'h14 == _T_594 ? welem[20] : _GEN_6549; // @[Execute.scala 117:10]
  assign _GEN_6551 = 6'h15 == _T_594 ? welem[21] : _GEN_6550; // @[Execute.scala 117:10]
  assign _GEN_6552 = 6'h16 == _T_594 ? welem[22] : _GEN_6551; // @[Execute.scala 117:10]
  assign _GEN_6553 = 6'h17 == _T_594 ? welem[23] : _GEN_6552; // @[Execute.scala 117:10]
  assign _GEN_6554 = 6'h18 == _T_594 ? welem[24] : _GEN_6553; // @[Execute.scala 117:10]
  assign _GEN_6555 = 6'h19 == _T_594 ? welem[25] : _GEN_6554; // @[Execute.scala 117:10]
  assign _GEN_6556 = 6'h1a == _T_594 ? welem[26] : _GEN_6555; // @[Execute.scala 117:10]
  assign _GEN_6557 = 6'h1b == _T_594 ? welem[27] : _GEN_6556; // @[Execute.scala 117:10]
  assign _GEN_6558 = 6'h1c == _T_594 ? welem[28] : _GEN_6557; // @[Execute.scala 117:10]
  assign _GEN_6559 = 6'h1d == _T_594 ? welem[29] : _GEN_6558; // @[Execute.scala 117:10]
  assign _GEN_6560 = 6'h1e == _T_594 ? welem[30] : _GEN_6559; // @[Execute.scala 117:10]
  assign _GEN_6561 = 6'h1f == _T_594 ? welem[31] : _GEN_6560; // @[Execute.scala 117:10]
  assign _GEN_6562 = 6'h20 == _T_594 ? welem[32] : _GEN_6561; // @[Execute.scala 117:10]
  assign _GEN_6563 = 6'h21 == _T_594 ? welem[33] : _GEN_6562; // @[Execute.scala 117:10]
  assign _GEN_6564 = 6'h22 == _T_594 ? welem[34] : _GEN_6563; // @[Execute.scala 117:10]
  assign _GEN_6565 = 6'h23 == _T_594 ? welem[35] : _GEN_6564; // @[Execute.scala 117:10]
  assign _GEN_6566 = 6'h24 == _T_594 ? welem[36] : _GEN_6565; // @[Execute.scala 117:10]
  assign _GEN_6567 = 6'h25 == _T_594 ? welem[37] : _GEN_6566; // @[Execute.scala 117:10]
  assign _GEN_6568 = 6'h26 == _T_594 ? welem[38] : _GEN_6567; // @[Execute.scala 117:10]
  assign _GEN_6569 = 6'h27 == _T_594 ? welem[39] : _GEN_6568; // @[Execute.scala 117:10]
  assign _GEN_6570 = 6'h28 == _T_594 ? welem[40] : _GEN_6569; // @[Execute.scala 117:10]
  assign _GEN_6571 = 6'h29 == _T_594 ? welem[41] : _GEN_6570; // @[Execute.scala 117:10]
  assign _GEN_6572 = 6'h2a == _T_594 ? welem[42] : _GEN_6571; // @[Execute.scala 117:10]
  assign _GEN_6573 = 6'h2b == _T_594 ? welem[43] : _GEN_6572; // @[Execute.scala 117:10]
  assign _GEN_6574 = 6'h2c == _T_594 ? welem[44] : _GEN_6573; // @[Execute.scala 117:10]
  assign _GEN_6575 = 6'h2d == _T_594 ? welem[45] : _GEN_6574; // @[Execute.scala 117:10]
  assign _GEN_6576 = 6'h2e == _T_594 ? welem[46] : _GEN_6575; // @[Execute.scala 117:10]
  assign _GEN_6577 = 6'h2f == _T_594 ? welem[47] : _GEN_6576; // @[Execute.scala 117:10]
  assign _GEN_6578 = 6'h30 == _T_594 ? welem[48] : _GEN_6577; // @[Execute.scala 117:10]
  assign _GEN_6579 = 6'h31 == _T_594 ? welem[49] : _GEN_6578; // @[Execute.scala 117:10]
  assign _GEN_6580 = 6'h32 == _T_594 ? welem[50] : _GEN_6579; // @[Execute.scala 117:10]
  assign _GEN_6581 = 6'h33 == _T_594 ? welem[51] : _GEN_6580; // @[Execute.scala 117:10]
  assign _GEN_6582 = 6'h34 == _T_594 ? welem[52] : _GEN_6581; // @[Execute.scala 117:10]
  assign _GEN_6583 = 6'h35 == _T_594 ? welem[53] : _GEN_6582; // @[Execute.scala 117:10]
  assign _GEN_6584 = 6'h36 == _T_594 ? welem[54] : _GEN_6583; // @[Execute.scala 117:10]
  assign _GEN_6585 = 6'h37 == _T_594 ? welem[55] : _GEN_6584; // @[Execute.scala 117:10]
  assign _GEN_6586 = 6'h38 == _T_594 ? welem[56] : _GEN_6585; // @[Execute.scala 117:10]
  assign _GEN_6587 = 6'h39 == _T_594 ? welem[57] : _GEN_6586; // @[Execute.scala 117:10]
  assign _GEN_6588 = 6'h3a == _T_594 ? welem[58] : _GEN_6587; // @[Execute.scala 117:10]
  assign _GEN_6589 = 6'h3b == _T_594 ? welem[59] : _GEN_6588; // @[Execute.scala 117:10]
  assign _GEN_6590 = 6'h3c == _T_594 ? welem[60] : _GEN_6589; // @[Execute.scala 117:10]
  assign _GEN_6591 = 6'h3d == _T_594 ? welem[61] : _GEN_6590; // @[Execute.scala 117:10]
  assign _GEN_6592 = 6'h3e == _T_594 ? welem[62] : _GEN_6591; // @[Execute.scala 117:10]
  assign _GEN_6593 = 6'h3f == _T_594 ? welem[63] : _GEN_6592; // @[Execute.scala 117:10]
  assign _GEN_6595 = 6'h1 == _T_598 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6596 = 6'h2 == _T_598 ? welem[2] : _GEN_6595; // @[Execute.scala 117:10]
  assign _GEN_6597 = 6'h3 == _T_598 ? welem[3] : _GEN_6596; // @[Execute.scala 117:10]
  assign _GEN_6598 = 6'h4 == _T_598 ? welem[4] : _GEN_6597; // @[Execute.scala 117:10]
  assign _GEN_6599 = 6'h5 == _T_598 ? welem[5] : _GEN_6598; // @[Execute.scala 117:10]
  assign _GEN_6600 = 6'h6 == _T_598 ? welem[6] : _GEN_6599; // @[Execute.scala 117:10]
  assign _GEN_6601 = 6'h7 == _T_598 ? welem[7] : _GEN_6600; // @[Execute.scala 117:10]
  assign _GEN_6602 = 6'h8 == _T_598 ? welem[8] : _GEN_6601; // @[Execute.scala 117:10]
  assign _GEN_6603 = 6'h9 == _T_598 ? welem[9] : _GEN_6602; // @[Execute.scala 117:10]
  assign _GEN_6604 = 6'ha == _T_598 ? welem[10] : _GEN_6603; // @[Execute.scala 117:10]
  assign _GEN_6605 = 6'hb == _T_598 ? welem[11] : _GEN_6604; // @[Execute.scala 117:10]
  assign _GEN_6606 = 6'hc == _T_598 ? welem[12] : _GEN_6605; // @[Execute.scala 117:10]
  assign _GEN_6607 = 6'hd == _T_598 ? welem[13] : _GEN_6606; // @[Execute.scala 117:10]
  assign _GEN_6608 = 6'he == _T_598 ? welem[14] : _GEN_6607; // @[Execute.scala 117:10]
  assign _GEN_6609 = 6'hf == _T_598 ? welem[15] : _GEN_6608; // @[Execute.scala 117:10]
  assign _GEN_6610 = 6'h10 == _T_598 ? welem[16] : _GEN_6609; // @[Execute.scala 117:10]
  assign _GEN_6611 = 6'h11 == _T_598 ? welem[17] : _GEN_6610; // @[Execute.scala 117:10]
  assign _GEN_6612 = 6'h12 == _T_598 ? welem[18] : _GEN_6611; // @[Execute.scala 117:10]
  assign _GEN_6613 = 6'h13 == _T_598 ? welem[19] : _GEN_6612; // @[Execute.scala 117:10]
  assign _GEN_6614 = 6'h14 == _T_598 ? welem[20] : _GEN_6613; // @[Execute.scala 117:10]
  assign _GEN_6615 = 6'h15 == _T_598 ? welem[21] : _GEN_6614; // @[Execute.scala 117:10]
  assign _GEN_6616 = 6'h16 == _T_598 ? welem[22] : _GEN_6615; // @[Execute.scala 117:10]
  assign _GEN_6617 = 6'h17 == _T_598 ? welem[23] : _GEN_6616; // @[Execute.scala 117:10]
  assign _GEN_6618 = 6'h18 == _T_598 ? welem[24] : _GEN_6617; // @[Execute.scala 117:10]
  assign _GEN_6619 = 6'h19 == _T_598 ? welem[25] : _GEN_6618; // @[Execute.scala 117:10]
  assign _GEN_6620 = 6'h1a == _T_598 ? welem[26] : _GEN_6619; // @[Execute.scala 117:10]
  assign _GEN_6621 = 6'h1b == _T_598 ? welem[27] : _GEN_6620; // @[Execute.scala 117:10]
  assign _GEN_6622 = 6'h1c == _T_598 ? welem[28] : _GEN_6621; // @[Execute.scala 117:10]
  assign _GEN_6623 = 6'h1d == _T_598 ? welem[29] : _GEN_6622; // @[Execute.scala 117:10]
  assign _GEN_6624 = 6'h1e == _T_598 ? welem[30] : _GEN_6623; // @[Execute.scala 117:10]
  assign _GEN_6625 = 6'h1f == _T_598 ? welem[31] : _GEN_6624; // @[Execute.scala 117:10]
  assign _GEN_6626 = 6'h20 == _T_598 ? welem[32] : _GEN_6625; // @[Execute.scala 117:10]
  assign _GEN_6627 = 6'h21 == _T_598 ? welem[33] : _GEN_6626; // @[Execute.scala 117:10]
  assign _GEN_6628 = 6'h22 == _T_598 ? welem[34] : _GEN_6627; // @[Execute.scala 117:10]
  assign _GEN_6629 = 6'h23 == _T_598 ? welem[35] : _GEN_6628; // @[Execute.scala 117:10]
  assign _GEN_6630 = 6'h24 == _T_598 ? welem[36] : _GEN_6629; // @[Execute.scala 117:10]
  assign _GEN_6631 = 6'h25 == _T_598 ? welem[37] : _GEN_6630; // @[Execute.scala 117:10]
  assign _GEN_6632 = 6'h26 == _T_598 ? welem[38] : _GEN_6631; // @[Execute.scala 117:10]
  assign _GEN_6633 = 6'h27 == _T_598 ? welem[39] : _GEN_6632; // @[Execute.scala 117:10]
  assign _GEN_6634 = 6'h28 == _T_598 ? welem[40] : _GEN_6633; // @[Execute.scala 117:10]
  assign _GEN_6635 = 6'h29 == _T_598 ? welem[41] : _GEN_6634; // @[Execute.scala 117:10]
  assign _GEN_6636 = 6'h2a == _T_598 ? welem[42] : _GEN_6635; // @[Execute.scala 117:10]
  assign _GEN_6637 = 6'h2b == _T_598 ? welem[43] : _GEN_6636; // @[Execute.scala 117:10]
  assign _GEN_6638 = 6'h2c == _T_598 ? welem[44] : _GEN_6637; // @[Execute.scala 117:10]
  assign _GEN_6639 = 6'h2d == _T_598 ? welem[45] : _GEN_6638; // @[Execute.scala 117:10]
  assign _GEN_6640 = 6'h2e == _T_598 ? welem[46] : _GEN_6639; // @[Execute.scala 117:10]
  assign _GEN_6641 = 6'h2f == _T_598 ? welem[47] : _GEN_6640; // @[Execute.scala 117:10]
  assign _GEN_6642 = 6'h30 == _T_598 ? welem[48] : _GEN_6641; // @[Execute.scala 117:10]
  assign _GEN_6643 = 6'h31 == _T_598 ? welem[49] : _GEN_6642; // @[Execute.scala 117:10]
  assign _GEN_6644 = 6'h32 == _T_598 ? welem[50] : _GEN_6643; // @[Execute.scala 117:10]
  assign _GEN_6645 = 6'h33 == _T_598 ? welem[51] : _GEN_6644; // @[Execute.scala 117:10]
  assign _GEN_6646 = 6'h34 == _T_598 ? welem[52] : _GEN_6645; // @[Execute.scala 117:10]
  assign _GEN_6647 = 6'h35 == _T_598 ? welem[53] : _GEN_6646; // @[Execute.scala 117:10]
  assign _GEN_6648 = 6'h36 == _T_598 ? welem[54] : _GEN_6647; // @[Execute.scala 117:10]
  assign _GEN_6649 = 6'h37 == _T_598 ? welem[55] : _GEN_6648; // @[Execute.scala 117:10]
  assign _GEN_6650 = 6'h38 == _T_598 ? welem[56] : _GEN_6649; // @[Execute.scala 117:10]
  assign _GEN_6651 = 6'h39 == _T_598 ? welem[57] : _GEN_6650; // @[Execute.scala 117:10]
  assign _GEN_6652 = 6'h3a == _T_598 ? welem[58] : _GEN_6651; // @[Execute.scala 117:10]
  assign _GEN_6653 = 6'h3b == _T_598 ? welem[59] : _GEN_6652; // @[Execute.scala 117:10]
  assign _GEN_6654 = 6'h3c == _T_598 ? welem[60] : _GEN_6653; // @[Execute.scala 117:10]
  assign _GEN_6655 = 6'h3d == _T_598 ? welem[61] : _GEN_6654; // @[Execute.scala 117:10]
  assign _GEN_6656 = 6'h3e == _T_598 ? welem[62] : _GEN_6655; // @[Execute.scala 117:10]
  assign _GEN_6657 = 6'h3f == _T_598 ? welem[63] : _GEN_6656; // @[Execute.scala 117:10]
  assign _T_601 = _T_592 ? _GEN_6593 : _GEN_6657; // @[Execute.scala 117:10]
  assign _T_602 = r < 6'hd; // @[Execute.scala 117:15]
  assign _T_604 = r - 6'hd; // @[Execute.scala 117:37]
  assign _T_608 = 6'h33 + r; // @[Execute.scala 117:60]
  assign _GEN_6659 = 6'h1 == _T_604 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6660 = 6'h2 == _T_604 ? welem[2] : _GEN_6659; // @[Execute.scala 117:10]
  assign _GEN_6661 = 6'h3 == _T_604 ? welem[3] : _GEN_6660; // @[Execute.scala 117:10]
  assign _GEN_6662 = 6'h4 == _T_604 ? welem[4] : _GEN_6661; // @[Execute.scala 117:10]
  assign _GEN_6663 = 6'h5 == _T_604 ? welem[5] : _GEN_6662; // @[Execute.scala 117:10]
  assign _GEN_6664 = 6'h6 == _T_604 ? welem[6] : _GEN_6663; // @[Execute.scala 117:10]
  assign _GEN_6665 = 6'h7 == _T_604 ? welem[7] : _GEN_6664; // @[Execute.scala 117:10]
  assign _GEN_6666 = 6'h8 == _T_604 ? welem[8] : _GEN_6665; // @[Execute.scala 117:10]
  assign _GEN_6667 = 6'h9 == _T_604 ? welem[9] : _GEN_6666; // @[Execute.scala 117:10]
  assign _GEN_6668 = 6'ha == _T_604 ? welem[10] : _GEN_6667; // @[Execute.scala 117:10]
  assign _GEN_6669 = 6'hb == _T_604 ? welem[11] : _GEN_6668; // @[Execute.scala 117:10]
  assign _GEN_6670 = 6'hc == _T_604 ? welem[12] : _GEN_6669; // @[Execute.scala 117:10]
  assign _GEN_6671 = 6'hd == _T_604 ? welem[13] : _GEN_6670; // @[Execute.scala 117:10]
  assign _GEN_6672 = 6'he == _T_604 ? welem[14] : _GEN_6671; // @[Execute.scala 117:10]
  assign _GEN_6673 = 6'hf == _T_604 ? welem[15] : _GEN_6672; // @[Execute.scala 117:10]
  assign _GEN_6674 = 6'h10 == _T_604 ? welem[16] : _GEN_6673; // @[Execute.scala 117:10]
  assign _GEN_6675 = 6'h11 == _T_604 ? welem[17] : _GEN_6674; // @[Execute.scala 117:10]
  assign _GEN_6676 = 6'h12 == _T_604 ? welem[18] : _GEN_6675; // @[Execute.scala 117:10]
  assign _GEN_6677 = 6'h13 == _T_604 ? welem[19] : _GEN_6676; // @[Execute.scala 117:10]
  assign _GEN_6678 = 6'h14 == _T_604 ? welem[20] : _GEN_6677; // @[Execute.scala 117:10]
  assign _GEN_6679 = 6'h15 == _T_604 ? welem[21] : _GEN_6678; // @[Execute.scala 117:10]
  assign _GEN_6680 = 6'h16 == _T_604 ? welem[22] : _GEN_6679; // @[Execute.scala 117:10]
  assign _GEN_6681 = 6'h17 == _T_604 ? welem[23] : _GEN_6680; // @[Execute.scala 117:10]
  assign _GEN_6682 = 6'h18 == _T_604 ? welem[24] : _GEN_6681; // @[Execute.scala 117:10]
  assign _GEN_6683 = 6'h19 == _T_604 ? welem[25] : _GEN_6682; // @[Execute.scala 117:10]
  assign _GEN_6684 = 6'h1a == _T_604 ? welem[26] : _GEN_6683; // @[Execute.scala 117:10]
  assign _GEN_6685 = 6'h1b == _T_604 ? welem[27] : _GEN_6684; // @[Execute.scala 117:10]
  assign _GEN_6686 = 6'h1c == _T_604 ? welem[28] : _GEN_6685; // @[Execute.scala 117:10]
  assign _GEN_6687 = 6'h1d == _T_604 ? welem[29] : _GEN_6686; // @[Execute.scala 117:10]
  assign _GEN_6688 = 6'h1e == _T_604 ? welem[30] : _GEN_6687; // @[Execute.scala 117:10]
  assign _GEN_6689 = 6'h1f == _T_604 ? welem[31] : _GEN_6688; // @[Execute.scala 117:10]
  assign _GEN_6690 = 6'h20 == _T_604 ? welem[32] : _GEN_6689; // @[Execute.scala 117:10]
  assign _GEN_6691 = 6'h21 == _T_604 ? welem[33] : _GEN_6690; // @[Execute.scala 117:10]
  assign _GEN_6692 = 6'h22 == _T_604 ? welem[34] : _GEN_6691; // @[Execute.scala 117:10]
  assign _GEN_6693 = 6'h23 == _T_604 ? welem[35] : _GEN_6692; // @[Execute.scala 117:10]
  assign _GEN_6694 = 6'h24 == _T_604 ? welem[36] : _GEN_6693; // @[Execute.scala 117:10]
  assign _GEN_6695 = 6'h25 == _T_604 ? welem[37] : _GEN_6694; // @[Execute.scala 117:10]
  assign _GEN_6696 = 6'h26 == _T_604 ? welem[38] : _GEN_6695; // @[Execute.scala 117:10]
  assign _GEN_6697 = 6'h27 == _T_604 ? welem[39] : _GEN_6696; // @[Execute.scala 117:10]
  assign _GEN_6698 = 6'h28 == _T_604 ? welem[40] : _GEN_6697; // @[Execute.scala 117:10]
  assign _GEN_6699 = 6'h29 == _T_604 ? welem[41] : _GEN_6698; // @[Execute.scala 117:10]
  assign _GEN_6700 = 6'h2a == _T_604 ? welem[42] : _GEN_6699; // @[Execute.scala 117:10]
  assign _GEN_6701 = 6'h2b == _T_604 ? welem[43] : _GEN_6700; // @[Execute.scala 117:10]
  assign _GEN_6702 = 6'h2c == _T_604 ? welem[44] : _GEN_6701; // @[Execute.scala 117:10]
  assign _GEN_6703 = 6'h2d == _T_604 ? welem[45] : _GEN_6702; // @[Execute.scala 117:10]
  assign _GEN_6704 = 6'h2e == _T_604 ? welem[46] : _GEN_6703; // @[Execute.scala 117:10]
  assign _GEN_6705 = 6'h2f == _T_604 ? welem[47] : _GEN_6704; // @[Execute.scala 117:10]
  assign _GEN_6706 = 6'h30 == _T_604 ? welem[48] : _GEN_6705; // @[Execute.scala 117:10]
  assign _GEN_6707 = 6'h31 == _T_604 ? welem[49] : _GEN_6706; // @[Execute.scala 117:10]
  assign _GEN_6708 = 6'h32 == _T_604 ? welem[50] : _GEN_6707; // @[Execute.scala 117:10]
  assign _GEN_6709 = 6'h33 == _T_604 ? welem[51] : _GEN_6708; // @[Execute.scala 117:10]
  assign _GEN_6710 = 6'h34 == _T_604 ? welem[52] : _GEN_6709; // @[Execute.scala 117:10]
  assign _GEN_6711 = 6'h35 == _T_604 ? welem[53] : _GEN_6710; // @[Execute.scala 117:10]
  assign _GEN_6712 = 6'h36 == _T_604 ? welem[54] : _GEN_6711; // @[Execute.scala 117:10]
  assign _GEN_6713 = 6'h37 == _T_604 ? welem[55] : _GEN_6712; // @[Execute.scala 117:10]
  assign _GEN_6714 = 6'h38 == _T_604 ? welem[56] : _GEN_6713; // @[Execute.scala 117:10]
  assign _GEN_6715 = 6'h39 == _T_604 ? welem[57] : _GEN_6714; // @[Execute.scala 117:10]
  assign _GEN_6716 = 6'h3a == _T_604 ? welem[58] : _GEN_6715; // @[Execute.scala 117:10]
  assign _GEN_6717 = 6'h3b == _T_604 ? welem[59] : _GEN_6716; // @[Execute.scala 117:10]
  assign _GEN_6718 = 6'h3c == _T_604 ? welem[60] : _GEN_6717; // @[Execute.scala 117:10]
  assign _GEN_6719 = 6'h3d == _T_604 ? welem[61] : _GEN_6718; // @[Execute.scala 117:10]
  assign _GEN_6720 = 6'h3e == _T_604 ? welem[62] : _GEN_6719; // @[Execute.scala 117:10]
  assign _GEN_6721 = 6'h3f == _T_604 ? welem[63] : _GEN_6720; // @[Execute.scala 117:10]
  assign _GEN_6723 = 6'h1 == _T_608 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6724 = 6'h2 == _T_608 ? welem[2] : _GEN_6723; // @[Execute.scala 117:10]
  assign _GEN_6725 = 6'h3 == _T_608 ? welem[3] : _GEN_6724; // @[Execute.scala 117:10]
  assign _GEN_6726 = 6'h4 == _T_608 ? welem[4] : _GEN_6725; // @[Execute.scala 117:10]
  assign _GEN_6727 = 6'h5 == _T_608 ? welem[5] : _GEN_6726; // @[Execute.scala 117:10]
  assign _GEN_6728 = 6'h6 == _T_608 ? welem[6] : _GEN_6727; // @[Execute.scala 117:10]
  assign _GEN_6729 = 6'h7 == _T_608 ? welem[7] : _GEN_6728; // @[Execute.scala 117:10]
  assign _GEN_6730 = 6'h8 == _T_608 ? welem[8] : _GEN_6729; // @[Execute.scala 117:10]
  assign _GEN_6731 = 6'h9 == _T_608 ? welem[9] : _GEN_6730; // @[Execute.scala 117:10]
  assign _GEN_6732 = 6'ha == _T_608 ? welem[10] : _GEN_6731; // @[Execute.scala 117:10]
  assign _GEN_6733 = 6'hb == _T_608 ? welem[11] : _GEN_6732; // @[Execute.scala 117:10]
  assign _GEN_6734 = 6'hc == _T_608 ? welem[12] : _GEN_6733; // @[Execute.scala 117:10]
  assign _GEN_6735 = 6'hd == _T_608 ? welem[13] : _GEN_6734; // @[Execute.scala 117:10]
  assign _GEN_6736 = 6'he == _T_608 ? welem[14] : _GEN_6735; // @[Execute.scala 117:10]
  assign _GEN_6737 = 6'hf == _T_608 ? welem[15] : _GEN_6736; // @[Execute.scala 117:10]
  assign _GEN_6738 = 6'h10 == _T_608 ? welem[16] : _GEN_6737; // @[Execute.scala 117:10]
  assign _GEN_6739 = 6'h11 == _T_608 ? welem[17] : _GEN_6738; // @[Execute.scala 117:10]
  assign _GEN_6740 = 6'h12 == _T_608 ? welem[18] : _GEN_6739; // @[Execute.scala 117:10]
  assign _GEN_6741 = 6'h13 == _T_608 ? welem[19] : _GEN_6740; // @[Execute.scala 117:10]
  assign _GEN_6742 = 6'h14 == _T_608 ? welem[20] : _GEN_6741; // @[Execute.scala 117:10]
  assign _GEN_6743 = 6'h15 == _T_608 ? welem[21] : _GEN_6742; // @[Execute.scala 117:10]
  assign _GEN_6744 = 6'h16 == _T_608 ? welem[22] : _GEN_6743; // @[Execute.scala 117:10]
  assign _GEN_6745 = 6'h17 == _T_608 ? welem[23] : _GEN_6744; // @[Execute.scala 117:10]
  assign _GEN_6746 = 6'h18 == _T_608 ? welem[24] : _GEN_6745; // @[Execute.scala 117:10]
  assign _GEN_6747 = 6'h19 == _T_608 ? welem[25] : _GEN_6746; // @[Execute.scala 117:10]
  assign _GEN_6748 = 6'h1a == _T_608 ? welem[26] : _GEN_6747; // @[Execute.scala 117:10]
  assign _GEN_6749 = 6'h1b == _T_608 ? welem[27] : _GEN_6748; // @[Execute.scala 117:10]
  assign _GEN_6750 = 6'h1c == _T_608 ? welem[28] : _GEN_6749; // @[Execute.scala 117:10]
  assign _GEN_6751 = 6'h1d == _T_608 ? welem[29] : _GEN_6750; // @[Execute.scala 117:10]
  assign _GEN_6752 = 6'h1e == _T_608 ? welem[30] : _GEN_6751; // @[Execute.scala 117:10]
  assign _GEN_6753 = 6'h1f == _T_608 ? welem[31] : _GEN_6752; // @[Execute.scala 117:10]
  assign _GEN_6754 = 6'h20 == _T_608 ? welem[32] : _GEN_6753; // @[Execute.scala 117:10]
  assign _GEN_6755 = 6'h21 == _T_608 ? welem[33] : _GEN_6754; // @[Execute.scala 117:10]
  assign _GEN_6756 = 6'h22 == _T_608 ? welem[34] : _GEN_6755; // @[Execute.scala 117:10]
  assign _GEN_6757 = 6'h23 == _T_608 ? welem[35] : _GEN_6756; // @[Execute.scala 117:10]
  assign _GEN_6758 = 6'h24 == _T_608 ? welem[36] : _GEN_6757; // @[Execute.scala 117:10]
  assign _GEN_6759 = 6'h25 == _T_608 ? welem[37] : _GEN_6758; // @[Execute.scala 117:10]
  assign _GEN_6760 = 6'h26 == _T_608 ? welem[38] : _GEN_6759; // @[Execute.scala 117:10]
  assign _GEN_6761 = 6'h27 == _T_608 ? welem[39] : _GEN_6760; // @[Execute.scala 117:10]
  assign _GEN_6762 = 6'h28 == _T_608 ? welem[40] : _GEN_6761; // @[Execute.scala 117:10]
  assign _GEN_6763 = 6'h29 == _T_608 ? welem[41] : _GEN_6762; // @[Execute.scala 117:10]
  assign _GEN_6764 = 6'h2a == _T_608 ? welem[42] : _GEN_6763; // @[Execute.scala 117:10]
  assign _GEN_6765 = 6'h2b == _T_608 ? welem[43] : _GEN_6764; // @[Execute.scala 117:10]
  assign _GEN_6766 = 6'h2c == _T_608 ? welem[44] : _GEN_6765; // @[Execute.scala 117:10]
  assign _GEN_6767 = 6'h2d == _T_608 ? welem[45] : _GEN_6766; // @[Execute.scala 117:10]
  assign _GEN_6768 = 6'h2e == _T_608 ? welem[46] : _GEN_6767; // @[Execute.scala 117:10]
  assign _GEN_6769 = 6'h2f == _T_608 ? welem[47] : _GEN_6768; // @[Execute.scala 117:10]
  assign _GEN_6770 = 6'h30 == _T_608 ? welem[48] : _GEN_6769; // @[Execute.scala 117:10]
  assign _GEN_6771 = 6'h31 == _T_608 ? welem[49] : _GEN_6770; // @[Execute.scala 117:10]
  assign _GEN_6772 = 6'h32 == _T_608 ? welem[50] : _GEN_6771; // @[Execute.scala 117:10]
  assign _GEN_6773 = 6'h33 == _T_608 ? welem[51] : _GEN_6772; // @[Execute.scala 117:10]
  assign _GEN_6774 = 6'h34 == _T_608 ? welem[52] : _GEN_6773; // @[Execute.scala 117:10]
  assign _GEN_6775 = 6'h35 == _T_608 ? welem[53] : _GEN_6774; // @[Execute.scala 117:10]
  assign _GEN_6776 = 6'h36 == _T_608 ? welem[54] : _GEN_6775; // @[Execute.scala 117:10]
  assign _GEN_6777 = 6'h37 == _T_608 ? welem[55] : _GEN_6776; // @[Execute.scala 117:10]
  assign _GEN_6778 = 6'h38 == _T_608 ? welem[56] : _GEN_6777; // @[Execute.scala 117:10]
  assign _GEN_6779 = 6'h39 == _T_608 ? welem[57] : _GEN_6778; // @[Execute.scala 117:10]
  assign _GEN_6780 = 6'h3a == _T_608 ? welem[58] : _GEN_6779; // @[Execute.scala 117:10]
  assign _GEN_6781 = 6'h3b == _T_608 ? welem[59] : _GEN_6780; // @[Execute.scala 117:10]
  assign _GEN_6782 = 6'h3c == _T_608 ? welem[60] : _GEN_6781; // @[Execute.scala 117:10]
  assign _GEN_6783 = 6'h3d == _T_608 ? welem[61] : _GEN_6782; // @[Execute.scala 117:10]
  assign _GEN_6784 = 6'h3e == _T_608 ? welem[62] : _GEN_6783; // @[Execute.scala 117:10]
  assign _GEN_6785 = 6'h3f == _T_608 ? welem[63] : _GEN_6784; // @[Execute.scala 117:10]
  assign _T_611 = _T_602 ? _GEN_6721 : _GEN_6785; // @[Execute.scala 117:10]
  assign _T_612 = r < 6'hc; // @[Execute.scala 117:15]
  assign _T_614 = r - 6'hc; // @[Execute.scala 117:37]
  assign _T_618 = 6'h34 + r; // @[Execute.scala 117:60]
  assign _GEN_6787 = 6'h1 == _T_614 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6788 = 6'h2 == _T_614 ? welem[2] : _GEN_6787; // @[Execute.scala 117:10]
  assign _GEN_6789 = 6'h3 == _T_614 ? welem[3] : _GEN_6788; // @[Execute.scala 117:10]
  assign _GEN_6790 = 6'h4 == _T_614 ? welem[4] : _GEN_6789; // @[Execute.scala 117:10]
  assign _GEN_6791 = 6'h5 == _T_614 ? welem[5] : _GEN_6790; // @[Execute.scala 117:10]
  assign _GEN_6792 = 6'h6 == _T_614 ? welem[6] : _GEN_6791; // @[Execute.scala 117:10]
  assign _GEN_6793 = 6'h7 == _T_614 ? welem[7] : _GEN_6792; // @[Execute.scala 117:10]
  assign _GEN_6794 = 6'h8 == _T_614 ? welem[8] : _GEN_6793; // @[Execute.scala 117:10]
  assign _GEN_6795 = 6'h9 == _T_614 ? welem[9] : _GEN_6794; // @[Execute.scala 117:10]
  assign _GEN_6796 = 6'ha == _T_614 ? welem[10] : _GEN_6795; // @[Execute.scala 117:10]
  assign _GEN_6797 = 6'hb == _T_614 ? welem[11] : _GEN_6796; // @[Execute.scala 117:10]
  assign _GEN_6798 = 6'hc == _T_614 ? welem[12] : _GEN_6797; // @[Execute.scala 117:10]
  assign _GEN_6799 = 6'hd == _T_614 ? welem[13] : _GEN_6798; // @[Execute.scala 117:10]
  assign _GEN_6800 = 6'he == _T_614 ? welem[14] : _GEN_6799; // @[Execute.scala 117:10]
  assign _GEN_6801 = 6'hf == _T_614 ? welem[15] : _GEN_6800; // @[Execute.scala 117:10]
  assign _GEN_6802 = 6'h10 == _T_614 ? welem[16] : _GEN_6801; // @[Execute.scala 117:10]
  assign _GEN_6803 = 6'h11 == _T_614 ? welem[17] : _GEN_6802; // @[Execute.scala 117:10]
  assign _GEN_6804 = 6'h12 == _T_614 ? welem[18] : _GEN_6803; // @[Execute.scala 117:10]
  assign _GEN_6805 = 6'h13 == _T_614 ? welem[19] : _GEN_6804; // @[Execute.scala 117:10]
  assign _GEN_6806 = 6'h14 == _T_614 ? welem[20] : _GEN_6805; // @[Execute.scala 117:10]
  assign _GEN_6807 = 6'h15 == _T_614 ? welem[21] : _GEN_6806; // @[Execute.scala 117:10]
  assign _GEN_6808 = 6'h16 == _T_614 ? welem[22] : _GEN_6807; // @[Execute.scala 117:10]
  assign _GEN_6809 = 6'h17 == _T_614 ? welem[23] : _GEN_6808; // @[Execute.scala 117:10]
  assign _GEN_6810 = 6'h18 == _T_614 ? welem[24] : _GEN_6809; // @[Execute.scala 117:10]
  assign _GEN_6811 = 6'h19 == _T_614 ? welem[25] : _GEN_6810; // @[Execute.scala 117:10]
  assign _GEN_6812 = 6'h1a == _T_614 ? welem[26] : _GEN_6811; // @[Execute.scala 117:10]
  assign _GEN_6813 = 6'h1b == _T_614 ? welem[27] : _GEN_6812; // @[Execute.scala 117:10]
  assign _GEN_6814 = 6'h1c == _T_614 ? welem[28] : _GEN_6813; // @[Execute.scala 117:10]
  assign _GEN_6815 = 6'h1d == _T_614 ? welem[29] : _GEN_6814; // @[Execute.scala 117:10]
  assign _GEN_6816 = 6'h1e == _T_614 ? welem[30] : _GEN_6815; // @[Execute.scala 117:10]
  assign _GEN_6817 = 6'h1f == _T_614 ? welem[31] : _GEN_6816; // @[Execute.scala 117:10]
  assign _GEN_6818 = 6'h20 == _T_614 ? welem[32] : _GEN_6817; // @[Execute.scala 117:10]
  assign _GEN_6819 = 6'h21 == _T_614 ? welem[33] : _GEN_6818; // @[Execute.scala 117:10]
  assign _GEN_6820 = 6'h22 == _T_614 ? welem[34] : _GEN_6819; // @[Execute.scala 117:10]
  assign _GEN_6821 = 6'h23 == _T_614 ? welem[35] : _GEN_6820; // @[Execute.scala 117:10]
  assign _GEN_6822 = 6'h24 == _T_614 ? welem[36] : _GEN_6821; // @[Execute.scala 117:10]
  assign _GEN_6823 = 6'h25 == _T_614 ? welem[37] : _GEN_6822; // @[Execute.scala 117:10]
  assign _GEN_6824 = 6'h26 == _T_614 ? welem[38] : _GEN_6823; // @[Execute.scala 117:10]
  assign _GEN_6825 = 6'h27 == _T_614 ? welem[39] : _GEN_6824; // @[Execute.scala 117:10]
  assign _GEN_6826 = 6'h28 == _T_614 ? welem[40] : _GEN_6825; // @[Execute.scala 117:10]
  assign _GEN_6827 = 6'h29 == _T_614 ? welem[41] : _GEN_6826; // @[Execute.scala 117:10]
  assign _GEN_6828 = 6'h2a == _T_614 ? welem[42] : _GEN_6827; // @[Execute.scala 117:10]
  assign _GEN_6829 = 6'h2b == _T_614 ? welem[43] : _GEN_6828; // @[Execute.scala 117:10]
  assign _GEN_6830 = 6'h2c == _T_614 ? welem[44] : _GEN_6829; // @[Execute.scala 117:10]
  assign _GEN_6831 = 6'h2d == _T_614 ? welem[45] : _GEN_6830; // @[Execute.scala 117:10]
  assign _GEN_6832 = 6'h2e == _T_614 ? welem[46] : _GEN_6831; // @[Execute.scala 117:10]
  assign _GEN_6833 = 6'h2f == _T_614 ? welem[47] : _GEN_6832; // @[Execute.scala 117:10]
  assign _GEN_6834 = 6'h30 == _T_614 ? welem[48] : _GEN_6833; // @[Execute.scala 117:10]
  assign _GEN_6835 = 6'h31 == _T_614 ? welem[49] : _GEN_6834; // @[Execute.scala 117:10]
  assign _GEN_6836 = 6'h32 == _T_614 ? welem[50] : _GEN_6835; // @[Execute.scala 117:10]
  assign _GEN_6837 = 6'h33 == _T_614 ? welem[51] : _GEN_6836; // @[Execute.scala 117:10]
  assign _GEN_6838 = 6'h34 == _T_614 ? welem[52] : _GEN_6837; // @[Execute.scala 117:10]
  assign _GEN_6839 = 6'h35 == _T_614 ? welem[53] : _GEN_6838; // @[Execute.scala 117:10]
  assign _GEN_6840 = 6'h36 == _T_614 ? welem[54] : _GEN_6839; // @[Execute.scala 117:10]
  assign _GEN_6841 = 6'h37 == _T_614 ? welem[55] : _GEN_6840; // @[Execute.scala 117:10]
  assign _GEN_6842 = 6'h38 == _T_614 ? welem[56] : _GEN_6841; // @[Execute.scala 117:10]
  assign _GEN_6843 = 6'h39 == _T_614 ? welem[57] : _GEN_6842; // @[Execute.scala 117:10]
  assign _GEN_6844 = 6'h3a == _T_614 ? welem[58] : _GEN_6843; // @[Execute.scala 117:10]
  assign _GEN_6845 = 6'h3b == _T_614 ? welem[59] : _GEN_6844; // @[Execute.scala 117:10]
  assign _GEN_6846 = 6'h3c == _T_614 ? welem[60] : _GEN_6845; // @[Execute.scala 117:10]
  assign _GEN_6847 = 6'h3d == _T_614 ? welem[61] : _GEN_6846; // @[Execute.scala 117:10]
  assign _GEN_6848 = 6'h3e == _T_614 ? welem[62] : _GEN_6847; // @[Execute.scala 117:10]
  assign _GEN_6849 = 6'h3f == _T_614 ? welem[63] : _GEN_6848; // @[Execute.scala 117:10]
  assign _GEN_6851 = 6'h1 == _T_618 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6852 = 6'h2 == _T_618 ? welem[2] : _GEN_6851; // @[Execute.scala 117:10]
  assign _GEN_6853 = 6'h3 == _T_618 ? welem[3] : _GEN_6852; // @[Execute.scala 117:10]
  assign _GEN_6854 = 6'h4 == _T_618 ? welem[4] : _GEN_6853; // @[Execute.scala 117:10]
  assign _GEN_6855 = 6'h5 == _T_618 ? welem[5] : _GEN_6854; // @[Execute.scala 117:10]
  assign _GEN_6856 = 6'h6 == _T_618 ? welem[6] : _GEN_6855; // @[Execute.scala 117:10]
  assign _GEN_6857 = 6'h7 == _T_618 ? welem[7] : _GEN_6856; // @[Execute.scala 117:10]
  assign _GEN_6858 = 6'h8 == _T_618 ? welem[8] : _GEN_6857; // @[Execute.scala 117:10]
  assign _GEN_6859 = 6'h9 == _T_618 ? welem[9] : _GEN_6858; // @[Execute.scala 117:10]
  assign _GEN_6860 = 6'ha == _T_618 ? welem[10] : _GEN_6859; // @[Execute.scala 117:10]
  assign _GEN_6861 = 6'hb == _T_618 ? welem[11] : _GEN_6860; // @[Execute.scala 117:10]
  assign _GEN_6862 = 6'hc == _T_618 ? welem[12] : _GEN_6861; // @[Execute.scala 117:10]
  assign _GEN_6863 = 6'hd == _T_618 ? welem[13] : _GEN_6862; // @[Execute.scala 117:10]
  assign _GEN_6864 = 6'he == _T_618 ? welem[14] : _GEN_6863; // @[Execute.scala 117:10]
  assign _GEN_6865 = 6'hf == _T_618 ? welem[15] : _GEN_6864; // @[Execute.scala 117:10]
  assign _GEN_6866 = 6'h10 == _T_618 ? welem[16] : _GEN_6865; // @[Execute.scala 117:10]
  assign _GEN_6867 = 6'h11 == _T_618 ? welem[17] : _GEN_6866; // @[Execute.scala 117:10]
  assign _GEN_6868 = 6'h12 == _T_618 ? welem[18] : _GEN_6867; // @[Execute.scala 117:10]
  assign _GEN_6869 = 6'h13 == _T_618 ? welem[19] : _GEN_6868; // @[Execute.scala 117:10]
  assign _GEN_6870 = 6'h14 == _T_618 ? welem[20] : _GEN_6869; // @[Execute.scala 117:10]
  assign _GEN_6871 = 6'h15 == _T_618 ? welem[21] : _GEN_6870; // @[Execute.scala 117:10]
  assign _GEN_6872 = 6'h16 == _T_618 ? welem[22] : _GEN_6871; // @[Execute.scala 117:10]
  assign _GEN_6873 = 6'h17 == _T_618 ? welem[23] : _GEN_6872; // @[Execute.scala 117:10]
  assign _GEN_6874 = 6'h18 == _T_618 ? welem[24] : _GEN_6873; // @[Execute.scala 117:10]
  assign _GEN_6875 = 6'h19 == _T_618 ? welem[25] : _GEN_6874; // @[Execute.scala 117:10]
  assign _GEN_6876 = 6'h1a == _T_618 ? welem[26] : _GEN_6875; // @[Execute.scala 117:10]
  assign _GEN_6877 = 6'h1b == _T_618 ? welem[27] : _GEN_6876; // @[Execute.scala 117:10]
  assign _GEN_6878 = 6'h1c == _T_618 ? welem[28] : _GEN_6877; // @[Execute.scala 117:10]
  assign _GEN_6879 = 6'h1d == _T_618 ? welem[29] : _GEN_6878; // @[Execute.scala 117:10]
  assign _GEN_6880 = 6'h1e == _T_618 ? welem[30] : _GEN_6879; // @[Execute.scala 117:10]
  assign _GEN_6881 = 6'h1f == _T_618 ? welem[31] : _GEN_6880; // @[Execute.scala 117:10]
  assign _GEN_6882 = 6'h20 == _T_618 ? welem[32] : _GEN_6881; // @[Execute.scala 117:10]
  assign _GEN_6883 = 6'h21 == _T_618 ? welem[33] : _GEN_6882; // @[Execute.scala 117:10]
  assign _GEN_6884 = 6'h22 == _T_618 ? welem[34] : _GEN_6883; // @[Execute.scala 117:10]
  assign _GEN_6885 = 6'h23 == _T_618 ? welem[35] : _GEN_6884; // @[Execute.scala 117:10]
  assign _GEN_6886 = 6'h24 == _T_618 ? welem[36] : _GEN_6885; // @[Execute.scala 117:10]
  assign _GEN_6887 = 6'h25 == _T_618 ? welem[37] : _GEN_6886; // @[Execute.scala 117:10]
  assign _GEN_6888 = 6'h26 == _T_618 ? welem[38] : _GEN_6887; // @[Execute.scala 117:10]
  assign _GEN_6889 = 6'h27 == _T_618 ? welem[39] : _GEN_6888; // @[Execute.scala 117:10]
  assign _GEN_6890 = 6'h28 == _T_618 ? welem[40] : _GEN_6889; // @[Execute.scala 117:10]
  assign _GEN_6891 = 6'h29 == _T_618 ? welem[41] : _GEN_6890; // @[Execute.scala 117:10]
  assign _GEN_6892 = 6'h2a == _T_618 ? welem[42] : _GEN_6891; // @[Execute.scala 117:10]
  assign _GEN_6893 = 6'h2b == _T_618 ? welem[43] : _GEN_6892; // @[Execute.scala 117:10]
  assign _GEN_6894 = 6'h2c == _T_618 ? welem[44] : _GEN_6893; // @[Execute.scala 117:10]
  assign _GEN_6895 = 6'h2d == _T_618 ? welem[45] : _GEN_6894; // @[Execute.scala 117:10]
  assign _GEN_6896 = 6'h2e == _T_618 ? welem[46] : _GEN_6895; // @[Execute.scala 117:10]
  assign _GEN_6897 = 6'h2f == _T_618 ? welem[47] : _GEN_6896; // @[Execute.scala 117:10]
  assign _GEN_6898 = 6'h30 == _T_618 ? welem[48] : _GEN_6897; // @[Execute.scala 117:10]
  assign _GEN_6899 = 6'h31 == _T_618 ? welem[49] : _GEN_6898; // @[Execute.scala 117:10]
  assign _GEN_6900 = 6'h32 == _T_618 ? welem[50] : _GEN_6899; // @[Execute.scala 117:10]
  assign _GEN_6901 = 6'h33 == _T_618 ? welem[51] : _GEN_6900; // @[Execute.scala 117:10]
  assign _GEN_6902 = 6'h34 == _T_618 ? welem[52] : _GEN_6901; // @[Execute.scala 117:10]
  assign _GEN_6903 = 6'h35 == _T_618 ? welem[53] : _GEN_6902; // @[Execute.scala 117:10]
  assign _GEN_6904 = 6'h36 == _T_618 ? welem[54] : _GEN_6903; // @[Execute.scala 117:10]
  assign _GEN_6905 = 6'h37 == _T_618 ? welem[55] : _GEN_6904; // @[Execute.scala 117:10]
  assign _GEN_6906 = 6'h38 == _T_618 ? welem[56] : _GEN_6905; // @[Execute.scala 117:10]
  assign _GEN_6907 = 6'h39 == _T_618 ? welem[57] : _GEN_6906; // @[Execute.scala 117:10]
  assign _GEN_6908 = 6'h3a == _T_618 ? welem[58] : _GEN_6907; // @[Execute.scala 117:10]
  assign _GEN_6909 = 6'h3b == _T_618 ? welem[59] : _GEN_6908; // @[Execute.scala 117:10]
  assign _GEN_6910 = 6'h3c == _T_618 ? welem[60] : _GEN_6909; // @[Execute.scala 117:10]
  assign _GEN_6911 = 6'h3d == _T_618 ? welem[61] : _GEN_6910; // @[Execute.scala 117:10]
  assign _GEN_6912 = 6'h3e == _T_618 ? welem[62] : _GEN_6911; // @[Execute.scala 117:10]
  assign _GEN_6913 = 6'h3f == _T_618 ? welem[63] : _GEN_6912; // @[Execute.scala 117:10]
  assign _T_621 = _T_612 ? _GEN_6849 : _GEN_6913; // @[Execute.scala 117:10]
  assign _T_622 = r < 6'hb; // @[Execute.scala 117:15]
  assign _T_624 = r - 6'hb; // @[Execute.scala 117:37]
  assign _T_628 = 6'h35 + r; // @[Execute.scala 117:60]
  assign _GEN_6915 = 6'h1 == _T_624 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6916 = 6'h2 == _T_624 ? welem[2] : _GEN_6915; // @[Execute.scala 117:10]
  assign _GEN_6917 = 6'h3 == _T_624 ? welem[3] : _GEN_6916; // @[Execute.scala 117:10]
  assign _GEN_6918 = 6'h4 == _T_624 ? welem[4] : _GEN_6917; // @[Execute.scala 117:10]
  assign _GEN_6919 = 6'h5 == _T_624 ? welem[5] : _GEN_6918; // @[Execute.scala 117:10]
  assign _GEN_6920 = 6'h6 == _T_624 ? welem[6] : _GEN_6919; // @[Execute.scala 117:10]
  assign _GEN_6921 = 6'h7 == _T_624 ? welem[7] : _GEN_6920; // @[Execute.scala 117:10]
  assign _GEN_6922 = 6'h8 == _T_624 ? welem[8] : _GEN_6921; // @[Execute.scala 117:10]
  assign _GEN_6923 = 6'h9 == _T_624 ? welem[9] : _GEN_6922; // @[Execute.scala 117:10]
  assign _GEN_6924 = 6'ha == _T_624 ? welem[10] : _GEN_6923; // @[Execute.scala 117:10]
  assign _GEN_6925 = 6'hb == _T_624 ? welem[11] : _GEN_6924; // @[Execute.scala 117:10]
  assign _GEN_6926 = 6'hc == _T_624 ? welem[12] : _GEN_6925; // @[Execute.scala 117:10]
  assign _GEN_6927 = 6'hd == _T_624 ? welem[13] : _GEN_6926; // @[Execute.scala 117:10]
  assign _GEN_6928 = 6'he == _T_624 ? welem[14] : _GEN_6927; // @[Execute.scala 117:10]
  assign _GEN_6929 = 6'hf == _T_624 ? welem[15] : _GEN_6928; // @[Execute.scala 117:10]
  assign _GEN_6930 = 6'h10 == _T_624 ? welem[16] : _GEN_6929; // @[Execute.scala 117:10]
  assign _GEN_6931 = 6'h11 == _T_624 ? welem[17] : _GEN_6930; // @[Execute.scala 117:10]
  assign _GEN_6932 = 6'h12 == _T_624 ? welem[18] : _GEN_6931; // @[Execute.scala 117:10]
  assign _GEN_6933 = 6'h13 == _T_624 ? welem[19] : _GEN_6932; // @[Execute.scala 117:10]
  assign _GEN_6934 = 6'h14 == _T_624 ? welem[20] : _GEN_6933; // @[Execute.scala 117:10]
  assign _GEN_6935 = 6'h15 == _T_624 ? welem[21] : _GEN_6934; // @[Execute.scala 117:10]
  assign _GEN_6936 = 6'h16 == _T_624 ? welem[22] : _GEN_6935; // @[Execute.scala 117:10]
  assign _GEN_6937 = 6'h17 == _T_624 ? welem[23] : _GEN_6936; // @[Execute.scala 117:10]
  assign _GEN_6938 = 6'h18 == _T_624 ? welem[24] : _GEN_6937; // @[Execute.scala 117:10]
  assign _GEN_6939 = 6'h19 == _T_624 ? welem[25] : _GEN_6938; // @[Execute.scala 117:10]
  assign _GEN_6940 = 6'h1a == _T_624 ? welem[26] : _GEN_6939; // @[Execute.scala 117:10]
  assign _GEN_6941 = 6'h1b == _T_624 ? welem[27] : _GEN_6940; // @[Execute.scala 117:10]
  assign _GEN_6942 = 6'h1c == _T_624 ? welem[28] : _GEN_6941; // @[Execute.scala 117:10]
  assign _GEN_6943 = 6'h1d == _T_624 ? welem[29] : _GEN_6942; // @[Execute.scala 117:10]
  assign _GEN_6944 = 6'h1e == _T_624 ? welem[30] : _GEN_6943; // @[Execute.scala 117:10]
  assign _GEN_6945 = 6'h1f == _T_624 ? welem[31] : _GEN_6944; // @[Execute.scala 117:10]
  assign _GEN_6946 = 6'h20 == _T_624 ? welem[32] : _GEN_6945; // @[Execute.scala 117:10]
  assign _GEN_6947 = 6'h21 == _T_624 ? welem[33] : _GEN_6946; // @[Execute.scala 117:10]
  assign _GEN_6948 = 6'h22 == _T_624 ? welem[34] : _GEN_6947; // @[Execute.scala 117:10]
  assign _GEN_6949 = 6'h23 == _T_624 ? welem[35] : _GEN_6948; // @[Execute.scala 117:10]
  assign _GEN_6950 = 6'h24 == _T_624 ? welem[36] : _GEN_6949; // @[Execute.scala 117:10]
  assign _GEN_6951 = 6'h25 == _T_624 ? welem[37] : _GEN_6950; // @[Execute.scala 117:10]
  assign _GEN_6952 = 6'h26 == _T_624 ? welem[38] : _GEN_6951; // @[Execute.scala 117:10]
  assign _GEN_6953 = 6'h27 == _T_624 ? welem[39] : _GEN_6952; // @[Execute.scala 117:10]
  assign _GEN_6954 = 6'h28 == _T_624 ? welem[40] : _GEN_6953; // @[Execute.scala 117:10]
  assign _GEN_6955 = 6'h29 == _T_624 ? welem[41] : _GEN_6954; // @[Execute.scala 117:10]
  assign _GEN_6956 = 6'h2a == _T_624 ? welem[42] : _GEN_6955; // @[Execute.scala 117:10]
  assign _GEN_6957 = 6'h2b == _T_624 ? welem[43] : _GEN_6956; // @[Execute.scala 117:10]
  assign _GEN_6958 = 6'h2c == _T_624 ? welem[44] : _GEN_6957; // @[Execute.scala 117:10]
  assign _GEN_6959 = 6'h2d == _T_624 ? welem[45] : _GEN_6958; // @[Execute.scala 117:10]
  assign _GEN_6960 = 6'h2e == _T_624 ? welem[46] : _GEN_6959; // @[Execute.scala 117:10]
  assign _GEN_6961 = 6'h2f == _T_624 ? welem[47] : _GEN_6960; // @[Execute.scala 117:10]
  assign _GEN_6962 = 6'h30 == _T_624 ? welem[48] : _GEN_6961; // @[Execute.scala 117:10]
  assign _GEN_6963 = 6'h31 == _T_624 ? welem[49] : _GEN_6962; // @[Execute.scala 117:10]
  assign _GEN_6964 = 6'h32 == _T_624 ? welem[50] : _GEN_6963; // @[Execute.scala 117:10]
  assign _GEN_6965 = 6'h33 == _T_624 ? welem[51] : _GEN_6964; // @[Execute.scala 117:10]
  assign _GEN_6966 = 6'h34 == _T_624 ? welem[52] : _GEN_6965; // @[Execute.scala 117:10]
  assign _GEN_6967 = 6'h35 == _T_624 ? welem[53] : _GEN_6966; // @[Execute.scala 117:10]
  assign _GEN_6968 = 6'h36 == _T_624 ? welem[54] : _GEN_6967; // @[Execute.scala 117:10]
  assign _GEN_6969 = 6'h37 == _T_624 ? welem[55] : _GEN_6968; // @[Execute.scala 117:10]
  assign _GEN_6970 = 6'h38 == _T_624 ? welem[56] : _GEN_6969; // @[Execute.scala 117:10]
  assign _GEN_6971 = 6'h39 == _T_624 ? welem[57] : _GEN_6970; // @[Execute.scala 117:10]
  assign _GEN_6972 = 6'h3a == _T_624 ? welem[58] : _GEN_6971; // @[Execute.scala 117:10]
  assign _GEN_6973 = 6'h3b == _T_624 ? welem[59] : _GEN_6972; // @[Execute.scala 117:10]
  assign _GEN_6974 = 6'h3c == _T_624 ? welem[60] : _GEN_6973; // @[Execute.scala 117:10]
  assign _GEN_6975 = 6'h3d == _T_624 ? welem[61] : _GEN_6974; // @[Execute.scala 117:10]
  assign _GEN_6976 = 6'h3e == _T_624 ? welem[62] : _GEN_6975; // @[Execute.scala 117:10]
  assign _GEN_6977 = 6'h3f == _T_624 ? welem[63] : _GEN_6976; // @[Execute.scala 117:10]
  assign _GEN_6979 = 6'h1 == _T_628 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_6980 = 6'h2 == _T_628 ? welem[2] : _GEN_6979; // @[Execute.scala 117:10]
  assign _GEN_6981 = 6'h3 == _T_628 ? welem[3] : _GEN_6980; // @[Execute.scala 117:10]
  assign _GEN_6982 = 6'h4 == _T_628 ? welem[4] : _GEN_6981; // @[Execute.scala 117:10]
  assign _GEN_6983 = 6'h5 == _T_628 ? welem[5] : _GEN_6982; // @[Execute.scala 117:10]
  assign _GEN_6984 = 6'h6 == _T_628 ? welem[6] : _GEN_6983; // @[Execute.scala 117:10]
  assign _GEN_6985 = 6'h7 == _T_628 ? welem[7] : _GEN_6984; // @[Execute.scala 117:10]
  assign _GEN_6986 = 6'h8 == _T_628 ? welem[8] : _GEN_6985; // @[Execute.scala 117:10]
  assign _GEN_6987 = 6'h9 == _T_628 ? welem[9] : _GEN_6986; // @[Execute.scala 117:10]
  assign _GEN_6988 = 6'ha == _T_628 ? welem[10] : _GEN_6987; // @[Execute.scala 117:10]
  assign _GEN_6989 = 6'hb == _T_628 ? welem[11] : _GEN_6988; // @[Execute.scala 117:10]
  assign _GEN_6990 = 6'hc == _T_628 ? welem[12] : _GEN_6989; // @[Execute.scala 117:10]
  assign _GEN_6991 = 6'hd == _T_628 ? welem[13] : _GEN_6990; // @[Execute.scala 117:10]
  assign _GEN_6992 = 6'he == _T_628 ? welem[14] : _GEN_6991; // @[Execute.scala 117:10]
  assign _GEN_6993 = 6'hf == _T_628 ? welem[15] : _GEN_6992; // @[Execute.scala 117:10]
  assign _GEN_6994 = 6'h10 == _T_628 ? welem[16] : _GEN_6993; // @[Execute.scala 117:10]
  assign _GEN_6995 = 6'h11 == _T_628 ? welem[17] : _GEN_6994; // @[Execute.scala 117:10]
  assign _GEN_6996 = 6'h12 == _T_628 ? welem[18] : _GEN_6995; // @[Execute.scala 117:10]
  assign _GEN_6997 = 6'h13 == _T_628 ? welem[19] : _GEN_6996; // @[Execute.scala 117:10]
  assign _GEN_6998 = 6'h14 == _T_628 ? welem[20] : _GEN_6997; // @[Execute.scala 117:10]
  assign _GEN_6999 = 6'h15 == _T_628 ? welem[21] : _GEN_6998; // @[Execute.scala 117:10]
  assign _GEN_7000 = 6'h16 == _T_628 ? welem[22] : _GEN_6999; // @[Execute.scala 117:10]
  assign _GEN_7001 = 6'h17 == _T_628 ? welem[23] : _GEN_7000; // @[Execute.scala 117:10]
  assign _GEN_7002 = 6'h18 == _T_628 ? welem[24] : _GEN_7001; // @[Execute.scala 117:10]
  assign _GEN_7003 = 6'h19 == _T_628 ? welem[25] : _GEN_7002; // @[Execute.scala 117:10]
  assign _GEN_7004 = 6'h1a == _T_628 ? welem[26] : _GEN_7003; // @[Execute.scala 117:10]
  assign _GEN_7005 = 6'h1b == _T_628 ? welem[27] : _GEN_7004; // @[Execute.scala 117:10]
  assign _GEN_7006 = 6'h1c == _T_628 ? welem[28] : _GEN_7005; // @[Execute.scala 117:10]
  assign _GEN_7007 = 6'h1d == _T_628 ? welem[29] : _GEN_7006; // @[Execute.scala 117:10]
  assign _GEN_7008 = 6'h1e == _T_628 ? welem[30] : _GEN_7007; // @[Execute.scala 117:10]
  assign _GEN_7009 = 6'h1f == _T_628 ? welem[31] : _GEN_7008; // @[Execute.scala 117:10]
  assign _GEN_7010 = 6'h20 == _T_628 ? welem[32] : _GEN_7009; // @[Execute.scala 117:10]
  assign _GEN_7011 = 6'h21 == _T_628 ? welem[33] : _GEN_7010; // @[Execute.scala 117:10]
  assign _GEN_7012 = 6'h22 == _T_628 ? welem[34] : _GEN_7011; // @[Execute.scala 117:10]
  assign _GEN_7013 = 6'h23 == _T_628 ? welem[35] : _GEN_7012; // @[Execute.scala 117:10]
  assign _GEN_7014 = 6'h24 == _T_628 ? welem[36] : _GEN_7013; // @[Execute.scala 117:10]
  assign _GEN_7015 = 6'h25 == _T_628 ? welem[37] : _GEN_7014; // @[Execute.scala 117:10]
  assign _GEN_7016 = 6'h26 == _T_628 ? welem[38] : _GEN_7015; // @[Execute.scala 117:10]
  assign _GEN_7017 = 6'h27 == _T_628 ? welem[39] : _GEN_7016; // @[Execute.scala 117:10]
  assign _GEN_7018 = 6'h28 == _T_628 ? welem[40] : _GEN_7017; // @[Execute.scala 117:10]
  assign _GEN_7019 = 6'h29 == _T_628 ? welem[41] : _GEN_7018; // @[Execute.scala 117:10]
  assign _GEN_7020 = 6'h2a == _T_628 ? welem[42] : _GEN_7019; // @[Execute.scala 117:10]
  assign _GEN_7021 = 6'h2b == _T_628 ? welem[43] : _GEN_7020; // @[Execute.scala 117:10]
  assign _GEN_7022 = 6'h2c == _T_628 ? welem[44] : _GEN_7021; // @[Execute.scala 117:10]
  assign _GEN_7023 = 6'h2d == _T_628 ? welem[45] : _GEN_7022; // @[Execute.scala 117:10]
  assign _GEN_7024 = 6'h2e == _T_628 ? welem[46] : _GEN_7023; // @[Execute.scala 117:10]
  assign _GEN_7025 = 6'h2f == _T_628 ? welem[47] : _GEN_7024; // @[Execute.scala 117:10]
  assign _GEN_7026 = 6'h30 == _T_628 ? welem[48] : _GEN_7025; // @[Execute.scala 117:10]
  assign _GEN_7027 = 6'h31 == _T_628 ? welem[49] : _GEN_7026; // @[Execute.scala 117:10]
  assign _GEN_7028 = 6'h32 == _T_628 ? welem[50] : _GEN_7027; // @[Execute.scala 117:10]
  assign _GEN_7029 = 6'h33 == _T_628 ? welem[51] : _GEN_7028; // @[Execute.scala 117:10]
  assign _GEN_7030 = 6'h34 == _T_628 ? welem[52] : _GEN_7029; // @[Execute.scala 117:10]
  assign _GEN_7031 = 6'h35 == _T_628 ? welem[53] : _GEN_7030; // @[Execute.scala 117:10]
  assign _GEN_7032 = 6'h36 == _T_628 ? welem[54] : _GEN_7031; // @[Execute.scala 117:10]
  assign _GEN_7033 = 6'h37 == _T_628 ? welem[55] : _GEN_7032; // @[Execute.scala 117:10]
  assign _GEN_7034 = 6'h38 == _T_628 ? welem[56] : _GEN_7033; // @[Execute.scala 117:10]
  assign _GEN_7035 = 6'h39 == _T_628 ? welem[57] : _GEN_7034; // @[Execute.scala 117:10]
  assign _GEN_7036 = 6'h3a == _T_628 ? welem[58] : _GEN_7035; // @[Execute.scala 117:10]
  assign _GEN_7037 = 6'h3b == _T_628 ? welem[59] : _GEN_7036; // @[Execute.scala 117:10]
  assign _GEN_7038 = 6'h3c == _T_628 ? welem[60] : _GEN_7037; // @[Execute.scala 117:10]
  assign _GEN_7039 = 6'h3d == _T_628 ? welem[61] : _GEN_7038; // @[Execute.scala 117:10]
  assign _GEN_7040 = 6'h3e == _T_628 ? welem[62] : _GEN_7039; // @[Execute.scala 117:10]
  assign _GEN_7041 = 6'h3f == _T_628 ? welem[63] : _GEN_7040; // @[Execute.scala 117:10]
  assign _T_631 = _T_622 ? _GEN_6977 : _GEN_7041; // @[Execute.scala 117:10]
  assign _T_632 = r < 6'ha; // @[Execute.scala 117:15]
  assign _T_634 = r - 6'ha; // @[Execute.scala 117:37]
  assign _T_638 = 6'h36 + r; // @[Execute.scala 117:60]
  assign _GEN_7043 = 6'h1 == _T_634 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7044 = 6'h2 == _T_634 ? welem[2] : _GEN_7043; // @[Execute.scala 117:10]
  assign _GEN_7045 = 6'h3 == _T_634 ? welem[3] : _GEN_7044; // @[Execute.scala 117:10]
  assign _GEN_7046 = 6'h4 == _T_634 ? welem[4] : _GEN_7045; // @[Execute.scala 117:10]
  assign _GEN_7047 = 6'h5 == _T_634 ? welem[5] : _GEN_7046; // @[Execute.scala 117:10]
  assign _GEN_7048 = 6'h6 == _T_634 ? welem[6] : _GEN_7047; // @[Execute.scala 117:10]
  assign _GEN_7049 = 6'h7 == _T_634 ? welem[7] : _GEN_7048; // @[Execute.scala 117:10]
  assign _GEN_7050 = 6'h8 == _T_634 ? welem[8] : _GEN_7049; // @[Execute.scala 117:10]
  assign _GEN_7051 = 6'h9 == _T_634 ? welem[9] : _GEN_7050; // @[Execute.scala 117:10]
  assign _GEN_7052 = 6'ha == _T_634 ? welem[10] : _GEN_7051; // @[Execute.scala 117:10]
  assign _GEN_7053 = 6'hb == _T_634 ? welem[11] : _GEN_7052; // @[Execute.scala 117:10]
  assign _GEN_7054 = 6'hc == _T_634 ? welem[12] : _GEN_7053; // @[Execute.scala 117:10]
  assign _GEN_7055 = 6'hd == _T_634 ? welem[13] : _GEN_7054; // @[Execute.scala 117:10]
  assign _GEN_7056 = 6'he == _T_634 ? welem[14] : _GEN_7055; // @[Execute.scala 117:10]
  assign _GEN_7057 = 6'hf == _T_634 ? welem[15] : _GEN_7056; // @[Execute.scala 117:10]
  assign _GEN_7058 = 6'h10 == _T_634 ? welem[16] : _GEN_7057; // @[Execute.scala 117:10]
  assign _GEN_7059 = 6'h11 == _T_634 ? welem[17] : _GEN_7058; // @[Execute.scala 117:10]
  assign _GEN_7060 = 6'h12 == _T_634 ? welem[18] : _GEN_7059; // @[Execute.scala 117:10]
  assign _GEN_7061 = 6'h13 == _T_634 ? welem[19] : _GEN_7060; // @[Execute.scala 117:10]
  assign _GEN_7062 = 6'h14 == _T_634 ? welem[20] : _GEN_7061; // @[Execute.scala 117:10]
  assign _GEN_7063 = 6'h15 == _T_634 ? welem[21] : _GEN_7062; // @[Execute.scala 117:10]
  assign _GEN_7064 = 6'h16 == _T_634 ? welem[22] : _GEN_7063; // @[Execute.scala 117:10]
  assign _GEN_7065 = 6'h17 == _T_634 ? welem[23] : _GEN_7064; // @[Execute.scala 117:10]
  assign _GEN_7066 = 6'h18 == _T_634 ? welem[24] : _GEN_7065; // @[Execute.scala 117:10]
  assign _GEN_7067 = 6'h19 == _T_634 ? welem[25] : _GEN_7066; // @[Execute.scala 117:10]
  assign _GEN_7068 = 6'h1a == _T_634 ? welem[26] : _GEN_7067; // @[Execute.scala 117:10]
  assign _GEN_7069 = 6'h1b == _T_634 ? welem[27] : _GEN_7068; // @[Execute.scala 117:10]
  assign _GEN_7070 = 6'h1c == _T_634 ? welem[28] : _GEN_7069; // @[Execute.scala 117:10]
  assign _GEN_7071 = 6'h1d == _T_634 ? welem[29] : _GEN_7070; // @[Execute.scala 117:10]
  assign _GEN_7072 = 6'h1e == _T_634 ? welem[30] : _GEN_7071; // @[Execute.scala 117:10]
  assign _GEN_7073 = 6'h1f == _T_634 ? welem[31] : _GEN_7072; // @[Execute.scala 117:10]
  assign _GEN_7074 = 6'h20 == _T_634 ? welem[32] : _GEN_7073; // @[Execute.scala 117:10]
  assign _GEN_7075 = 6'h21 == _T_634 ? welem[33] : _GEN_7074; // @[Execute.scala 117:10]
  assign _GEN_7076 = 6'h22 == _T_634 ? welem[34] : _GEN_7075; // @[Execute.scala 117:10]
  assign _GEN_7077 = 6'h23 == _T_634 ? welem[35] : _GEN_7076; // @[Execute.scala 117:10]
  assign _GEN_7078 = 6'h24 == _T_634 ? welem[36] : _GEN_7077; // @[Execute.scala 117:10]
  assign _GEN_7079 = 6'h25 == _T_634 ? welem[37] : _GEN_7078; // @[Execute.scala 117:10]
  assign _GEN_7080 = 6'h26 == _T_634 ? welem[38] : _GEN_7079; // @[Execute.scala 117:10]
  assign _GEN_7081 = 6'h27 == _T_634 ? welem[39] : _GEN_7080; // @[Execute.scala 117:10]
  assign _GEN_7082 = 6'h28 == _T_634 ? welem[40] : _GEN_7081; // @[Execute.scala 117:10]
  assign _GEN_7083 = 6'h29 == _T_634 ? welem[41] : _GEN_7082; // @[Execute.scala 117:10]
  assign _GEN_7084 = 6'h2a == _T_634 ? welem[42] : _GEN_7083; // @[Execute.scala 117:10]
  assign _GEN_7085 = 6'h2b == _T_634 ? welem[43] : _GEN_7084; // @[Execute.scala 117:10]
  assign _GEN_7086 = 6'h2c == _T_634 ? welem[44] : _GEN_7085; // @[Execute.scala 117:10]
  assign _GEN_7087 = 6'h2d == _T_634 ? welem[45] : _GEN_7086; // @[Execute.scala 117:10]
  assign _GEN_7088 = 6'h2e == _T_634 ? welem[46] : _GEN_7087; // @[Execute.scala 117:10]
  assign _GEN_7089 = 6'h2f == _T_634 ? welem[47] : _GEN_7088; // @[Execute.scala 117:10]
  assign _GEN_7090 = 6'h30 == _T_634 ? welem[48] : _GEN_7089; // @[Execute.scala 117:10]
  assign _GEN_7091 = 6'h31 == _T_634 ? welem[49] : _GEN_7090; // @[Execute.scala 117:10]
  assign _GEN_7092 = 6'h32 == _T_634 ? welem[50] : _GEN_7091; // @[Execute.scala 117:10]
  assign _GEN_7093 = 6'h33 == _T_634 ? welem[51] : _GEN_7092; // @[Execute.scala 117:10]
  assign _GEN_7094 = 6'h34 == _T_634 ? welem[52] : _GEN_7093; // @[Execute.scala 117:10]
  assign _GEN_7095 = 6'h35 == _T_634 ? welem[53] : _GEN_7094; // @[Execute.scala 117:10]
  assign _GEN_7096 = 6'h36 == _T_634 ? welem[54] : _GEN_7095; // @[Execute.scala 117:10]
  assign _GEN_7097 = 6'h37 == _T_634 ? welem[55] : _GEN_7096; // @[Execute.scala 117:10]
  assign _GEN_7098 = 6'h38 == _T_634 ? welem[56] : _GEN_7097; // @[Execute.scala 117:10]
  assign _GEN_7099 = 6'h39 == _T_634 ? welem[57] : _GEN_7098; // @[Execute.scala 117:10]
  assign _GEN_7100 = 6'h3a == _T_634 ? welem[58] : _GEN_7099; // @[Execute.scala 117:10]
  assign _GEN_7101 = 6'h3b == _T_634 ? welem[59] : _GEN_7100; // @[Execute.scala 117:10]
  assign _GEN_7102 = 6'h3c == _T_634 ? welem[60] : _GEN_7101; // @[Execute.scala 117:10]
  assign _GEN_7103 = 6'h3d == _T_634 ? welem[61] : _GEN_7102; // @[Execute.scala 117:10]
  assign _GEN_7104 = 6'h3e == _T_634 ? welem[62] : _GEN_7103; // @[Execute.scala 117:10]
  assign _GEN_7105 = 6'h3f == _T_634 ? welem[63] : _GEN_7104; // @[Execute.scala 117:10]
  assign _GEN_7107 = 6'h1 == _T_638 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7108 = 6'h2 == _T_638 ? welem[2] : _GEN_7107; // @[Execute.scala 117:10]
  assign _GEN_7109 = 6'h3 == _T_638 ? welem[3] : _GEN_7108; // @[Execute.scala 117:10]
  assign _GEN_7110 = 6'h4 == _T_638 ? welem[4] : _GEN_7109; // @[Execute.scala 117:10]
  assign _GEN_7111 = 6'h5 == _T_638 ? welem[5] : _GEN_7110; // @[Execute.scala 117:10]
  assign _GEN_7112 = 6'h6 == _T_638 ? welem[6] : _GEN_7111; // @[Execute.scala 117:10]
  assign _GEN_7113 = 6'h7 == _T_638 ? welem[7] : _GEN_7112; // @[Execute.scala 117:10]
  assign _GEN_7114 = 6'h8 == _T_638 ? welem[8] : _GEN_7113; // @[Execute.scala 117:10]
  assign _GEN_7115 = 6'h9 == _T_638 ? welem[9] : _GEN_7114; // @[Execute.scala 117:10]
  assign _GEN_7116 = 6'ha == _T_638 ? welem[10] : _GEN_7115; // @[Execute.scala 117:10]
  assign _GEN_7117 = 6'hb == _T_638 ? welem[11] : _GEN_7116; // @[Execute.scala 117:10]
  assign _GEN_7118 = 6'hc == _T_638 ? welem[12] : _GEN_7117; // @[Execute.scala 117:10]
  assign _GEN_7119 = 6'hd == _T_638 ? welem[13] : _GEN_7118; // @[Execute.scala 117:10]
  assign _GEN_7120 = 6'he == _T_638 ? welem[14] : _GEN_7119; // @[Execute.scala 117:10]
  assign _GEN_7121 = 6'hf == _T_638 ? welem[15] : _GEN_7120; // @[Execute.scala 117:10]
  assign _GEN_7122 = 6'h10 == _T_638 ? welem[16] : _GEN_7121; // @[Execute.scala 117:10]
  assign _GEN_7123 = 6'h11 == _T_638 ? welem[17] : _GEN_7122; // @[Execute.scala 117:10]
  assign _GEN_7124 = 6'h12 == _T_638 ? welem[18] : _GEN_7123; // @[Execute.scala 117:10]
  assign _GEN_7125 = 6'h13 == _T_638 ? welem[19] : _GEN_7124; // @[Execute.scala 117:10]
  assign _GEN_7126 = 6'h14 == _T_638 ? welem[20] : _GEN_7125; // @[Execute.scala 117:10]
  assign _GEN_7127 = 6'h15 == _T_638 ? welem[21] : _GEN_7126; // @[Execute.scala 117:10]
  assign _GEN_7128 = 6'h16 == _T_638 ? welem[22] : _GEN_7127; // @[Execute.scala 117:10]
  assign _GEN_7129 = 6'h17 == _T_638 ? welem[23] : _GEN_7128; // @[Execute.scala 117:10]
  assign _GEN_7130 = 6'h18 == _T_638 ? welem[24] : _GEN_7129; // @[Execute.scala 117:10]
  assign _GEN_7131 = 6'h19 == _T_638 ? welem[25] : _GEN_7130; // @[Execute.scala 117:10]
  assign _GEN_7132 = 6'h1a == _T_638 ? welem[26] : _GEN_7131; // @[Execute.scala 117:10]
  assign _GEN_7133 = 6'h1b == _T_638 ? welem[27] : _GEN_7132; // @[Execute.scala 117:10]
  assign _GEN_7134 = 6'h1c == _T_638 ? welem[28] : _GEN_7133; // @[Execute.scala 117:10]
  assign _GEN_7135 = 6'h1d == _T_638 ? welem[29] : _GEN_7134; // @[Execute.scala 117:10]
  assign _GEN_7136 = 6'h1e == _T_638 ? welem[30] : _GEN_7135; // @[Execute.scala 117:10]
  assign _GEN_7137 = 6'h1f == _T_638 ? welem[31] : _GEN_7136; // @[Execute.scala 117:10]
  assign _GEN_7138 = 6'h20 == _T_638 ? welem[32] : _GEN_7137; // @[Execute.scala 117:10]
  assign _GEN_7139 = 6'h21 == _T_638 ? welem[33] : _GEN_7138; // @[Execute.scala 117:10]
  assign _GEN_7140 = 6'h22 == _T_638 ? welem[34] : _GEN_7139; // @[Execute.scala 117:10]
  assign _GEN_7141 = 6'h23 == _T_638 ? welem[35] : _GEN_7140; // @[Execute.scala 117:10]
  assign _GEN_7142 = 6'h24 == _T_638 ? welem[36] : _GEN_7141; // @[Execute.scala 117:10]
  assign _GEN_7143 = 6'h25 == _T_638 ? welem[37] : _GEN_7142; // @[Execute.scala 117:10]
  assign _GEN_7144 = 6'h26 == _T_638 ? welem[38] : _GEN_7143; // @[Execute.scala 117:10]
  assign _GEN_7145 = 6'h27 == _T_638 ? welem[39] : _GEN_7144; // @[Execute.scala 117:10]
  assign _GEN_7146 = 6'h28 == _T_638 ? welem[40] : _GEN_7145; // @[Execute.scala 117:10]
  assign _GEN_7147 = 6'h29 == _T_638 ? welem[41] : _GEN_7146; // @[Execute.scala 117:10]
  assign _GEN_7148 = 6'h2a == _T_638 ? welem[42] : _GEN_7147; // @[Execute.scala 117:10]
  assign _GEN_7149 = 6'h2b == _T_638 ? welem[43] : _GEN_7148; // @[Execute.scala 117:10]
  assign _GEN_7150 = 6'h2c == _T_638 ? welem[44] : _GEN_7149; // @[Execute.scala 117:10]
  assign _GEN_7151 = 6'h2d == _T_638 ? welem[45] : _GEN_7150; // @[Execute.scala 117:10]
  assign _GEN_7152 = 6'h2e == _T_638 ? welem[46] : _GEN_7151; // @[Execute.scala 117:10]
  assign _GEN_7153 = 6'h2f == _T_638 ? welem[47] : _GEN_7152; // @[Execute.scala 117:10]
  assign _GEN_7154 = 6'h30 == _T_638 ? welem[48] : _GEN_7153; // @[Execute.scala 117:10]
  assign _GEN_7155 = 6'h31 == _T_638 ? welem[49] : _GEN_7154; // @[Execute.scala 117:10]
  assign _GEN_7156 = 6'h32 == _T_638 ? welem[50] : _GEN_7155; // @[Execute.scala 117:10]
  assign _GEN_7157 = 6'h33 == _T_638 ? welem[51] : _GEN_7156; // @[Execute.scala 117:10]
  assign _GEN_7158 = 6'h34 == _T_638 ? welem[52] : _GEN_7157; // @[Execute.scala 117:10]
  assign _GEN_7159 = 6'h35 == _T_638 ? welem[53] : _GEN_7158; // @[Execute.scala 117:10]
  assign _GEN_7160 = 6'h36 == _T_638 ? welem[54] : _GEN_7159; // @[Execute.scala 117:10]
  assign _GEN_7161 = 6'h37 == _T_638 ? welem[55] : _GEN_7160; // @[Execute.scala 117:10]
  assign _GEN_7162 = 6'h38 == _T_638 ? welem[56] : _GEN_7161; // @[Execute.scala 117:10]
  assign _GEN_7163 = 6'h39 == _T_638 ? welem[57] : _GEN_7162; // @[Execute.scala 117:10]
  assign _GEN_7164 = 6'h3a == _T_638 ? welem[58] : _GEN_7163; // @[Execute.scala 117:10]
  assign _GEN_7165 = 6'h3b == _T_638 ? welem[59] : _GEN_7164; // @[Execute.scala 117:10]
  assign _GEN_7166 = 6'h3c == _T_638 ? welem[60] : _GEN_7165; // @[Execute.scala 117:10]
  assign _GEN_7167 = 6'h3d == _T_638 ? welem[61] : _GEN_7166; // @[Execute.scala 117:10]
  assign _GEN_7168 = 6'h3e == _T_638 ? welem[62] : _GEN_7167; // @[Execute.scala 117:10]
  assign _GEN_7169 = 6'h3f == _T_638 ? welem[63] : _GEN_7168; // @[Execute.scala 117:10]
  assign _T_641 = _T_632 ? _GEN_7105 : _GEN_7169; // @[Execute.scala 117:10]
  assign _T_642 = r < 6'h9; // @[Execute.scala 117:15]
  assign _T_644 = r - 6'h9; // @[Execute.scala 117:37]
  assign _T_648 = 6'h37 + r; // @[Execute.scala 117:60]
  assign _GEN_7171 = 6'h1 == _T_644 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7172 = 6'h2 == _T_644 ? welem[2] : _GEN_7171; // @[Execute.scala 117:10]
  assign _GEN_7173 = 6'h3 == _T_644 ? welem[3] : _GEN_7172; // @[Execute.scala 117:10]
  assign _GEN_7174 = 6'h4 == _T_644 ? welem[4] : _GEN_7173; // @[Execute.scala 117:10]
  assign _GEN_7175 = 6'h5 == _T_644 ? welem[5] : _GEN_7174; // @[Execute.scala 117:10]
  assign _GEN_7176 = 6'h6 == _T_644 ? welem[6] : _GEN_7175; // @[Execute.scala 117:10]
  assign _GEN_7177 = 6'h7 == _T_644 ? welem[7] : _GEN_7176; // @[Execute.scala 117:10]
  assign _GEN_7178 = 6'h8 == _T_644 ? welem[8] : _GEN_7177; // @[Execute.scala 117:10]
  assign _GEN_7179 = 6'h9 == _T_644 ? welem[9] : _GEN_7178; // @[Execute.scala 117:10]
  assign _GEN_7180 = 6'ha == _T_644 ? welem[10] : _GEN_7179; // @[Execute.scala 117:10]
  assign _GEN_7181 = 6'hb == _T_644 ? welem[11] : _GEN_7180; // @[Execute.scala 117:10]
  assign _GEN_7182 = 6'hc == _T_644 ? welem[12] : _GEN_7181; // @[Execute.scala 117:10]
  assign _GEN_7183 = 6'hd == _T_644 ? welem[13] : _GEN_7182; // @[Execute.scala 117:10]
  assign _GEN_7184 = 6'he == _T_644 ? welem[14] : _GEN_7183; // @[Execute.scala 117:10]
  assign _GEN_7185 = 6'hf == _T_644 ? welem[15] : _GEN_7184; // @[Execute.scala 117:10]
  assign _GEN_7186 = 6'h10 == _T_644 ? welem[16] : _GEN_7185; // @[Execute.scala 117:10]
  assign _GEN_7187 = 6'h11 == _T_644 ? welem[17] : _GEN_7186; // @[Execute.scala 117:10]
  assign _GEN_7188 = 6'h12 == _T_644 ? welem[18] : _GEN_7187; // @[Execute.scala 117:10]
  assign _GEN_7189 = 6'h13 == _T_644 ? welem[19] : _GEN_7188; // @[Execute.scala 117:10]
  assign _GEN_7190 = 6'h14 == _T_644 ? welem[20] : _GEN_7189; // @[Execute.scala 117:10]
  assign _GEN_7191 = 6'h15 == _T_644 ? welem[21] : _GEN_7190; // @[Execute.scala 117:10]
  assign _GEN_7192 = 6'h16 == _T_644 ? welem[22] : _GEN_7191; // @[Execute.scala 117:10]
  assign _GEN_7193 = 6'h17 == _T_644 ? welem[23] : _GEN_7192; // @[Execute.scala 117:10]
  assign _GEN_7194 = 6'h18 == _T_644 ? welem[24] : _GEN_7193; // @[Execute.scala 117:10]
  assign _GEN_7195 = 6'h19 == _T_644 ? welem[25] : _GEN_7194; // @[Execute.scala 117:10]
  assign _GEN_7196 = 6'h1a == _T_644 ? welem[26] : _GEN_7195; // @[Execute.scala 117:10]
  assign _GEN_7197 = 6'h1b == _T_644 ? welem[27] : _GEN_7196; // @[Execute.scala 117:10]
  assign _GEN_7198 = 6'h1c == _T_644 ? welem[28] : _GEN_7197; // @[Execute.scala 117:10]
  assign _GEN_7199 = 6'h1d == _T_644 ? welem[29] : _GEN_7198; // @[Execute.scala 117:10]
  assign _GEN_7200 = 6'h1e == _T_644 ? welem[30] : _GEN_7199; // @[Execute.scala 117:10]
  assign _GEN_7201 = 6'h1f == _T_644 ? welem[31] : _GEN_7200; // @[Execute.scala 117:10]
  assign _GEN_7202 = 6'h20 == _T_644 ? welem[32] : _GEN_7201; // @[Execute.scala 117:10]
  assign _GEN_7203 = 6'h21 == _T_644 ? welem[33] : _GEN_7202; // @[Execute.scala 117:10]
  assign _GEN_7204 = 6'h22 == _T_644 ? welem[34] : _GEN_7203; // @[Execute.scala 117:10]
  assign _GEN_7205 = 6'h23 == _T_644 ? welem[35] : _GEN_7204; // @[Execute.scala 117:10]
  assign _GEN_7206 = 6'h24 == _T_644 ? welem[36] : _GEN_7205; // @[Execute.scala 117:10]
  assign _GEN_7207 = 6'h25 == _T_644 ? welem[37] : _GEN_7206; // @[Execute.scala 117:10]
  assign _GEN_7208 = 6'h26 == _T_644 ? welem[38] : _GEN_7207; // @[Execute.scala 117:10]
  assign _GEN_7209 = 6'h27 == _T_644 ? welem[39] : _GEN_7208; // @[Execute.scala 117:10]
  assign _GEN_7210 = 6'h28 == _T_644 ? welem[40] : _GEN_7209; // @[Execute.scala 117:10]
  assign _GEN_7211 = 6'h29 == _T_644 ? welem[41] : _GEN_7210; // @[Execute.scala 117:10]
  assign _GEN_7212 = 6'h2a == _T_644 ? welem[42] : _GEN_7211; // @[Execute.scala 117:10]
  assign _GEN_7213 = 6'h2b == _T_644 ? welem[43] : _GEN_7212; // @[Execute.scala 117:10]
  assign _GEN_7214 = 6'h2c == _T_644 ? welem[44] : _GEN_7213; // @[Execute.scala 117:10]
  assign _GEN_7215 = 6'h2d == _T_644 ? welem[45] : _GEN_7214; // @[Execute.scala 117:10]
  assign _GEN_7216 = 6'h2e == _T_644 ? welem[46] : _GEN_7215; // @[Execute.scala 117:10]
  assign _GEN_7217 = 6'h2f == _T_644 ? welem[47] : _GEN_7216; // @[Execute.scala 117:10]
  assign _GEN_7218 = 6'h30 == _T_644 ? welem[48] : _GEN_7217; // @[Execute.scala 117:10]
  assign _GEN_7219 = 6'h31 == _T_644 ? welem[49] : _GEN_7218; // @[Execute.scala 117:10]
  assign _GEN_7220 = 6'h32 == _T_644 ? welem[50] : _GEN_7219; // @[Execute.scala 117:10]
  assign _GEN_7221 = 6'h33 == _T_644 ? welem[51] : _GEN_7220; // @[Execute.scala 117:10]
  assign _GEN_7222 = 6'h34 == _T_644 ? welem[52] : _GEN_7221; // @[Execute.scala 117:10]
  assign _GEN_7223 = 6'h35 == _T_644 ? welem[53] : _GEN_7222; // @[Execute.scala 117:10]
  assign _GEN_7224 = 6'h36 == _T_644 ? welem[54] : _GEN_7223; // @[Execute.scala 117:10]
  assign _GEN_7225 = 6'h37 == _T_644 ? welem[55] : _GEN_7224; // @[Execute.scala 117:10]
  assign _GEN_7226 = 6'h38 == _T_644 ? welem[56] : _GEN_7225; // @[Execute.scala 117:10]
  assign _GEN_7227 = 6'h39 == _T_644 ? welem[57] : _GEN_7226; // @[Execute.scala 117:10]
  assign _GEN_7228 = 6'h3a == _T_644 ? welem[58] : _GEN_7227; // @[Execute.scala 117:10]
  assign _GEN_7229 = 6'h3b == _T_644 ? welem[59] : _GEN_7228; // @[Execute.scala 117:10]
  assign _GEN_7230 = 6'h3c == _T_644 ? welem[60] : _GEN_7229; // @[Execute.scala 117:10]
  assign _GEN_7231 = 6'h3d == _T_644 ? welem[61] : _GEN_7230; // @[Execute.scala 117:10]
  assign _GEN_7232 = 6'h3e == _T_644 ? welem[62] : _GEN_7231; // @[Execute.scala 117:10]
  assign _GEN_7233 = 6'h3f == _T_644 ? welem[63] : _GEN_7232; // @[Execute.scala 117:10]
  assign _GEN_7235 = 6'h1 == _T_648 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7236 = 6'h2 == _T_648 ? welem[2] : _GEN_7235; // @[Execute.scala 117:10]
  assign _GEN_7237 = 6'h3 == _T_648 ? welem[3] : _GEN_7236; // @[Execute.scala 117:10]
  assign _GEN_7238 = 6'h4 == _T_648 ? welem[4] : _GEN_7237; // @[Execute.scala 117:10]
  assign _GEN_7239 = 6'h5 == _T_648 ? welem[5] : _GEN_7238; // @[Execute.scala 117:10]
  assign _GEN_7240 = 6'h6 == _T_648 ? welem[6] : _GEN_7239; // @[Execute.scala 117:10]
  assign _GEN_7241 = 6'h7 == _T_648 ? welem[7] : _GEN_7240; // @[Execute.scala 117:10]
  assign _GEN_7242 = 6'h8 == _T_648 ? welem[8] : _GEN_7241; // @[Execute.scala 117:10]
  assign _GEN_7243 = 6'h9 == _T_648 ? welem[9] : _GEN_7242; // @[Execute.scala 117:10]
  assign _GEN_7244 = 6'ha == _T_648 ? welem[10] : _GEN_7243; // @[Execute.scala 117:10]
  assign _GEN_7245 = 6'hb == _T_648 ? welem[11] : _GEN_7244; // @[Execute.scala 117:10]
  assign _GEN_7246 = 6'hc == _T_648 ? welem[12] : _GEN_7245; // @[Execute.scala 117:10]
  assign _GEN_7247 = 6'hd == _T_648 ? welem[13] : _GEN_7246; // @[Execute.scala 117:10]
  assign _GEN_7248 = 6'he == _T_648 ? welem[14] : _GEN_7247; // @[Execute.scala 117:10]
  assign _GEN_7249 = 6'hf == _T_648 ? welem[15] : _GEN_7248; // @[Execute.scala 117:10]
  assign _GEN_7250 = 6'h10 == _T_648 ? welem[16] : _GEN_7249; // @[Execute.scala 117:10]
  assign _GEN_7251 = 6'h11 == _T_648 ? welem[17] : _GEN_7250; // @[Execute.scala 117:10]
  assign _GEN_7252 = 6'h12 == _T_648 ? welem[18] : _GEN_7251; // @[Execute.scala 117:10]
  assign _GEN_7253 = 6'h13 == _T_648 ? welem[19] : _GEN_7252; // @[Execute.scala 117:10]
  assign _GEN_7254 = 6'h14 == _T_648 ? welem[20] : _GEN_7253; // @[Execute.scala 117:10]
  assign _GEN_7255 = 6'h15 == _T_648 ? welem[21] : _GEN_7254; // @[Execute.scala 117:10]
  assign _GEN_7256 = 6'h16 == _T_648 ? welem[22] : _GEN_7255; // @[Execute.scala 117:10]
  assign _GEN_7257 = 6'h17 == _T_648 ? welem[23] : _GEN_7256; // @[Execute.scala 117:10]
  assign _GEN_7258 = 6'h18 == _T_648 ? welem[24] : _GEN_7257; // @[Execute.scala 117:10]
  assign _GEN_7259 = 6'h19 == _T_648 ? welem[25] : _GEN_7258; // @[Execute.scala 117:10]
  assign _GEN_7260 = 6'h1a == _T_648 ? welem[26] : _GEN_7259; // @[Execute.scala 117:10]
  assign _GEN_7261 = 6'h1b == _T_648 ? welem[27] : _GEN_7260; // @[Execute.scala 117:10]
  assign _GEN_7262 = 6'h1c == _T_648 ? welem[28] : _GEN_7261; // @[Execute.scala 117:10]
  assign _GEN_7263 = 6'h1d == _T_648 ? welem[29] : _GEN_7262; // @[Execute.scala 117:10]
  assign _GEN_7264 = 6'h1e == _T_648 ? welem[30] : _GEN_7263; // @[Execute.scala 117:10]
  assign _GEN_7265 = 6'h1f == _T_648 ? welem[31] : _GEN_7264; // @[Execute.scala 117:10]
  assign _GEN_7266 = 6'h20 == _T_648 ? welem[32] : _GEN_7265; // @[Execute.scala 117:10]
  assign _GEN_7267 = 6'h21 == _T_648 ? welem[33] : _GEN_7266; // @[Execute.scala 117:10]
  assign _GEN_7268 = 6'h22 == _T_648 ? welem[34] : _GEN_7267; // @[Execute.scala 117:10]
  assign _GEN_7269 = 6'h23 == _T_648 ? welem[35] : _GEN_7268; // @[Execute.scala 117:10]
  assign _GEN_7270 = 6'h24 == _T_648 ? welem[36] : _GEN_7269; // @[Execute.scala 117:10]
  assign _GEN_7271 = 6'h25 == _T_648 ? welem[37] : _GEN_7270; // @[Execute.scala 117:10]
  assign _GEN_7272 = 6'h26 == _T_648 ? welem[38] : _GEN_7271; // @[Execute.scala 117:10]
  assign _GEN_7273 = 6'h27 == _T_648 ? welem[39] : _GEN_7272; // @[Execute.scala 117:10]
  assign _GEN_7274 = 6'h28 == _T_648 ? welem[40] : _GEN_7273; // @[Execute.scala 117:10]
  assign _GEN_7275 = 6'h29 == _T_648 ? welem[41] : _GEN_7274; // @[Execute.scala 117:10]
  assign _GEN_7276 = 6'h2a == _T_648 ? welem[42] : _GEN_7275; // @[Execute.scala 117:10]
  assign _GEN_7277 = 6'h2b == _T_648 ? welem[43] : _GEN_7276; // @[Execute.scala 117:10]
  assign _GEN_7278 = 6'h2c == _T_648 ? welem[44] : _GEN_7277; // @[Execute.scala 117:10]
  assign _GEN_7279 = 6'h2d == _T_648 ? welem[45] : _GEN_7278; // @[Execute.scala 117:10]
  assign _GEN_7280 = 6'h2e == _T_648 ? welem[46] : _GEN_7279; // @[Execute.scala 117:10]
  assign _GEN_7281 = 6'h2f == _T_648 ? welem[47] : _GEN_7280; // @[Execute.scala 117:10]
  assign _GEN_7282 = 6'h30 == _T_648 ? welem[48] : _GEN_7281; // @[Execute.scala 117:10]
  assign _GEN_7283 = 6'h31 == _T_648 ? welem[49] : _GEN_7282; // @[Execute.scala 117:10]
  assign _GEN_7284 = 6'h32 == _T_648 ? welem[50] : _GEN_7283; // @[Execute.scala 117:10]
  assign _GEN_7285 = 6'h33 == _T_648 ? welem[51] : _GEN_7284; // @[Execute.scala 117:10]
  assign _GEN_7286 = 6'h34 == _T_648 ? welem[52] : _GEN_7285; // @[Execute.scala 117:10]
  assign _GEN_7287 = 6'h35 == _T_648 ? welem[53] : _GEN_7286; // @[Execute.scala 117:10]
  assign _GEN_7288 = 6'h36 == _T_648 ? welem[54] : _GEN_7287; // @[Execute.scala 117:10]
  assign _GEN_7289 = 6'h37 == _T_648 ? welem[55] : _GEN_7288; // @[Execute.scala 117:10]
  assign _GEN_7290 = 6'h38 == _T_648 ? welem[56] : _GEN_7289; // @[Execute.scala 117:10]
  assign _GEN_7291 = 6'h39 == _T_648 ? welem[57] : _GEN_7290; // @[Execute.scala 117:10]
  assign _GEN_7292 = 6'h3a == _T_648 ? welem[58] : _GEN_7291; // @[Execute.scala 117:10]
  assign _GEN_7293 = 6'h3b == _T_648 ? welem[59] : _GEN_7292; // @[Execute.scala 117:10]
  assign _GEN_7294 = 6'h3c == _T_648 ? welem[60] : _GEN_7293; // @[Execute.scala 117:10]
  assign _GEN_7295 = 6'h3d == _T_648 ? welem[61] : _GEN_7294; // @[Execute.scala 117:10]
  assign _GEN_7296 = 6'h3e == _T_648 ? welem[62] : _GEN_7295; // @[Execute.scala 117:10]
  assign _GEN_7297 = 6'h3f == _T_648 ? welem[63] : _GEN_7296; // @[Execute.scala 117:10]
  assign _T_651 = _T_642 ? _GEN_7233 : _GEN_7297; // @[Execute.scala 117:10]
  assign _T_652 = r < 6'h8; // @[Execute.scala 117:15]
  assign _T_654 = r - 6'h8; // @[Execute.scala 117:37]
  assign _T_658 = 6'h38 + r; // @[Execute.scala 117:60]
  assign _GEN_7299 = 6'h1 == _T_654 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7300 = 6'h2 == _T_654 ? welem[2] : _GEN_7299; // @[Execute.scala 117:10]
  assign _GEN_7301 = 6'h3 == _T_654 ? welem[3] : _GEN_7300; // @[Execute.scala 117:10]
  assign _GEN_7302 = 6'h4 == _T_654 ? welem[4] : _GEN_7301; // @[Execute.scala 117:10]
  assign _GEN_7303 = 6'h5 == _T_654 ? welem[5] : _GEN_7302; // @[Execute.scala 117:10]
  assign _GEN_7304 = 6'h6 == _T_654 ? welem[6] : _GEN_7303; // @[Execute.scala 117:10]
  assign _GEN_7305 = 6'h7 == _T_654 ? welem[7] : _GEN_7304; // @[Execute.scala 117:10]
  assign _GEN_7306 = 6'h8 == _T_654 ? welem[8] : _GEN_7305; // @[Execute.scala 117:10]
  assign _GEN_7307 = 6'h9 == _T_654 ? welem[9] : _GEN_7306; // @[Execute.scala 117:10]
  assign _GEN_7308 = 6'ha == _T_654 ? welem[10] : _GEN_7307; // @[Execute.scala 117:10]
  assign _GEN_7309 = 6'hb == _T_654 ? welem[11] : _GEN_7308; // @[Execute.scala 117:10]
  assign _GEN_7310 = 6'hc == _T_654 ? welem[12] : _GEN_7309; // @[Execute.scala 117:10]
  assign _GEN_7311 = 6'hd == _T_654 ? welem[13] : _GEN_7310; // @[Execute.scala 117:10]
  assign _GEN_7312 = 6'he == _T_654 ? welem[14] : _GEN_7311; // @[Execute.scala 117:10]
  assign _GEN_7313 = 6'hf == _T_654 ? welem[15] : _GEN_7312; // @[Execute.scala 117:10]
  assign _GEN_7314 = 6'h10 == _T_654 ? welem[16] : _GEN_7313; // @[Execute.scala 117:10]
  assign _GEN_7315 = 6'h11 == _T_654 ? welem[17] : _GEN_7314; // @[Execute.scala 117:10]
  assign _GEN_7316 = 6'h12 == _T_654 ? welem[18] : _GEN_7315; // @[Execute.scala 117:10]
  assign _GEN_7317 = 6'h13 == _T_654 ? welem[19] : _GEN_7316; // @[Execute.scala 117:10]
  assign _GEN_7318 = 6'h14 == _T_654 ? welem[20] : _GEN_7317; // @[Execute.scala 117:10]
  assign _GEN_7319 = 6'h15 == _T_654 ? welem[21] : _GEN_7318; // @[Execute.scala 117:10]
  assign _GEN_7320 = 6'h16 == _T_654 ? welem[22] : _GEN_7319; // @[Execute.scala 117:10]
  assign _GEN_7321 = 6'h17 == _T_654 ? welem[23] : _GEN_7320; // @[Execute.scala 117:10]
  assign _GEN_7322 = 6'h18 == _T_654 ? welem[24] : _GEN_7321; // @[Execute.scala 117:10]
  assign _GEN_7323 = 6'h19 == _T_654 ? welem[25] : _GEN_7322; // @[Execute.scala 117:10]
  assign _GEN_7324 = 6'h1a == _T_654 ? welem[26] : _GEN_7323; // @[Execute.scala 117:10]
  assign _GEN_7325 = 6'h1b == _T_654 ? welem[27] : _GEN_7324; // @[Execute.scala 117:10]
  assign _GEN_7326 = 6'h1c == _T_654 ? welem[28] : _GEN_7325; // @[Execute.scala 117:10]
  assign _GEN_7327 = 6'h1d == _T_654 ? welem[29] : _GEN_7326; // @[Execute.scala 117:10]
  assign _GEN_7328 = 6'h1e == _T_654 ? welem[30] : _GEN_7327; // @[Execute.scala 117:10]
  assign _GEN_7329 = 6'h1f == _T_654 ? welem[31] : _GEN_7328; // @[Execute.scala 117:10]
  assign _GEN_7330 = 6'h20 == _T_654 ? welem[32] : _GEN_7329; // @[Execute.scala 117:10]
  assign _GEN_7331 = 6'h21 == _T_654 ? welem[33] : _GEN_7330; // @[Execute.scala 117:10]
  assign _GEN_7332 = 6'h22 == _T_654 ? welem[34] : _GEN_7331; // @[Execute.scala 117:10]
  assign _GEN_7333 = 6'h23 == _T_654 ? welem[35] : _GEN_7332; // @[Execute.scala 117:10]
  assign _GEN_7334 = 6'h24 == _T_654 ? welem[36] : _GEN_7333; // @[Execute.scala 117:10]
  assign _GEN_7335 = 6'h25 == _T_654 ? welem[37] : _GEN_7334; // @[Execute.scala 117:10]
  assign _GEN_7336 = 6'h26 == _T_654 ? welem[38] : _GEN_7335; // @[Execute.scala 117:10]
  assign _GEN_7337 = 6'h27 == _T_654 ? welem[39] : _GEN_7336; // @[Execute.scala 117:10]
  assign _GEN_7338 = 6'h28 == _T_654 ? welem[40] : _GEN_7337; // @[Execute.scala 117:10]
  assign _GEN_7339 = 6'h29 == _T_654 ? welem[41] : _GEN_7338; // @[Execute.scala 117:10]
  assign _GEN_7340 = 6'h2a == _T_654 ? welem[42] : _GEN_7339; // @[Execute.scala 117:10]
  assign _GEN_7341 = 6'h2b == _T_654 ? welem[43] : _GEN_7340; // @[Execute.scala 117:10]
  assign _GEN_7342 = 6'h2c == _T_654 ? welem[44] : _GEN_7341; // @[Execute.scala 117:10]
  assign _GEN_7343 = 6'h2d == _T_654 ? welem[45] : _GEN_7342; // @[Execute.scala 117:10]
  assign _GEN_7344 = 6'h2e == _T_654 ? welem[46] : _GEN_7343; // @[Execute.scala 117:10]
  assign _GEN_7345 = 6'h2f == _T_654 ? welem[47] : _GEN_7344; // @[Execute.scala 117:10]
  assign _GEN_7346 = 6'h30 == _T_654 ? welem[48] : _GEN_7345; // @[Execute.scala 117:10]
  assign _GEN_7347 = 6'h31 == _T_654 ? welem[49] : _GEN_7346; // @[Execute.scala 117:10]
  assign _GEN_7348 = 6'h32 == _T_654 ? welem[50] : _GEN_7347; // @[Execute.scala 117:10]
  assign _GEN_7349 = 6'h33 == _T_654 ? welem[51] : _GEN_7348; // @[Execute.scala 117:10]
  assign _GEN_7350 = 6'h34 == _T_654 ? welem[52] : _GEN_7349; // @[Execute.scala 117:10]
  assign _GEN_7351 = 6'h35 == _T_654 ? welem[53] : _GEN_7350; // @[Execute.scala 117:10]
  assign _GEN_7352 = 6'h36 == _T_654 ? welem[54] : _GEN_7351; // @[Execute.scala 117:10]
  assign _GEN_7353 = 6'h37 == _T_654 ? welem[55] : _GEN_7352; // @[Execute.scala 117:10]
  assign _GEN_7354 = 6'h38 == _T_654 ? welem[56] : _GEN_7353; // @[Execute.scala 117:10]
  assign _GEN_7355 = 6'h39 == _T_654 ? welem[57] : _GEN_7354; // @[Execute.scala 117:10]
  assign _GEN_7356 = 6'h3a == _T_654 ? welem[58] : _GEN_7355; // @[Execute.scala 117:10]
  assign _GEN_7357 = 6'h3b == _T_654 ? welem[59] : _GEN_7356; // @[Execute.scala 117:10]
  assign _GEN_7358 = 6'h3c == _T_654 ? welem[60] : _GEN_7357; // @[Execute.scala 117:10]
  assign _GEN_7359 = 6'h3d == _T_654 ? welem[61] : _GEN_7358; // @[Execute.scala 117:10]
  assign _GEN_7360 = 6'h3e == _T_654 ? welem[62] : _GEN_7359; // @[Execute.scala 117:10]
  assign _GEN_7361 = 6'h3f == _T_654 ? welem[63] : _GEN_7360; // @[Execute.scala 117:10]
  assign _GEN_7363 = 6'h1 == _T_658 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7364 = 6'h2 == _T_658 ? welem[2] : _GEN_7363; // @[Execute.scala 117:10]
  assign _GEN_7365 = 6'h3 == _T_658 ? welem[3] : _GEN_7364; // @[Execute.scala 117:10]
  assign _GEN_7366 = 6'h4 == _T_658 ? welem[4] : _GEN_7365; // @[Execute.scala 117:10]
  assign _GEN_7367 = 6'h5 == _T_658 ? welem[5] : _GEN_7366; // @[Execute.scala 117:10]
  assign _GEN_7368 = 6'h6 == _T_658 ? welem[6] : _GEN_7367; // @[Execute.scala 117:10]
  assign _GEN_7369 = 6'h7 == _T_658 ? welem[7] : _GEN_7368; // @[Execute.scala 117:10]
  assign _GEN_7370 = 6'h8 == _T_658 ? welem[8] : _GEN_7369; // @[Execute.scala 117:10]
  assign _GEN_7371 = 6'h9 == _T_658 ? welem[9] : _GEN_7370; // @[Execute.scala 117:10]
  assign _GEN_7372 = 6'ha == _T_658 ? welem[10] : _GEN_7371; // @[Execute.scala 117:10]
  assign _GEN_7373 = 6'hb == _T_658 ? welem[11] : _GEN_7372; // @[Execute.scala 117:10]
  assign _GEN_7374 = 6'hc == _T_658 ? welem[12] : _GEN_7373; // @[Execute.scala 117:10]
  assign _GEN_7375 = 6'hd == _T_658 ? welem[13] : _GEN_7374; // @[Execute.scala 117:10]
  assign _GEN_7376 = 6'he == _T_658 ? welem[14] : _GEN_7375; // @[Execute.scala 117:10]
  assign _GEN_7377 = 6'hf == _T_658 ? welem[15] : _GEN_7376; // @[Execute.scala 117:10]
  assign _GEN_7378 = 6'h10 == _T_658 ? welem[16] : _GEN_7377; // @[Execute.scala 117:10]
  assign _GEN_7379 = 6'h11 == _T_658 ? welem[17] : _GEN_7378; // @[Execute.scala 117:10]
  assign _GEN_7380 = 6'h12 == _T_658 ? welem[18] : _GEN_7379; // @[Execute.scala 117:10]
  assign _GEN_7381 = 6'h13 == _T_658 ? welem[19] : _GEN_7380; // @[Execute.scala 117:10]
  assign _GEN_7382 = 6'h14 == _T_658 ? welem[20] : _GEN_7381; // @[Execute.scala 117:10]
  assign _GEN_7383 = 6'h15 == _T_658 ? welem[21] : _GEN_7382; // @[Execute.scala 117:10]
  assign _GEN_7384 = 6'h16 == _T_658 ? welem[22] : _GEN_7383; // @[Execute.scala 117:10]
  assign _GEN_7385 = 6'h17 == _T_658 ? welem[23] : _GEN_7384; // @[Execute.scala 117:10]
  assign _GEN_7386 = 6'h18 == _T_658 ? welem[24] : _GEN_7385; // @[Execute.scala 117:10]
  assign _GEN_7387 = 6'h19 == _T_658 ? welem[25] : _GEN_7386; // @[Execute.scala 117:10]
  assign _GEN_7388 = 6'h1a == _T_658 ? welem[26] : _GEN_7387; // @[Execute.scala 117:10]
  assign _GEN_7389 = 6'h1b == _T_658 ? welem[27] : _GEN_7388; // @[Execute.scala 117:10]
  assign _GEN_7390 = 6'h1c == _T_658 ? welem[28] : _GEN_7389; // @[Execute.scala 117:10]
  assign _GEN_7391 = 6'h1d == _T_658 ? welem[29] : _GEN_7390; // @[Execute.scala 117:10]
  assign _GEN_7392 = 6'h1e == _T_658 ? welem[30] : _GEN_7391; // @[Execute.scala 117:10]
  assign _GEN_7393 = 6'h1f == _T_658 ? welem[31] : _GEN_7392; // @[Execute.scala 117:10]
  assign _GEN_7394 = 6'h20 == _T_658 ? welem[32] : _GEN_7393; // @[Execute.scala 117:10]
  assign _GEN_7395 = 6'h21 == _T_658 ? welem[33] : _GEN_7394; // @[Execute.scala 117:10]
  assign _GEN_7396 = 6'h22 == _T_658 ? welem[34] : _GEN_7395; // @[Execute.scala 117:10]
  assign _GEN_7397 = 6'h23 == _T_658 ? welem[35] : _GEN_7396; // @[Execute.scala 117:10]
  assign _GEN_7398 = 6'h24 == _T_658 ? welem[36] : _GEN_7397; // @[Execute.scala 117:10]
  assign _GEN_7399 = 6'h25 == _T_658 ? welem[37] : _GEN_7398; // @[Execute.scala 117:10]
  assign _GEN_7400 = 6'h26 == _T_658 ? welem[38] : _GEN_7399; // @[Execute.scala 117:10]
  assign _GEN_7401 = 6'h27 == _T_658 ? welem[39] : _GEN_7400; // @[Execute.scala 117:10]
  assign _GEN_7402 = 6'h28 == _T_658 ? welem[40] : _GEN_7401; // @[Execute.scala 117:10]
  assign _GEN_7403 = 6'h29 == _T_658 ? welem[41] : _GEN_7402; // @[Execute.scala 117:10]
  assign _GEN_7404 = 6'h2a == _T_658 ? welem[42] : _GEN_7403; // @[Execute.scala 117:10]
  assign _GEN_7405 = 6'h2b == _T_658 ? welem[43] : _GEN_7404; // @[Execute.scala 117:10]
  assign _GEN_7406 = 6'h2c == _T_658 ? welem[44] : _GEN_7405; // @[Execute.scala 117:10]
  assign _GEN_7407 = 6'h2d == _T_658 ? welem[45] : _GEN_7406; // @[Execute.scala 117:10]
  assign _GEN_7408 = 6'h2e == _T_658 ? welem[46] : _GEN_7407; // @[Execute.scala 117:10]
  assign _GEN_7409 = 6'h2f == _T_658 ? welem[47] : _GEN_7408; // @[Execute.scala 117:10]
  assign _GEN_7410 = 6'h30 == _T_658 ? welem[48] : _GEN_7409; // @[Execute.scala 117:10]
  assign _GEN_7411 = 6'h31 == _T_658 ? welem[49] : _GEN_7410; // @[Execute.scala 117:10]
  assign _GEN_7412 = 6'h32 == _T_658 ? welem[50] : _GEN_7411; // @[Execute.scala 117:10]
  assign _GEN_7413 = 6'h33 == _T_658 ? welem[51] : _GEN_7412; // @[Execute.scala 117:10]
  assign _GEN_7414 = 6'h34 == _T_658 ? welem[52] : _GEN_7413; // @[Execute.scala 117:10]
  assign _GEN_7415 = 6'h35 == _T_658 ? welem[53] : _GEN_7414; // @[Execute.scala 117:10]
  assign _GEN_7416 = 6'h36 == _T_658 ? welem[54] : _GEN_7415; // @[Execute.scala 117:10]
  assign _GEN_7417 = 6'h37 == _T_658 ? welem[55] : _GEN_7416; // @[Execute.scala 117:10]
  assign _GEN_7418 = 6'h38 == _T_658 ? welem[56] : _GEN_7417; // @[Execute.scala 117:10]
  assign _GEN_7419 = 6'h39 == _T_658 ? welem[57] : _GEN_7418; // @[Execute.scala 117:10]
  assign _GEN_7420 = 6'h3a == _T_658 ? welem[58] : _GEN_7419; // @[Execute.scala 117:10]
  assign _GEN_7421 = 6'h3b == _T_658 ? welem[59] : _GEN_7420; // @[Execute.scala 117:10]
  assign _GEN_7422 = 6'h3c == _T_658 ? welem[60] : _GEN_7421; // @[Execute.scala 117:10]
  assign _GEN_7423 = 6'h3d == _T_658 ? welem[61] : _GEN_7422; // @[Execute.scala 117:10]
  assign _GEN_7424 = 6'h3e == _T_658 ? welem[62] : _GEN_7423; // @[Execute.scala 117:10]
  assign _GEN_7425 = 6'h3f == _T_658 ? welem[63] : _GEN_7424; // @[Execute.scala 117:10]
  assign _T_661 = _T_652 ? _GEN_7361 : _GEN_7425; // @[Execute.scala 117:10]
  assign _T_662 = r < 6'h7; // @[Execute.scala 117:15]
  assign _T_664 = r - 6'h7; // @[Execute.scala 117:37]
  assign _T_668 = 6'h39 + r; // @[Execute.scala 117:60]
  assign _GEN_7427 = 6'h1 == _T_664 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7428 = 6'h2 == _T_664 ? welem[2] : _GEN_7427; // @[Execute.scala 117:10]
  assign _GEN_7429 = 6'h3 == _T_664 ? welem[3] : _GEN_7428; // @[Execute.scala 117:10]
  assign _GEN_7430 = 6'h4 == _T_664 ? welem[4] : _GEN_7429; // @[Execute.scala 117:10]
  assign _GEN_7431 = 6'h5 == _T_664 ? welem[5] : _GEN_7430; // @[Execute.scala 117:10]
  assign _GEN_7432 = 6'h6 == _T_664 ? welem[6] : _GEN_7431; // @[Execute.scala 117:10]
  assign _GEN_7433 = 6'h7 == _T_664 ? welem[7] : _GEN_7432; // @[Execute.scala 117:10]
  assign _GEN_7434 = 6'h8 == _T_664 ? welem[8] : _GEN_7433; // @[Execute.scala 117:10]
  assign _GEN_7435 = 6'h9 == _T_664 ? welem[9] : _GEN_7434; // @[Execute.scala 117:10]
  assign _GEN_7436 = 6'ha == _T_664 ? welem[10] : _GEN_7435; // @[Execute.scala 117:10]
  assign _GEN_7437 = 6'hb == _T_664 ? welem[11] : _GEN_7436; // @[Execute.scala 117:10]
  assign _GEN_7438 = 6'hc == _T_664 ? welem[12] : _GEN_7437; // @[Execute.scala 117:10]
  assign _GEN_7439 = 6'hd == _T_664 ? welem[13] : _GEN_7438; // @[Execute.scala 117:10]
  assign _GEN_7440 = 6'he == _T_664 ? welem[14] : _GEN_7439; // @[Execute.scala 117:10]
  assign _GEN_7441 = 6'hf == _T_664 ? welem[15] : _GEN_7440; // @[Execute.scala 117:10]
  assign _GEN_7442 = 6'h10 == _T_664 ? welem[16] : _GEN_7441; // @[Execute.scala 117:10]
  assign _GEN_7443 = 6'h11 == _T_664 ? welem[17] : _GEN_7442; // @[Execute.scala 117:10]
  assign _GEN_7444 = 6'h12 == _T_664 ? welem[18] : _GEN_7443; // @[Execute.scala 117:10]
  assign _GEN_7445 = 6'h13 == _T_664 ? welem[19] : _GEN_7444; // @[Execute.scala 117:10]
  assign _GEN_7446 = 6'h14 == _T_664 ? welem[20] : _GEN_7445; // @[Execute.scala 117:10]
  assign _GEN_7447 = 6'h15 == _T_664 ? welem[21] : _GEN_7446; // @[Execute.scala 117:10]
  assign _GEN_7448 = 6'h16 == _T_664 ? welem[22] : _GEN_7447; // @[Execute.scala 117:10]
  assign _GEN_7449 = 6'h17 == _T_664 ? welem[23] : _GEN_7448; // @[Execute.scala 117:10]
  assign _GEN_7450 = 6'h18 == _T_664 ? welem[24] : _GEN_7449; // @[Execute.scala 117:10]
  assign _GEN_7451 = 6'h19 == _T_664 ? welem[25] : _GEN_7450; // @[Execute.scala 117:10]
  assign _GEN_7452 = 6'h1a == _T_664 ? welem[26] : _GEN_7451; // @[Execute.scala 117:10]
  assign _GEN_7453 = 6'h1b == _T_664 ? welem[27] : _GEN_7452; // @[Execute.scala 117:10]
  assign _GEN_7454 = 6'h1c == _T_664 ? welem[28] : _GEN_7453; // @[Execute.scala 117:10]
  assign _GEN_7455 = 6'h1d == _T_664 ? welem[29] : _GEN_7454; // @[Execute.scala 117:10]
  assign _GEN_7456 = 6'h1e == _T_664 ? welem[30] : _GEN_7455; // @[Execute.scala 117:10]
  assign _GEN_7457 = 6'h1f == _T_664 ? welem[31] : _GEN_7456; // @[Execute.scala 117:10]
  assign _GEN_7458 = 6'h20 == _T_664 ? welem[32] : _GEN_7457; // @[Execute.scala 117:10]
  assign _GEN_7459 = 6'h21 == _T_664 ? welem[33] : _GEN_7458; // @[Execute.scala 117:10]
  assign _GEN_7460 = 6'h22 == _T_664 ? welem[34] : _GEN_7459; // @[Execute.scala 117:10]
  assign _GEN_7461 = 6'h23 == _T_664 ? welem[35] : _GEN_7460; // @[Execute.scala 117:10]
  assign _GEN_7462 = 6'h24 == _T_664 ? welem[36] : _GEN_7461; // @[Execute.scala 117:10]
  assign _GEN_7463 = 6'h25 == _T_664 ? welem[37] : _GEN_7462; // @[Execute.scala 117:10]
  assign _GEN_7464 = 6'h26 == _T_664 ? welem[38] : _GEN_7463; // @[Execute.scala 117:10]
  assign _GEN_7465 = 6'h27 == _T_664 ? welem[39] : _GEN_7464; // @[Execute.scala 117:10]
  assign _GEN_7466 = 6'h28 == _T_664 ? welem[40] : _GEN_7465; // @[Execute.scala 117:10]
  assign _GEN_7467 = 6'h29 == _T_664 ? welem[41] : _GEN_7466; // @[Execute.scala 117:10]
  assign _GEN_7468 = 6'h2a == _T_664 ? welem[42] : _GEN_7467; // @[Execute.scala 117:10]
  assign _GEN_7469 = 6'h2b == _T_664 ? welem[43] : _GEN_7468; // @[Execute.scala 117:10]
  assign _GEN_7470 = 6'h2c == _T_664 ? welem[44] : _GEN_7469; // @[Execute.scala 117:10]
  assign _GEN_7471 = 6'h2d == _T_664 ? welem[45] : _GEN_7470; // @[Execute.scala 117:10]
  assign _GEN_7472 = 6'h2e == _T_664 ? welem[46] : _GEN_7471; // @[Execute.scala 117:10]
  assign _GEN_7473 = 6'h2f == _T_664 ? welem[47] : _GEN_7472; // @[Execute.scala 117:10]
  assign _GEN_7474 = 6'h30 == _T_664 ? welem[48] : _GEN_7473; // @[Execute.scala 117:10]
  assign _GEN_7475 = 6'h31 == _T_664 ? welem[49] : _GEN_7474; // @[Execute.scala 117:10]
  assign _GEN_7476 = 6'h32 == _T_664 ? welem[50] : _GEN_7475; // @[Execute.scala 117:10]
  assign _GEN_7477 = 6'h33 == _T_664 ? welem[51] : _GEN_7476; // @[Execute.scala 117:10]
  assign _GEN_7478 = 6'h34 == _T_664 ? welem[52] : _GEN_7477; // @[Execute.scala 117:10]
  assign _GEN_7479 = 6'h35 == _T_664 ? welem[53] : _GEN_7478; // @[Execute.scala 117:10]
  assign _GEN_7480 = 6'h36 == _T_664 ? welem[54] : _GEN_7479; // @[Execute.scala 117:10]
  assign _GEN_7481 = 6'h37 == _T_664 ? welem[55] : _GEN_7480; // @[Execute.scala 117:10]
  assign _GEN_7482 = 6'h38 == _T_664 ? welem[56] : _GEN_7481; // @[Execute.scala 117:10]
  assign _GEN_7483 = 6'h39 == _T_664 ? welem[57] : _GEN_7482; // @[Execute.scala 117:10]
  assign _GEN_7484 = 6'h3a == _T_664 ? welem[58] : _GEN_7483; // @[Execute.scala 117:10]
  assign _GEN_7485 = 6'h3b == _T_664 ? welem[59] : _GEN_7484; // @[Execute.scala 117:10]
  assign _GEN_7486 = 6'h3c == _T_664 ? welem[60] : _GEN_7485; // @[Execute.scala 117:10]
  assign _GEN_7487 = 6'h3d == _T_664 ? welem[61] : _GEN_7486; // @[Execute.scala 117:10]
  assign _GEN_7488 = 6'h3e == _T_664 ? welem[62] : _GEN_7487; // @[Execute.scala 117:10]
  assign _GEN_7489 = 6'h3f == _T_664 ? welem[63] : _GEN_7488; // @[Execute.scala 117:10]
  assign _GEN_7491 = 6'h1 == _T_668 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7492 = 6'h2 == _T_668 ? welem[2] : _GEN_7491; // @[Execute.scala 117:10]
  assign _GEN_7493 = 6'h3 == _T_668 ? welem[3] : _GEN_7492; // @[Execute.scala 117:10]
  assign _GEN_7494 = 6'h4 == _T_668 ? welem[4] : _GEN_7493; // @[Execute.scala 117:10]
  assign _GEN_7495 = 6'h5 == _T_668 ? welem[5] : _GEN_7494; // @[Execute.scala 117:10]
  assign _GEN_7496 = 6'h6 == _T_668 ? welem[6] : _GEN_7495; // @[Execute.scala 117:10]
  assign _GEN_7497 = 6'h7 == _T_668 ? welem[7] : _GEN_7496; // @[Execute.scala 117:10]
  assign _GEN_7498 = 6'h8 == _T_668 ? welem[8] : _GEN_7497; // @[Execute.scala 117:10]
  assign _GEN_7499 = 6'h9 == _T_668 ? welem[9] : _GEN_7498; // @[Execute.scala 117:10]
  assign _GEN_7500 = 6'ha == _T_668 ? welem[10] : _GEN_7499; // @[Execute.scala 117:10]
  assign _GEN_7501 = 6'hb == _T_668 ? welem[11] : _GEN_7500; // @[Execute.scala 117:10]
  assign _GEN_7502 = 6'hc == _T_668 ? welem[12] : _GEN_7501; // @[Execute.scala 117:10]
  assign _GEN_7503 = 6'hd == _T_668 ? welem[13] : _GEN_7502; // @[Execute.scala 117:10]
  assign _GEN_7504 = 6'he == _T_668 ? welem[14] : _GEN_7503; // @[Execute.scala 117:10]
  assign _GEN_7505 = 6'hf == _T_668 ? welem[15] : _GEN_7504; // @[Execute.scala 117:10]
  assign _GEN_7506 = 6'h10 == _T_668 ? welem[16] : _GEN_7505; // @[Execute.scala 117:10]
  assign _GEN_7507 = 6'h11 == _T_668 ? welem[17] : _GEN_7506; // @[Execute.scala 117:10]
  assign _GEN_7508 = 6'h12 == _T_668 ? welem[18] : _GEN_7507; // @[Execute.scala 117:10]
  assign _GEN_7509 = 6'h13 == _T_668 ? welem[19] : _GEN_7508; // @[Execute.scala 117:10]
  assign _GEN_7510 = 6'h14 == _T_668 ? welem[20] : _GEN_7509; // @[Execute.scala 117:10]
  assign _GEN_7511 = 6'h15 == _T_668 ? welem[21] : _GEN_7510; // @[Execute.scala 117:10]
  assign _GEN_7512 = 6'h16 == _T_668 ? welem[22] : _GEN_7511; // @[Execute.scala 117:10]
  assign _GEN_7513 = 6'h17 == _T_668 ? welem[23] : _GEN_7512; // @[Execute.scala 117:10]
  assign _GEN_7514 = 6'h18 == _T_668 ? welem[24] : _GEN_7513; // @[Execute.scala 117:10]
  assign _GEN_7515 = 6'h19 == _T_668 ? welem[25] : _GEN_7514; // @[Execute.scala 117:10]
  assign _GEN_7516 = 6'h1a == _T_668 ? welem[26] : _GEN_7515; // @[Execute.scala 117:10]
  assign _GEN_7517 = 6'h1b == _T_668 ? welem[27] : _GEN_7516; // @[Execute.scala 117:10]
  assign _GEN_7518 = 6'h1c == _T_668 ? welem[28] : _GEN_7517; // @[Execute.scala 117:10]
  assign _GEN_7519 = 6'h1d == _T_668 ? welem[29] : _GEN_7518; // @[Execute.scala 117:10]
  assign _GEN_7520 = 6'h1e == _T_668 ? welem[30] : _GEN_7519; // @[Execute.scala 117:10]
  assign _GEN_7521 = 6'h1f == _T_668 ? welem[31] : _GEN_7520; // @[Execute.scala 117:10]
  assign _GEN_7522 = 6'h20 == _T_668 ? welem[32] : _GEN_7521; // @[Execute.scala 117:10]
  assign _GEN_7523 = 6'h21 == _T_668 ? welem[33] : _GEN_7522; // @[Execute.scala 117:10]
  assign _GEN_7524 = 6'h22 == _T_668 ? welem[34] : _GEN_7523; // @[Execute.scala 117:10]
  assign _GEN_7525 = 6'h23 == _T_668 ? welem[35] : _GEN_7524; // @[Execute.scala 117:10]
  assign _GEN_7526 = 6'h24 == _T_668 ? welem[36] : _GEN_7525; // @[Execute.scala 117:10]
  assign _GEN_7527 = 6'h25 == _T_668 ? welem[37] : _GEN_7526; // @[Execute.scala 117:10]
  assign _GEN_7528 = 6'h26 == _T_668 ? welem[38] : _GEN_7527; // @[Execute.scala 117:10]
  assign _GEN_7529 = 6'h27 == _T_668 ? welem[39] : _GEN_7528; // @[Execute.scala 117:10]
  assign _GEN_7530 = 6'h28 == _T_668 ? welem[40] : _GEN_7529; // @[Execute.scala 117:10]
  assign _GEN_7531 = 6'h29 == _T_668 ? welem[41] : _GEN_7530; // @[Execute.scala 117:10]
  assign _GEN_7532 = 6'h2a == _T_668 ? welem[42] : _GEN_7531; // @[Execute.scala 117:10]
  assign _GEN_7533 = 6'h2b == _T_668 ? welem[43] : _GEN_7532; // @[Execute.scala 117:10]
  assign _GEN_7534 = 6'h2c == _T_668 ? welem[44] : _GEN_7533; // @[Execute.scala 117:10]
  assign _GEN_7535 = 6'h2d == _T_668 ? welem[45] : _GEN_7534; // @[Execute.scala 117:10]
  assign _GEN_7536 = 6'h2e == _T_668 ? welem[46] : _GEN_7535; // @[Execute.scala 117:10]
  assign _GEN_7537 = 6'h2f == _T_668 ? welem[47] : _GEN_7536; // @[Execute.scala 117:10]
  assign _GEN_7538 = 6'h30 == _T_668 ? welem[48] : _GEN_7537; // @[Execute.scala 117:10]
  assign _GEN_7539 = 6'h31 == _T_668 ? welem[49] : _GEN_7538; // @[Execute.scala 117:10]
  assign _GEN_7540 = 6'h32 == _T_668 ? welem[50] : _GEN_7539; // @[Execute.scala 117:10]
  assign _GEN_7541 = 6'h33 == _T_668 ? welem[51] : _GEN_7540; // @[Execute.scala 117:10]
  assign _GEN_7542 = 6'h34 == _T_668 ? welem[52] : _GEN_7541; // @[Execute.scala 117:10]
  assign _GEN_7543 = 6'h35 == _T_668 ? welem[53] : _GEN_7542; // @[Execute.scala 117:10]
  assign _GEN_7544 = 6'h36 == _T_668 ? welem[54] : _GEN_7543; // @[Execute.scala 117:10]
  assign _GEN_7545 = 6'h37 == _T_668 ? welem[55] : _GEN_7544; // @[Execute.scala 117:10]
  assign _GEN_7546 = 6'h38 == _T_668 ? welem[56] : _GEN_7545; // @[Execute.scala 117:10]
  assign _GEN_7547 = 6'h39 == _T_668 ? welem[57] : _GEN_7546; // @[Execute.scala 117:10]
  assign _GEN_7548 = 6'h3a == _T_668 ? welem[58] : _GEN_7547; // @[Execute.scala 117:10]
  assign _GEN_7549 = 6'h3b == _T_668 ? welem[59] : _GEN_7548; // @[Execute.scala 117:10]
  assign _GEN_7550 = 6'h3c == _T_668 ? welem[60] : _GEN_7549; // @[Execute.scala 117:10]
  assign _GEN_7551 = 6'h3d == _T_668 ? welem[61] : _GEN_7550; // @[Execute.scala 117:10]
  assign _GEN_7552 = 6'h3e == _T_668 ? welem[62] : _GEN_7551; // @[Execute.scala 117:10]
  assign _GEN_7553 = 6'h3f == _T_668 ? welem[63] : _GEN_7552; // @[Execute.scala 117:10]
  assign _T_671 = _T_662 ? _GEN_7489 : _GEN_7553; // @[Execute.scala 117:10]
  assign _T_672 = r < 6'h6; // @[Execute.scala 117:15]
  assign _T_674 = r - 6'h6; // @[Execute.scala 117:37]
  assign _T_678 = 6'h3a + r; // @[Execute.scala 117:60]
  assign _GEN_7555 = 6'h1 == _T_674 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7556 = 6'h2 == _T_674 ? welem[2] : _GEN_7555; // @[Execute.scala 117:10]
  assign _GEN_7557 = 6'h3 == _T_674 ? welem[3] : _GEN_7556; // @[Execute.scala 117:10]
  assign _GEN_7558 = 6'h4 == _T_674 ? welem[4] : _GEN_7557; // @[Execute.scala 117:10]
  assign _GEN_7559 = 6'h5 == _T_674 ? welem[5] : _GEN_7558; // @[Execute.scala 117:10]
  assign _GEN_7560 = 6'h6 == _T_674 ? welem[6] : _GEN_7559; // @[Execute.scala 117:10]
  assign _GEN_7561 = 6'h7 == _T_674 ? welem[7] : _GEN_7560; // @[Execute.scala 117:10]
  assign _GEN_7562 = 6'h8 == _T_674 ? welem[8] : _GEN_7561; // @[Execute.scala 117:10]
  assign _GEN_7563 = 6'h9 == _T_674 ? welem[9] : _GEN_7562; // @[Execute.scala 117:10]
  assign _GEN_7564 = 6'ha == _T_674 ? welem[10] : _GEN_7563; // @[Execute.scala 117:10]
  assign _GEN_7565 = 6'hb == _T_674 ? welem[11] : _GEN_7564; // @[Execute.scala 117:10]
  assign _GEN_7566 = 6'hc == _T_674 ? welem[12] : _GEN_7565; // @[Execute.scala 117:10]
  assign _GEN_7567 = 6'hd == _T_674 ? welem[13] : _GEN_7566; // @[Execute.scala 117:10]
  assign _GEN_7568 = 6'he == _T_674 ? welem[14] : _GEN_7567; // @[Execute.scala 117:10]
  assign _GEN_7569 = 6'hf == _T_674 ? welem[15] : _GEN_7568; // @[Execute.scala 117:10]
  assign _GEN_7570 = 6'h10 == _T_674 ? welem[16] : _GEN_7569; // @[Execute.scala 117:10]
  assign _GEN_7571 = 6'h11 == _T_674 ? welem[17] : _GEN_7570; // @[Execute.scala 117:10]
  assign _GEN_7572 = 6'h12 == _T_674 ? welem[18] : _GEN_7571; // @[Execute.scala 117:10]
  assign _GEN_7573 = 6'h13 == _T_674 ? welem[19] : _GEN_7572; // @[Execute.scala 117:10]
  assign _GEN_7574 = 6'h14 == _T_674 ? welem[20] : _GEN_7573; // @[Execute.scala 117:10]
  assign _GEN_7575 = 6'h15 == _T_674 ? welem[21] : _GEN_7574; // @[Execute.scala 117:10]
  assign _GEN_7576 = 6'h16 == _T_674 ? welem[22] : _GEN_7575; // @[Execute.scala 117:10]
  assign _GEN_7577 = 6'h17 == _T_674 ? welem[23] : _GEN_7576; // @[Execute.scala 117:10]
  assign _GEN_7578 = 6'h18 == _T_674 ? welem[24] : _GEN_7577; // @[Execute.scala 117:10]
  assign _GEN_7579 = 6'h19 == _T_674 ? welem[25] : _GEN_7578; // @[Execute.scala 117:10]
  assign _GEN_7580 = 6'h1a == _T_674 ? welem[26] : _GEN_7579; // @[Execute.scala 117:10]
  assign _GEN_7581 = 6'h1b == _T_674 ? welem[27] : _GEN_7580; // @[Execute.scala 117:10]
  assign _GEN_7582 = 6'h1c == _T_674 ? welem[28] : _GEN_7581; // @[Execute.scala 117:10]
  assign _GEN_7583 = 6'h1d == _T_674 ? welem[29] : _GEN_7582; // @[Execute.scala 117:10]
  assign _GEN_7584 = 6'h1e == _T_674 ? welem[30] : _GEN_7583; // @[Execute.scala 117:10]
  assign _GEN_7585 = 6'h1f == _T_674 ? welem[31] : _GEN_7584; // @[Execute.scala 117:10]
  assign _GEN_7586 = 6'h20 == _T_674 ? welem[32] : _GEN_7585; // @[Execute.scala 117:10]
  assign _GEN_7587 = 6'h21 == _T_674 ? welem[33] : _GEN_7586; // @[Execute.scala 117:10]
  assign _GEN_7588 = 6'h22 == _T_674 ? welem[34] : _GEN_7587; // @[Execute.scala 117:10]
  assign _GEN_7589 = 6'h23 == _T_674 ? welem[35] : _GEN_7588; // @[Execute.scala 117:10]
  assign _GEN_7590 = 6'h24 == _T_674 ? welem[36] : _GEN_7589; // @[Execute.scala 117:10]
  assign _GEN_7591 = 6'h25 == _T_674 ? welem[37] : _GEN_7590; // @[Execute.scala 117:10]
  assign _GEN_7592 = 6'h26 == _T_674 ? welem[38] : _GEN_7591; // @[Execute.scala 117:10]
  assign _GEN_7593 = 6'h27 == _T_674 ? welem[39] : _GEN_7592; // @[Execute.scala 117:10]
  assign _GEN_7594 = 6'h28 == _T_674 ? welem[40] : _GEN_7593; // @[Execute.scala 117:10]
  assign _GEN_7595 = 6'h29 == _T_674 ? welem[41] : _GEN_7594; // @[Execute.scala 117:10]
  assign _GEN_7596 = 6'h2a == _T_674 ? welem[42] : _GEN_7595; // @[Execute.scala 117:10]
  assign _GEN_7597 = 6'h2b == _T_674 ? welem[43] : _GEN_7596; // @[Execute.scala 117:10]
  assign _GEN_7598 = 6'h2c == _T_674 ? welem[44] : _GEN_7597; // @[Execute.scala 117:10]
  assign _GEN_7599 = 6'h2d == _T_674 ? welem[45] : _GEN_7598; // @[Execute.scala 117:10]
  assign _GEN_7600 = 6'h2e == _T_674 ? welem[46] : _GEN_7599; // @[Execute.scala 117:10]
  assign _GEN_7601 = 6'h2f == _T_674 ? welem[47] : _GEN_7600; // @[Execute.scala 117:10]
  assign _GEN_7602 = 6'h30 == _T_674 ? welem[48] : _GEN_7601; // @[Execute.scala 117:10]
  assign _GEN_7603 = 6'h31 == _T_674 ? welem[49] : _GEN_7602; // @[Execute.scala 117:10]
  assign _GEN_7604 = 6'h32 == _T_674 ? welem[50] : _GEN_7603; // @[Execute.scala 117:10]
  assign _GEN_7605 = 6'h33 == _T_674 ? welem[51] : _GEN_7604; // @[Execute.scala 117:10]
  assign _GEN_7606 = 6'h34 == _T_674 ? welem[52] : _GEN_7605; // @[Execute.scala 117:10]
  assign _GEN_7607 = 6'h35 == _T_674 ? welem[53] : _GEN_7606; // @[Execute.scala 117:10]
  assign _GEN_7608 = 6'h36 == _T_674 ? welem[54] : _GEN_7607; // @[Execute.scala 117:10]
  assign _GEN_7609 = 6'h37 == _T_674 ? welem[55] : _GEN_7608; // @[Execute.scala 117:10]
  assign _GEN_7610 = 6'h38 == _T_674 ? welem[56] : _GEN_7609; // @[Execute.scala 117:10]
  assign _GEN_7611 = 6'h39 == _T_674 ? welem[57] : _GEN_7610; // @[Execute.scala 117:10]
  assign _GEN_7612 = 6'h3a == _T_674 ? welem[58] : _GEN_7611; // @[Execute.scala 117:10]
  assign _GEN_7613 = 6'h3b == _T_674 ? welem[59] : _GEN_7612; // @[Execute.scala 117:10]
  assign _GEN_7614 = 6'h3c == _T_674 ? welem[60] : _GEN_7613; // @[Execute.scala 117:10]
  assign _GEN_7615 = 6'h3d == _T_674 ? welem[61] : _GEN_7614; // @[Execute.scala 117:10]
  assign _GEN_7616 = 6'h3e == _T_674 ? welem[62] : _GEN_7615; // @[Execute.scala 117:10]
  assign _GEN_7617 = 6'h3f == _T_674 ? welem[63] : _GEN_7616; // @[Execute.scala 117:10]
  assign _GEN_7619 = 6'h1 == _T_678 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7620 = 6'h2 == _T_678 ? welem[2] : _GEN_7619; // @[Execute.scala 117:10]
  assign _GEN_7621 = 6'h3 == _T_678 ? welem[3] : _GEN_7620; // @[Execute.scala 117:10]
  assign _GEN_7622 = 6'h4 == _T_678 ? welem[4] : _GEN_7621; // @[Execute.scala 117:10]
  assign _GEN_7623 = 6'h5 == _T_678 ? welem[5] : _GEN_7622; // @[Execute.scala 117:10]
  assign _GEN_7624 = 6'h6 == _T_678 ? welem[6] : _GEN_7623; // @[Execute.scala 117:10]
  assign _GEN_7625 = 6'h7 == _T_678 ? welem[7] : _GEN_7624; // @[Execute.scala 117:10]
  assign _GEN_7626 = 6'h8 == _T_678 ? welem[8] : _GEN_7625; // @[Execute.scala 117:10]
  assign _GEN_7627 = 6'h9 == _T_678 ? welem[9] : _GEN_7626; // @[Execute.scala 117:10]
  assign _GEN_7628 = 6'ha == _T_678 ? welem[10] : _GEN_7627; // @[Execute.scala 117:10]
  assign _GEN_7629 = 6'hb == _T_678 ? welem[11] : _GEN_7628; // @[Execute.scala 117:10]
  assign _GEN_7630 = 6'hc == _T_678 ? welem[12] : _GEN_7629; // @[Execute.scala 117:10]
  assign _GEN_7631 = 6'hd == _T_678 ? welem[13] : _GEN_7630; // @[Execute.scala 117:10]
  assign _GEN_7632 = 6'he == _T_678 ? welem[14] : _GEN_7631; // @[Execute.scala 117:10]
  assign _GEN_7633 = 6'hf == _T_678 ? welem[15] : _GEN_7632; // @[Execute.scala 117:10]
  assign _GEN_7634 = 6'h10 == _T_678 ? welem[16] : _GEN_7633; // @[Execute.scala 117:10]
  assign _GEN_7635 = 6'h11 == _T_678 ? welem[17] : _GEN_7634; // @[Execute.scala 117:10]
  assign _GEN_7636 = 6'h12 == _T_678 ? welem[18] : _GEN_7635; // @[Execute.scala 117:10]
  assign _GEN_7637 = 6'h13 == _T_678 ? welem[19] : _GEN_7636; // @[Execute.scala 117:10]
  assign _GEN_7638 = 6'h14 == _T_678 ? welem[20] : _GEN_7637; // @[Execute.scala 117:10]
  assign _GEN_7639 = 6'h15 == _T_678 ? welem[21] : _GEN_7638; // @[Execute.scala 117:10]
  assign _GEN_7640 = 6'h16 == _T_678 ? welem[22] : _GEN_7639; // @[Execute.scala 117:10]
  assign _GEN_7641 = 6'h17 == _T_678 ? welem[23] : _GEN_7640; // @[Execute.scala 117:10]
  assign _GEN_7642 = 6'h18 == _T_678 ? welem[24] : _GEN_7641; // @[Execute.scala 117:10]
  assign _GEN_7643 = 6'h19 == _T_678 ? welem[25] : _GEN_7642; // @[Execute.scala 117:10]
  assign _GEN_7644 = 6'h1a == _T_678 ? welem[26] : _GEN_7643; // @[Execute.scala 117:10]
  assign _GEN_7645 = 6'h1b == _T_678 ? welem[27] : _GEN_7644; // @[Execute.scala 117:10]
  assign _GEN_7646 = 6'h1c == _T_678 ? welem[28] : _GEN_7645; // @[Execute.scala 117:10]
  assign _GEN_7647 = 6'h1d == _T_678 ? welem[29] : _GEN_7646; // @[Execute.scala 117:10]
  assign _GEN_7648 = 6'h1e == _T_678 ? welem[30] : _GEN_7647; // @[Execute.scala 117:10]
  assign _GEN_7649 = 6'h1f == _T_678 ? welem[31] : _GEN_7648; // @[Execute.scala 117:10]
  assign _GEN_7650 = 6'h20 == _T_678 ? welem[32] : _GEN_7649; // @[Execute.scala 117:10]
  assign _GEN_7651 = 6'h21 == _T_678 ? welem[33] : _GEN_7650; // @[Execute.scala 117:10]
  assign _GEN_7652 = 6'h22 == _T_678 ? welem[34] : _GEN_7651; // @[Execute.scala 117:10]
  assign _GEN_7653 = 6'h23 == _T_678 ? welem[35] : _GEN_7652; // @[Execute.scala 117:10]
  assign _GEN_7654 = 6'h24 == _T_678 ? welem[36] : _GEN_7653; // @[Execute.scala 117:10]
  assign _GEN_7655 = 6'h25 == _T_678 ? welem[37] : _GEN_7654; // @[Execute.scala 117:10]
  assign _GEN_7656 = 6'h26 == _T_678 ? welem[38] : _GEN_7655; // @[Execute.scala 117:10]
  assign _GEN_7657 = 6'h27 == _T_678 ? welem[39] : _GEN_7656; // @[Execute.scala 117:10]
  assign _GEN_7658 = 6'h28 == _T_678 ? welem[40] : _GEN_7657; // @[Execute.scala 117:10]
  assign _GEN_7659 = 6'h29 == _T_678 ? welem[41] : _GEN_7658; // @[Execute.scala 117:10]
  assign _GEN_7660 = 6'h2a == _T_678 ? welem[42] : _GEN_7659; // @[Execute.scala 117:10]
  assign _GEN_7661 = 6'h2b == _T_678 ? welem[43] : _GEN_7660; // @[Execute.scala 117:10]
  assign _GEN_7662 = 6'h2c == _T_678 ? welem[44] : _GEN_7661; // @[Execute.scala 117:10]
  assign _GEN_7663 = 6'h2d == _T_678 ? welem[45] : _GEN_7662; // @[Execute.scala 117:10]
  assign _GEN_7664 = 6'h2e == _T_678 ? welem[46] : _GEN_7663; // @[Execute.scala 117:10]
  assign _GEN_7665 = 6'h2f == _T_678 ? welem[47] : _GEN_7664; // @[Execute.scala 117:10]
  assign _GEN_7666 = 6'h30 == _T_678 ? welem[48] : _GEN_7665; // @[Execute.scala 117:10]
  assign _GEN_7667 = 6'h31 == _T_678 ? welem[49] : _GEN_7666; // @[Execute.scala 117:10]
  assign _GEN_7668 = 6'h32 == _T_678 ? welem[50] : _GEN_7667; // @[Execute.scala 117:10]
  assign _GEN_7669 = 6'h33 == _T_678 ? welem[51] : _GEN_7668; // @[Execute.scala 117:10]
  assign _GEN_7670 = 6'h34 == _T_678 ? welem[52] : _GEN_7669; // @[Execute.scala 117:10]
  assign _GEN_7671 = 6'h35 == _T_678 ? welem[53] : _GEN_7670; // @[Execute.scala 117:10]
  assign _GEN_7672 = 6'h36 == _T_678 ? welem[54] : _GEN_7671; // @[Execute.scala 117:10]
  assign _GEN_7673 = 6'h37 == _T_678 ? welem[55] : _GEN_7672; // @[Execute.scala 117:10]
  assign _GEN_7674 = 6'h38 == _T_678 ? welem[56] : _GEN_7673; // @[Execute.scala 117:10]
  assign _GEN_7675 = 6'h39 == _T_678 ? welem[57] : _GEN_7674; // @[Execute.scala 117:10]
  assign _GEN_7676 = 6'h3a == _T_678 ? welem[58] : _GEN_7675; // @[Execute.scala 117:10]
  assign _GEN_7677 = 6'h3b == _T_678 ? welem[59] : _GEN_7676; // @[Execute.scala 117:10]
  assign _GEN_7678 = 6'h3c == _T_678 ? welem[60] : _GEN_7677; // @[Execute.scala 117:10]
  assign _GEN_7679 = 6'h3d == _T_678 ? welem[61] : _GEN_7678; // @[Execute.scala 117:10]
  assign _GEN_7680 = 6'h3e == _T_678 ? welem[62] : _GEN_7679; // @[Execute.scala 117:10]
  assign _GEN_7681 = 6'h3f == _T_678 ? welem[63] : _GEN_7680; // @[Execute.scala 117:10]
  assign _T_681 = _T_672 ? _GEN_7617 : _GEN_7681; // @[Execute.scala 117:10]
  assign _T_682 = r < 6'h5; // @[Execute.scala 117:15]
  assign _T_684 = r - 6'h5; // @[Execute.scala 117:37]
  assign _T_688 = 6'h3b + r; // @[Execute.scala 117:60]
  assign _GEN_7683 = 6'h1 == _T_684 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7684 = 6'h2 == _T_684 ? welem[2] : _GEN_7683; // @[Execute.scala 117:10]
  assign _GEN_7685 = 6'h3 == _T_684 ? welem[3] : _GEN_7684; // @[Execute.scala 117:10]
  assign _GEN_7686 = 6'h4 == _T_684 ? welem[4] : _GEN_7685; // @[Execute.scala 117:10]
  assign _GEN_7687 = 6'h5 == _T_684 ? welem[5] : _GEN_7686; // @[Execute.scala 117:10]
  assign _GEN_7688 = 6'h6 == _T_684 ? welem[6] : _GEN_7687; // @[Execute.scala 117:10]
  assign _GEN_7689 = 6'h7 == _T_684 ? welem[7] : _GEN_7688; // @[Execute.scala 117:10]
  assign _GEN_7690 = 6'h8 == _T_684 ? welem[8] : _GEN_7689; // @[Execute.scala 117:10]
  assign _GEN_7691 = 6'h9 == _T_684 ? welem[9] : _GEN_7690; // @[Execute.scala 117:10]
  assign _GEN_7692 = 6'ha == _T_684 ? welem[10] : _GEN_7691; // @[Execute.scala 117:10]
  assign _GEN_7693 = 6'hb == _T_684 ? welem[11] : _GEN_7692; // @[Execute.scala 117:10]
  assign _GEN_7694 = 6'hc == _T_684 ? welem[12] : _GEN_7693; // @[Execute.scala 117:10]
  assign _GEN_7695 = 6'hd == _T_684 ? welem[13] : _GEN_7694; // @[Execute.scala 117:10]
  assign _GEN_7696 = 6'he == _T_684 ? welem[14] : _GEN_7695; // @[Execute.scala 117:10]
  assign _GEN_7697 = 6'hf == _T_684 ? welem[15] : _GEN_7696; // @[Execute.scala 117:10]
  assign _GEN_7698 = 6'h10 == _T_684 ? welem[16] : _GEN_7697; // @[Execute.scala 117:10]
  assign _GEN_7699 = 6'h11 == _T_684 ? welem[17] : _GEN_7698; // @[Execute.scala 117:10]
  assign _GEN_7700 = 6'h12 == _T_684 ? welem[18] : _GEN_7699; // @[Execute.scala 117:10]
  assign _GEN_7701 = 6'h13 == _T_684 ? welem[19] : _GEN_7700; // @[Execute.scala 117:10]
  assign _GEN_7702 = 6'h14 == _T_684 ? welem[20] : _GEN_7701; // @[Execute.scala 117:10]
  assign _GEN_7703 = 6'h15 == _T_684 ? welem[21] : _GEN_7702; // @[Execute.scala 117:10]
  assign _GEN_7704 = 6'h16 == _T_684 ? welem[22] : _GEN_7703; // @[Execute.scala 117:10]
  assign _GEN_7705 = 6'h17 == _T_684 ? welem[23] : _GEN_7704; // @[Execute.scala 117:10]
  assign _GEN_7706 = 6'h18 == _T_684 ? welem[24] : _GEN_7705; // @[Execute.scala 117:10]
  assign _GEN_7707 = 6'h19 == _T_684 ? welem[25] : _GEN_7706; // @[Execute.scala 117:10]
  assign _GEN_7708 = 6'h1a == _T_684 ? welem[26] : _GEN_7707; // @[Execute.scala 117:10]
  assign _GEN_7709 = 6'h1b == _T_684 ? welem[27] : _GEN_7708; // @[Execute.scala 117:10]
  assign _GEN_7710 = 6'h1c == _T_684 ? welem[28] : _GEN_7709; // @[Execute.scala 117:10]
  assign _GEN_7711 = 6'h1d == _T_684 ? welem[29] : _GEN_7710; // @[Execute.scala 117:10]
  assign _GEN_7712 = 6'h1e == _T_684 ? welem[30] : _GEN_7711; // @[Execute.scala 117:10]
  assign _GEN_7713 = 6'h1f == _T_684 ? welem[31] : _GEN_7712; // @[Execute.scala 117:10]
  assign _GEN_7714 = 6'h20 == _T_684 ? welem[32] : _GEN_7713; // @[Execute.scala 117:10]
  assign _GEN_7715 = 6'h21 == _T_684 ? welem[33] : _GEN_7714; // @[Execute.scala 117:10]
  assign _GEN_7716 = 6'h22 == _T_684 ? welem[34] : _GEN_7715; // @[Execute.scala 117:10]
  assign _GEN_7717 = 6'h23 == _T_684 ? welem[35] : _GEN_7716; // @[Execute.scala 117:10]
  assign _GEN_7718 = 6'h24 == _T_684 ? welem[36] : _GEN_7717; // @[Execute.scala 117:10]
  assign _GEN_7719 = 6'h25 == _T_684 ? welem[37] : _GEN_7718; // @[Execute.scala 117:10]
  assign _GEN_7720 = 6'h26 == _T_684 ? welem[38] : _GEN_7719; // @[Execute.scala 117:10]
  assign _GEN_7721 = 6'h27 == _T_684 ? welem[39] : _GEN_7720; // @[Execute.scala 117:10]
  assign _GEN_7722 = 6'h28 == _T_684 ? welem[40] : _GEN_7721; // @[Execute.scala 117:10]
  assign _GEN_7723 = 6'h29 == _T_684 ? welem[41] : _GEN_7722; // @[Execute.scala 117:10]
  assign _GEN_7724 = 6'h2a == _T_684 ? welem[42] : _GEN_7723; // @[Execute.scala 117:10]
  assign _GEN_7725 = 6'h2b == _T_684 ? welem[43] : _GEN_7724; // @[Execute.scala 117:10]
  assign _GEN_7726 = 6'h2c == _T_684 ? welem[44] : _GEN_7725; // @[Execute.scala 117:10]
  assign _GEN_7727 = 6'h2d == _T_684 ? welem[45] : _GEN_7726; // @[Execute.scala 117:10]
  assign _GEN_7728 = 6'h2e == _T_684 ? welem[46] : _GEN_7727; // @[Execute.scala 117:10]
  assign _GEN_7729 = 6'h2f == _T_684 ? welem[47] : _GEN_7728; // @[Execute.scala 117:10]
  assign _GEN_7730 = 6'h30 == _T_684 ? welem[48] : _GEN_7729; // @[Execute.scala 117:10]
  assign _GEN_7731 = 6'h31 == _T_684 ? welem[49] : _GEN_7730; // @[Execute.scala 117:10]
  assign _GEN_7732 = 6'h32 == _T_684 ? welem[50] : _GEN_7731; // @[Execute.scala 117:10]
  assign _GEN_7733 = 6'h33 == _T_684 ? welem[51] : _GEN_7732; // @[Execute.scala 117:10]
  assign _GEN_7734 = 6'h34 == _T_684 ? welem[52] : _GEN_7733; // @[Execute.scala 117:10]
  assign _GEN_7735 = 6'h35 == _T_684 ? welem[53] : _GEN_7734; // @[Execute.scala 117:10]
  assign _GEN_7736 = 6'h36 == _T_684 ? welem[54] : _GEN_7735; // @[Execute.scala 117:10]
  assign _GEN_7737 = 6'h37 == _T_684 ? welem[55] : _GEN_7736; // @[Execute.scala 117:10]
  assign _GEN_7738 = 6'h38 == _T_684 ? welem[56] : _GEN_7737; // @[Execute.scala 117:10]
  assign _GEN_7739 = 6'h39 == _T_684 ? welem[57] : _GEN_7738; // @[Execute.scala 117:10]
  assign _GEN_7740 = 6'h3a == _T_684 ? welem[58] : _GEN_7739; // @[Execute.scala 117:10]
  assign _GEN_7741 = 6'h3b == _T_684 ? welem[59] : _GEN_7740; // @[Execute.scala 117:10]
  assign _GEN_7742 = 6'h3c == _T_684 ? welem[60] : _GEN_7741; // @[Execute.scala 117:10]
  assign _GEN_7743 = 6'h3d == _T_684 ? welem[61] : _GEN_7742; // @[Execute.scala 117:10]
  assign _GEN_7744 = 6'h3e == _T_684 ? welem[62] : _GEN_7743; // @[Execute.scala 117:10]
  assign _GEN_7745 = 6'h3f == _T_684 ? welem[63] : _GEN_7744; // @[Execute.scala 117:10]
  assign _GEN_7747 = 6'h1 == _T_688 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7748 = 6'h2 == _T_688 ? welem[2] : _GEN_7747; // @[Execute.scala 117:10]
  assign _GEN_7749 = 6'h3 == _T_688 ? welem[3] : _GEN_7748; // @[Execute.scala 117:10]
  assign _GEN_7750 = 6'h4 == _T_688 ? welem[4] : _GEN_7749; // @[Execute.scala 117:10]
  assign _GEN_7751 = 6'h5 == _T_688 ? welem[5] : _GEN_7750; // @[Execute.scala 117:10]
  assign _GEN_7752 = 6'h6 == _T_688 ? welem[6] : _GEN_7751; // @[Execute.scala 117:10]
  assign _GEN_7753 = 6'h7 == _T_688 ? welem[7] : _GEN_7752; // @[Execute.scala 117:10]
  assign _GEN_7754 = 6'h8 == _T_688 ? welem[8] : _GEN_7753; // @[Execute.scala 117:10]
  assign _GEN_7755 = 6'h9 == _T_688 ? welem[9] : _GEN_7754; // @[Execute.scala 117:10]
  assign _GEN_7756 = 6'ha == _T_688 ? welem[10] : _GEN_7755; // @[Execute.scala 117:10]
  assign _GEN_7757 = 6'hb == _T_688 ? welem[11] : _GEN_7756; // @[Execute.scala 117:10]
  assign _GEN_7758 = 6'hc == _T_688 ? welem[12] : _GEN_7757; // @[Execute.scala 117:10]
  assign _GEN_7759 = 6'hd == _T_688 ? welem[13] : _GEN_7758; // @[Execute.scala 117:10]
  assign _GEN_7760 = 6'he == _T_688 ? welem[14] : _GEN_7759; // @[Execute.scala 117:10]
  assign _GEN_7761 = 6'hf == _T_688 ? welem[15] : _GEN_7760; // @[Execute.scala 117:10]
  assign _GEN_7762 = 6'h10 == _T_688 ? welem[16] : _GEN_7761; // @[Execute.scala 117:10]
  assign _GEN_7763 = 6'h11 == _T_688 ? welem[17] : _GEN_7762; // @[Execute.scala 117:10]
  assign _GEN_7764 = 6'h12 == _T_688 ? welem[18] : _GEN_7763; // @[Execute.scala 117:10]
  assign _GEN_7765 = 6'h13 == _T_688 ? welem[19] : _GEN_7764; // @[Execute.scala 117:10]
  assign _GEN_7766 = 6'h14 == _T_688 ? welem[20] : _GEN_7765; // @[Execute.scala 117:10]
  assign _GEN_7767 = 6'h15 == _T_688 ? welem[21] : _GEN_7766; // @[Execute.scala 117:10]
  assign _GEN_7768 = 6'h16 == _T_688 ? welem[22] : _GEN_7767; // @[Execute.scala 117:10]
  assign _GEN_7769 = 6'h17 == _T_688 ? welem[23] : _GEN_7768; // @[Execute.scala 117:10]
  assign _GEN_7770 = 6'h18 == _T_688 ? welem[24] : _GEN_7769; // @[Execute.scala 117:10]
  assign _GEN_7771 = 6'h19 == _T_688 ? welem[25] : _GEN_7770; // @[Execute.scala 117:10]
  assign _GEN_7772 = 6'h1a == _T_688 ? welem[26] : _GEN_7771; // @[Execute.scala 117:10]
  assign _GEN_7773 = 6'h1b == _T_688 ? welem[27] : _GEN_7772; // @[Execute.scala 117:10]
  assign _GEN_7774 = 6'h1c == _T_688 ? welem[28] : _GEN_7773; // @[Execute.scala 117:10]
  assign _GEN_7775 = 6'h1d == _T_688 ? welem[29] : _GEN_7774; // @[Execute.scala 117:10]
  assign _GEN_7776 = 6'h1e == _T_688 ? welem[30] : _GEN_7775; // @[Execute.scala 117:10]
  assign _GEN_7777 = 6'h1f == _T_688 ? welem[31] : _GEN_7776; // @[Execute.scala 117:10]
  assign _GEN_7778 = 6'h20 == _T_688 ? welem[32] : _GEN_7777; // @[Execute.scala 117:10]
  assign _GEN_7779 = 6'h21 == _T_688 ? welem[33] : _GEN_7778; // @[Execute.scala 117:10]
  assign _GEN_7780 = 6'h22 == _T_688 ? welem[34] : _GEN_7779; // @[Execute.scala 117:10]
  assign _GEN_7781 = 6'h23 == _T_688 ? welem[35] : _GEN_7780; // @[Execute.scala 117:10]
  assign _GEN_7782 = 6'h24 == _T_688 ? welem[36] : _GEN_7781; // @[Execute.scala 117:10]
  assign _GEN_7783 = 6'h25 == _T_688 ? welem[37] : _GEN_7782; // @[Execute.scala 117:10]
  assign _GEN_7784 = 6'h26 == _T_688 ? welem[38] : _GEN_7783; // @[Execute.scala 117:10]
  assign _GEN_7785 = 6'h27 == _T_688 ? welem[39] : _GEN_7784; // @[Execute.scala 117:10]
  assign _GEN_7786 = 6'h28 == _T_688 ? welem[40] : _GEN_7785; // @[Execute.scala 117:10]
  assign _GEN_7787 = 6'h29 == _T_688 ? welem[41] : _GEN_7786; // @[Execute.scala 117:10]
  assign _GEN_7788 = 6'h2a == _T_688 ? welem[42] : _GEN_7787; // @[Execute.scala 117:10]
  assign _GEN_7789 = 6'h2b == _T_688 ? welem[43] : _GEN_7788; // @[Execute.scala 117:10]
  assign _GEN_7790 = 6'h2c == _T_688 ? welem[44] : _GEN_7789; // @[Execute.scala 117:10]
  assign _GEN_7791 = 6'h2d == _T_688 ? welem[45] : _GEN_7790; // @[Execute.scala 117:10]
  assign _GEN_7792 = 6'h2e == _T_688 ? welem[46] : _GEN_7791; // @[Execute.scala 117:10]
  assign _GEN_7793 = 6'h2f == _T_688 ? welem[47] : _GEN_7792; // @[Execute.scala 117:10]
  assign _GEN_7794 = 6'h30 == _T_688 ? welem[48] : _GEN_7793; // @[Execute.scala 117:10]
  assign _GEN_7795 = 6'h31 == _T_688 ? welem[49] : _GEN_7794; // @[Execute.scala 117:10]
  assign _GEN_7796 = 6'h32 == _T_688 ? welem[50] : _GEN_7795; // @[Execute.scala 117:10]
  assign _GEN_7797 = 6'h33 == _T_688 ? welem[51] : _GEN_7796; // @[Execute.scala 117:10]
  assign _GEN_7798 = 6'h34 == _T_688 ? welem[52] : _GEN_7797; // @[Execute.scala 117:10]
  assign _GEN_7799 = 6'h35 == _T_688 ? welem[53] : _GEN_7798; // @[Execute.scala 117:10]
  assign _GEN_7800 = 6'h36 == _T_688 ? welem[54] : _GEN_7799; // @[Execute.scala 117:10]
  assign _GEN_7801 = 6'h37 == _T_688 ? welem[55] : _GEN_7800; // @[Execute.scala 117:10]
  assign _GEN_7802 = 6'h38 == _T_688 ? welem[56] : _GEN_7801; // @[Execute.scala 117:10]
  assign _GEN_7803 = 6'h39 == _T_688 ? welem[57] : _GEN_7802; // @[Execute.scala 117:10]
  assign _GEN_7804 = 6'h3a == _T_688 ? welem[58] : _GEN_7803; // @[Execute.scala 117:10]
  assign _GEN_7805 = 6'h3b == _T_688 ? welem[59] : _GEN_7804; // @[Execute.scala 117:10]
  assign _GEN_7806 = 6'h3c == _T_688 ? welem[60] : _GEN_7805; // @[Execute.scala 117:10]
  assign _GEN_7807 = 6'h3d == _T_688 ? welem[61] : _GEN_7806; // @[Execute.scala 117:10]
  assign _GEN_7808 = 6'h3e == _T_688 ? welem[62] : _GEN_7807; // @[Execute.scala 117:10]
  assign _GEN_7809 = 6'h3f == _T_688 ? welem[63] : _GEN_7808; // @[Execute.scala 117:10]
  assign _T_691 = _T_682 ? _GEN_7745 : _GEN_7809; // @[Execute.scala 117:10]
  assign _T_692 = r < 6'h4; // @[Execute.scala 117:15]
  assign _T_694 = r - 6'h4; // @[Execute.scala 117:37]
  assign _T_698 = 6'h3c + r; // @[Execute.scala 117:60]
  assign _GEN_7811 = 6'h1 == _T_694 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7812 = 6'h2 == _T_694 ? welem[2] : _GEN_7811; // @[Execute.scala 117:10]
  assign _GEN_7813 = 6'h3 == _T_694 ? welem[3] : _GEN_7812; // @[Execute.scala 117:10]
  assign _GEN_7814 = 6'h4 == _T_694 ? welem[4] : _GEN_7813; // @[Execute.scala 117:10]
  assign _GEN_7815 = 6'h5 == _T_694 ? welem[5] : _GEN_7814; // @[Execute.scala 117:10]
  assign _GEN_7816 = 6'h6 == _T_694 ? welem[6] : _GEN_7815; // @[Execute.scala 117:10]
  assign _GEN_7817 = 6'h7 == _T_694 ? welem[7] : _GEN_7816; // @[Execute.scala 117:10]
  assign _GEN_7818 = 6'h8 == _T_694 ? welem[8] : _GEN_7817; // @[Execute.scala 117:10]
  assign _GEN_7819 = 6'h9 == _T_694 ? welem[9] : _GEN_7818; // @[Execute.scala 117:10]
  assign _GEN_7820 = 6'ha == _T_694 ? welem[10] : _GEN_7819; // @[Execute.scala 117:10]
  assign _GEN_7821 = 6'hb == _T_694 ? welem[11] : _GEN_7820; // @[Execute.scala 117:10]
  assign _GEN_7822 = 6'hc == _T_694 ? welem[12] : _GEN_7821; // @[Execute.scala 117:10]
  assign _GEN_7823 = 6'hd == _T_694 ? welem[13] : _GEN_7822; // @[Execute.scala 117:10]
  assign _GEN_7824 = 6'he == _T_694 ? welem[14] : _GEN_7823; // @[Execute.scala 117:10]
  assign _GEN_7825 = 6'hf == _T_694 ? welem[15] : _GEN_7824; // @[Execute.scala 117:10]
  assign _GEN_7826 = 6'h10 == _T_694 ? welem[16] : _GEN_7825; // @[Execute.scala 117:10]
  assign _GEN_7827 = 6'h11 == _T_694 ? welem[17] : _GEN_7826; // @[Execute.scala 117:10]
  assign _GEN_7828 = 6'h12 == _T_694 ? welem[18] : _GEN_7827; // @[Execute.scala 117:10]
  assign _GEN_7829 = 6'h13 == _T_694 ? welem[19] : _GEN_7828; // @[Execute.scala 117:10]
  assign _GEN_7830 = 6'h14 == _T_694 ? welem[20] : _GEN_7829; // @[Execute.scala 117:10]
  assign _GEN_7831 = 6'h15 == _T_694 ? welem[21] : _GEN_7830; // @[Execute.scala 117:10]
  assign _GEN_7832 = 6'h16 == _T_694 ? welem[22] : _GEN_7831; // @[Execute.scala 117:10]
  assign _GEN_7833 = 6'h17 == _T_694 ? welem[23] : _GEN_7832; // @[Execute.scala 117:10]
  assign _GEN_7834 = 6'h18 == _T_694 ? welem[24] : _GEN_7833; // @[Execute.scala 117:10]
  assign _GEN_7835 = 6'h19 == _T_694 ? welem[25] : _GEN_7834; // @[Execute.scala 117:10]
  assign _GEN_7836 = 6'h1a == _T_694 ? welem[26] : _GEN_7835; // @[Execute.scala 117:10]
  assign _GEN_7837 = 6'h1b == _T_694 ? welem[27] : _GEN_7836; // @[Execute.scala 117:10]
  assign _GEN_7838 = 6'h1c == _T_694 ? welem[28] : _GEN_7837; // @[Execute.scala 117:10]
  assign _GEN_7839 = 6'h1d == _T_694 ? welem[29] : _GEN_7838; // @[Execute.scala 117:10]
  assign _GEN_7840 = 6'h1e == _T_694 ? welem[30] : _GEN_7839; // @[Execute.scala 117:10]
  assign _GEN_7841 = 6'h1f == _T_694 ? welem[31] : _GEN_7840; // @[Execute.scala 117:10]
  assign _GEN_7842 = 6'h20 == _T_694 ? welem[32] : _GEN_7841; // @[Execute.scala 117:10]
  assign _GEN_7843 = 6'h21 == _T_694 ? welem[33] : _GEN_7842; // @[Execute.scala 117:10]
  assign _GEN_7844 = 6'h22 == _T_694 ? welem[34] : _GEN_7843; // @[Execute.scala 117:10]
  assign _GEN_7845 = 6'h23 == _T_694 ? welem[35] : _GEN_7844; // @[Execute.scala 117:10]
  assign _GEN_7846 = 6'h24 == _T_694 ? welem[36] : _GEN_7845; // @[Execute.scala 117:10]
  assign _GEN_7847 = 6'h25 == _T_694 ? welem[37] : _GEN_7846; // @[Execute.scala 117:10]
  assign _GEN_7848 = 6'h26 == _T_694 ? welem[38] : _GEN_7847; // @[Execute.scala 117:10]
  assign _GEN_7849 = 6'h27 == _T_694 ? welem[39] : _GEN_7848; // @[Execute.scala 117:10]
  assign _GEN_7850 = 6'h28 == _T_694 ? welem[40] : _GEN_7849; // @[Execute.scala 117:10]
  assign _GEN_7851 = 6'h29 == _T_694 ? welem[41] : _GEN_7850; // @[Execute.scala 117:10]
  assign _GEN_7852 = 6'h2a == _T_694 ? welem[42] : _GEN_7851; // @[Execute.scala 117:10]
  assign _GEN_7853 = 6'h2b == _T_694 ? welem[43] : _GEN_7852; // @[Execute.scala 117:10]
  assign _GEN_7854 = 6'h2c == _T_694 ? welem[44] : _GEN_7853; // @[Execute.scala 117:10]
  assign _GEN_7855 = 6'h2d == _T_694 ? welem[45] : _GEN_7854; // @[Execute.scala 117:10]
  assign _GEN_7856 = 6'h2e == _T_694 ? welem[46] : _GEN_7855; // @[Execute.scala 117:10]
  assign _GEN_7857 = 6'h2f == _T_694 ? welem[47] : _GEN_7856; // @[Execute.scala 117:10]
  assign _GEN_7858 = 6'h30 == _T_694 ? welem[48] : _GEN_7857; // @[Execute.scala 117:10]
  assign _GEN_7859 = 6'h31 == _T_694 ? welem[49] : _GEN_7858; // @[Execute.scala 117:10]
  assign _GEN_7860 = 6'h32 == _T_694 ? welem[50] : _GEN_7859; // @[Execute.scala 117:10]
  assign _GEN_7861 = 6'h33 == _T_694 ? welem[51] : _GEN_7860; // @[Execute.scala 117:10]
  assign _GEN_7862 = 6'h34 == _T_694 ? welem[52] : _GEN_7861; // @[Execute.scala 117:10]
  assign _GEN_7863 = 6'h35 == _T_694 ? welem[53] : _GEN_7862; // @[Execute.scala 117:10]
  assign _GEN_7864 = 6'h36 == _T_694 ? welem[54] : _GEN_7863; // @[Execute.scala 117:10]
  assign _GEN_7865 = 6'h37 == _T_694 ? welem[55] : _GEN_7864; // @[Execute.scala 117:10]
  assign _GEN_7866 = 6'h38 == _T_694 ? welem[56] : _GEN_7865; // @[Execute.scala 117:10]
  assign _GEN_7867 = 6'h39 == _T_694 ? welem[57] : _GEN_7866; // @[Execute.scala 117:10]
  assign _GEN_7868 = 6'h3a == _T_694 ? welem[58] : _GEN_7867; // @[Execute.scala 117:10]
  assign _GEN_7869 = 6'h3b == _T_694 ? welem[59] : _GEN_7868; // @[Execute.scala 117:10]
  assign _GEN_7870 = 6'h3c == _T_694 ? welem[60] : _GEN_7869; // @[Execute.scala 117:10]
  assign _GEN_7871 = 6'h3d == _T_694 ? welem[61] : _GEN_7870; // @[Execute.scala 117:10]
  assign _GEN_7872 = 6'h3e == _T_694 ? welem[62] : _GEN_7871; // @[Execute.scala 117:10]
  assign _GEN_7873 = 6'h3f == _T_694 ? welem[63] : _GEN_7872; // @[Execute.scala 117:10]
  assign _GEN_7875 = 6'h1 == _T_698 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7876 = 6'h2 == _T_698 ? welem[2] : _GEN_7875; // @[Execute.scala 117:10]
  assign _GEN_7877 = 6'h3 == _T_698 ? welem[3] : _GEN_7876; // @[Execute.scala 117:10]
  assign _GEN_7878 = 6'h4 == _T_698 ? welem[4] : _GEN_7877; // @[Execute.scala 117:10]
  assign _GEN_7879 = 6'h5 == _T_698 ? welem[5] : _GEN_7878; // @[Execute.scala 117:10]
  assign _GEN_7880 = 6'h6 == _T_698 ? welem[6] : _GEN_7879; // @[Execute.scala 117:10]
  assign _GEN_7881 = 6'h7 == _T_698 ? welem[7] : _GEN_7880; // @[Execute.scala 117:10]
  assign _GEN_7882 = 6'h8 == _T_698 ? welem[8] : _GEN_7881; // @[Execute.scala 117:10]
  assign _GEN_7883 = 6'h9 == _T_698 ? welem[9] : _GEN_7882; // @[Execute.scala 117:10]
  assign _GEN_7884 = 6'ha == _T_698 ? welem[10] : _GEN_7883; // @[Execute.scala 117:10]
  assign _GEN_7885 = 6'hb == _T_698 ? welem[11] : _GEN_7884; // @[Execute.scala 117:10]
  assign _GEN_7886 = 6'hc == _T_698 ? welem[12] : _GEN_7885; // @[Execute.scala 117:10]
  assign _GEN_7887 = 6'hd == _T_698 ? welem[13] : _GEN_7886; // @[Execute.scala 117:10]
  assign _GEN_7888 = 6'he == _T_698 ? welem[14] : _GEN_7887; // @[Execute.scala 117:10]
  assign _GEN_7889 = 6'hf == _T_698 ? welem[15] : _GEN_7888; // @[Execute.scala 117:10]
  assign _GEN_7890 = 6'h10 == _T_698 ? welem[16] : _GEN_7889; // @[Execute.scala 117:10]
  assign _GEN_7891 = 6'h11 == _T_698 ? welem[17] : _GEN_7890; // @[Execute.scala 117:10]
  assign _GEN_7892 = 6'h12 == _T_698 ? welem[18] : _GEN_7891; // @[Execute.scala 117:10]
  assign _GEN_7893 = 6'h13 == _T_698 ? welem[19] : _GEN_7892; // @[Execute.scala 117:10]
  assign _GEN_7894 = 6'h14 == _T_698 ? welem[20] : _GEN_7893; // @[Execute.scala 117:10]
  assign _GEN_7895 = 6'h15 == _T_698 ? welem[21] : _GEN_7894; // @[Execute.scala 117:10]
  assign _GEN_7896 = 6'h16 == _T_698 ? welem[22] : _GEN_7895; // @[Execute.scala 117:10]
  assign _GEN_7897 = 6'h17 == _T_698 ? welem[23] : _GEN_7896; // @[Execute.scala 117:10]
  assign _GEN_7898 = 6'h18 == _T_698 ? welem[24] : _GEN_7897; // @[Execute.scala 117:10]
  assign _GEN_7899 = 6'h19 == _T_698 ? welem[25] : _GEN_7898; // @[Execute.scala 117:10]
  assign _GEN_7900 = 6'h1a == _T_698 ? welem[26] : _GEN_7899; // @[Execute.scala 117:10]
  assign _GEN_7901 = 6'h1b == _T_698 ? welem[27] : _GEN_7900; // @[Execute.scala 117:10]
  assign _GEN_7902 = 6'h1c == _T_698 ? welem[28] : _GEN_7901; // @[Execute.scala 117:10]
  assign _GEN_7903 = 6'h1d == _T_698 ? welem[29] : _GEN_7902; // @[Execute.scala 117:10]
  assign _GEN_7904 = 6'h1e == _T_698 ? welem[30] : _GEN_7903; // @[Execute.scala 117:10]
  assign _GEN_7905 = 6'h1f == _T_698 ? welem[31] : _GEN_7904; // @[Execute.scala 117:10]
  assign _GEN_7906 = 6'h20 == _T_698 ? welem[32] : _GEN_7905; // @[Execute.scala 117:10]
  assign _GEN_7907 = 6'h21 == _T_698 ? welem[33] : _GEN_7906; // @[Execute.scala 117:10]
  assign _GEN_7908 = 6'h22 == _T_698 ? welem[34] : _GEN_7907; // @[Execute.scala 117:10]
  assign _GEN_7909 = 6'h23 == _T_698 ? welem[35] : _GEN_7908; // @[Execute.scala 117:10]
  assign _GEN_7910 = 6'h24 == _T_698 ? welem[36] : _GEN_7909; // @[Execute.scala 117:10]
  assign _GEN_7911 = 6'h25 == _T_698 ? welem[37] : _GEN_7910; // @[Execute.scala 117:10]
  assign _GEN_7912 = 6'h26 == _T_698 ? welem[38] : _GEN_7911; // @[Execute.scala 117:10]
  assign _GEN_7913 = 6'h27 == _T_698 ? welem[39] : _GEN_7912; // @[Execute.scala 117:10]
  assign _GEN_7914 = 6'h28 == _T_698 ? welem[40] : _GEN_7913; // @[Execute.scala 117:10]
  assign _GEN_7915 = 6'h29 == _T_698 ? welem[41] : _GEN_7914; // @[Execute.scala 117:10]
  assign _GEN_7916 = 6'h2a == _T_698 ? welem[42] : _GEN_7915; // @[Execute.scala 117:10]
  assign _GEN_7917 = 6'h2b == _T_698 ? welem[43] : _GEN_7916; // @[Execute.scala 117:10]
  assign _GEN_7918 = 6'h2c == _T_698 ? welem[44] : _GEN_7917; // @[Execute.scala 117:10]
  assign _GEN_7919 = 6'h2d == _T_698 ? welem[45] : _GEN_7918; // @[Execute.scala 117:10]
  assign _GEN_7920 = 6'h2e == _T_698 ? welem[46] : _GEN_7919; // @[Execute.scala 117:10]
  assign _GEN_7921 = 6'h2f == _T_698 ? welem[47] : _GEN_7920; // @[Execute.scala 117:10]
  assign _GEN_7922 = 6'h30 == _T_698 ? welem[48] : _GEN_7921; // @[Execute.scala 117:10]
  assign _GEN_7923 = 6'h31 == _T_698 ? welem[49] : _GEN_7922; // @[Execute.scala 117:10]
  assign _GEN_7924 = 6'h32 == _T_698 ? welem[50] : _GEN_7923; // @[Execute.scala 117:10]
  assign _GEN_7925 = 6'h33 == _T_698 ? welem[51] : _GEN_7924; // @[Execute.scala 117:10]
  assign _GEN_7926 = 6'h34 == _T_698 ? welem[52] : _GEN_7925; // @[Execute.scala 117:10]
  assign _GEN_7927 = 6'h35 == _T_698 ? welem[53] : _GEN_7926; // @[Execute.scala 117:10]
  assign _GEN_7928 = 6'h36 == _T_698 ? welem[54] : _GEN_7927; // @[Execute.scala 117:10]
  assign _GEN_7929 = 6'h37 == _T_698 ? welem[55] : _GEN_7928; // @[Execute.scala 117:10]
  assign _GEN_7930 = 6'h38 == _T_698 ? welem[56] : _GEN_7929; // @[Execute.scala 117:10]
  assign _GEN_7931 = 6'h39 == _T_698 ? welem[57] : _GEN_7930; // @[Execute.scala 117:10]
  assign _GEN_7932 = 6'h3a == _T_698 ? welem[58] : _GEN_7931; // @[Execute.scala 117:10]
  assign _GEN_7933 = 6'h3b == _T_698 ? welem[59] : _GEN_7932; // @[Execute.scala 117:10]
  assign _GEN_7934 = 6'h3c == _T_698 ? welem[60] : _GEN_7933; // @[Execute.scala 117:10]
  assign _GEN_7935 = 6'h3d == _T_698 ? welem[61] : _GEN_7934; // @[Execute.scala 117:10]
  assign _GEN_7936 = 6'h3e == _T_698 ? welem[62] : _GEN_7935; // @[Execute.scala 117:10]
  assign _GEN_7937 = 6'h3f == _T_698 ? welem[63] : _GEN_7936; // @[Execute.scala 117:10]
  assign _T_701 = _T_692 ? _GEN_7873 : _GEN_7937; // @[Execute.scala 117:10]
  assign _T_702 = r < 6'h3; // @[Execute.scala 117:15]
  assign _T_704 = r - 6'h3; // @[Execute.scala 117:37]
  assign _T_708 = 6'h3d + r; // @[Execute.scala 117:60]
  assign _GEN_7939 = 6'h1 == _T_704 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_7940 = 6'h2 == _T_704 ? welem[2] : _GEN_7939; // @[Execute.scala 117:10]
  assign _GEN_7941 = 6'h3 == _T_704 ? welem[3] : _GEN_7940; // @[Execute.scala 117:10]
  assign _GEN_7942 = 6'h4 == _T_704 ? welem[4] : _GEN_7941; // @[Execute.scala 117:10]
  assign _GEN_7943 = 6'h5 == _T_704 ? welem[5] : _GEN_7942; // @[Execute.scala 117:10]
  assign _GEN_7944 = 6'h6 == _T_704 ? welem[6] : _GEN_7943; // @[Execute.scala 117:10]
  assign _GEN_7945 = 6'h7 == _T_704 ? welem[7] : _GEN_7944; // @[Execute.scala 117:10]
  assign _GEN_7946 = 6'h8 == _T_704 ? welem[8] : _GEN_7945; // @[Execute.scala 117:10]
  assign _GEN_7947 = 6'h9 == _T_704 ? welem[9] : _GEN_7946; // @[Execute.scala 117:10]
  assign _GEN_7948 = 6'ha == _T_704 ? welem[10] : _GEN_7947; // @[Execute.scala 117:10]
  assign _GEN_7949 = 6'hb == _T_704 ? welem[11] : _GEN_7948; // @[Execute.scala 117:10]
  assign _GEN_7950 = 6'hc == _T_704 ? welem[12] : _GEN_7949; // @[Execute.scala 117:10]
  assign _GEN_7951 = 6'hd == _T_704 ? welem[13] : _GEN_7950; // @[Execute.scala 117:10]
  assign _GEN_7952 = 6'he == _T_704 ? welem[14] : _GEN_7951; // @[Execute.scala 117:10]
  assign _GEN_7953 = 6'hf == _T_704 ? welem[15] : _GEN_7952; // @[Execute.scala 117:10]
  assign _GEN_7954 = 6'h10 == _T_704 ? welem[16] : _GEN_7953; // @[Execute.scala 117:10]
  assign _GEN_7955 = 6'h11 == _T_704 ? welem[17] : _GEN_7954; // @[Execute.scala 117:10]
  assign _GEN_7956 = 6'h12 == _T_704 ? welem[18] : _GEN_7955; // @[Execute.scala 117:10]
  assign _GEN_7957 = 6'h13 == _T_704 ? welem[19] : _GEN_7956; // @[Execute.scala 117:10]
  assign _GEN_7958 = 6'h14 == _T_704 ? welem[20] : _GEN_7957; // @[Execute.scala 117:10]
  assign _GEN_7959 = 6'h15 == _T_704 ? welem[21] : _GEN_7958; // @[Execute.scala 117:10]
  assign _GEN_7960 = 6'h16 == _T_704 ? welem[22] : _GEN_7959; // @[Execute.scala 117:10]
  assign _GEN_7961 = 6'h17 == _T_704 ? welem[23] : _GEN_7960; // @[Execute.scala 117:10]
  assign _GEN_7962 = 6'h18 == _T_704 ? welem[24] : _GEN_7961; // @[Execute.scala 117:10]
  assign _GEN_7963 = 6'h19 == _T_704 ? welem[25] : _GEN_7962; // @[Execute.scala 117:10]
  assign _GEN_7964 = 6'h1a == _T_704 ? welem[26] : _GEN_7963; // @[Execute.scala 117:10]
  assign _GEN_7965 = 6'h1b == _T_704 ? welem[27] : _GEN_7964; // @[Execute.scala 117:10]
  assign _GEN_7966 = 6'h1c == _T_704 ? welem[28] : _GEN_7965; // @[Execute.scala 117:10]
  assign _GEN_7967 = 6'h1d == _T_704 ? welem[29] : _GEN_7966; // @[Execute.scala 117:10]
  assign _GEN_7968 = 6'h1e == _T_704 ? welem[30] : _GEN_7967; // @[Execute.scala 117:10]
  assign _GEN_7969 = 6'h1f == _T_704 ? welem[31] : _GEN_7968; // @[Execute.scala 117:10]
  assign _GEN_7970 = 6'h20 == _T_704 ? welem[32] : _GEN_7969; // @[Execute.scala 117:10]
  assign _GEN_7971 = 6'h21 == _T_704 ? welem[33] : _GEN_7970; // @[Execute.scala 117:10]
  assign _GEN_7972 = 6'h22 == _T_704 ? welem[34] : _GEN_7971; // @[Execute.scala 117:10]
  assign _GEN_7973 = 6'h23 == _T_704 ? welem[35] : _GEN_7972; // @[Execute.scala 117:10]
  assign _GEN_7974 = 6'h24 == _T_704 ? welem[36] : _GEN_7973; // @[Execute.scala 117:10]
  assign _GEN_7975 = 6'h25 == _T_704 ? welem[37] : _GEN_7974; // @[Execute.scala 117:10]
  assign _GEN_7976 = 6'h26 == _T_704 ? welem[38] : _GEN_7975; // @[Execute.scala 117:10]
  assign _GEN_7977 = 6'h27 == _T_704 ? welem[39] : _GEN_7976; // @[Execute.scala 117:10]
  assign _GEN_7978 = 6'h28 == _T_704 ? welem[40] : _GEN_7977; // @[Execute.scala 117:10]
  assign _GEN_7979 = 6'h29 == _T_704 ? welem[41] : _GEN_7978; // @[Execute.scala 117:10]
  assign _GEN_7980 = 6'h2a == _T_704 ? welem[42] : _GEN_7979; // @[Execute.scala 117:10]
  assign _GEN_7981 = 6'h2b == _T_704 ? welem[43] : _GEN_7980; // @[Execute.scala 117:10]
  assign _GEN_7982 = 6'h2c == _T_704 ? welem[44] : _GEN_7981; // @[Execute.scala 117:10]
  assign _GEN_7983 = 6'h2d == _T_704 ? welem[45] : _GEN_7982; // @[Execute.scala 117:10]
  assign _GEN_7984 = 6'h2e == _T_704 ? welem[46] : _GEN_7983; // @[Execute.scala 117:10]
  assign _GEN_7985 = 6'h2f == _T_704 ? welem[47] : _GEN_7984; // @[Execute.scala 117:10]
  assign _GEN_7986 = 6'h30 == _T_704 ? welem[48] : _GEN_7985; // @[Execute.scala 117:10]
  assign _GEN_7987 = 6'h31 == _T_704 ? welem[49] : _GEN_7986; // @[Execute.scala 117:10]
  assign _GEN_7988 = 6'h32 == _T_704 ? welem[50] : _GEN_7987; // @[Execute.scala 117:10]
  assign _GEN_7989 = 6'h33 == _T_704 ? welem[51] : _GEN_7988; // @[Execute.scala 117:10]
  assign _GEN_7990 = 6'h34 == _T_704 ? welem[52] : _GEN_7989; // @[Execute.scala 117:10]
  assign _GEN_7991 = 6'h35 == _T_704 ? welem[53] : _GEN_7990; // @[Execute.scala 117:10]
  assign _GEN_7992 = 6'h36 == _T_704 ? welem[54] : _GEN_7991; // @[Execute.scala 117:10]
  assign _GEN_7993 = 6'h37 == _T_704 ? welem[55] : _GEN_7992; // @[Execute.scala 117:10]
  assign _GEN_7994 = 6'h38 == _T_704 ? welem[56] : _GEN_7993; // @[Execute.scala 117:10]
  assign _GEN_7995 = 6'h39 == _T_704 ? welem[57] : _GEN_7994; // @[Execute.scala 117:10]
  assign _GEN_7996 = 6'h3a == _T_704 ? welem[58] : _GEN_7995; // @[Execute.scala 117:10]
  assign _GEN_7997 = 6'h3b == _T_704 ? welem[59] : _GEN_7996; // @[Execute.scala 117:10]
  assign _GEN_7998 = 6'h3c == _T_704 ? welem[60] : _GEN_7997; // @[Execute.scala 117:10]
  assign _GEN_7999 = 6'h3d == _T_704 ? welem[61] : _GEN_7998; // @[Execute.scala 117:10]
  assign _GEN_8000 = 6'h3e == _T_704 ? welem[62] : _GEN_7999; // @[Execute.scala 117:10]
  assign _GEN_8001 = 6'h3f == _T_704 ? welem[63] : _GEN_8000; // @[Execute.scala 117:10]
  assign _GEN_8003 = 6'h1 == _T_708 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8004 = 6'h2 == _T_708 ? welem[2] : _GEN_8003; // @[Execute.scala 117:10]
  assign _GEN_8005 = 6'h3 == _T_708 ? welem[3] : _GEN_8004; // @[Execute.scala 117:10]
  assign _GEN_8006 = 6'h4 == _T_708 ? welem[4] : _GEN_8005; // @[Execute.scala 117:10]
  assign _GEN_8007 = 6'h5 == _T_708 ? welem[5] : _GEN_8006; // @[Execute.scala 117:10]
  assign _GEN_8008 = 6'h6 == _T_708 ? welem[6] : _GEN_8007; // @[Execute.scala 117:10]
  assign _GEN_8009 = 6'h7 == _T_708 ? welem[7] : _GEN_8008; // @[Execute.scala 117:10]
  assign _GEN_8010 = 6'h8 == _T_708 ? welem[8] : _GEN_8009; // @[Execute.scala 117:10]
  assign _GEN_8011 = 6'h9 == _T_708 ? welem[9] : _GEN_8010; // @[Execute.scala 117:10]
  assign _GEN_8012 = 6'ha == _T_708 ? welem[10] : _GEN_8011; // @[Execute.scala 117:10]
  assign _GEN_8013 = 6'hb == _T_708 ? welem[11] : _GEN_8012; // @[Execute.scala 117:10]
  assign _GEN_8014 = 6'hc == _T_708 ? welem[12] : _GEN_8013; // @[Execute.scala 117:10]
  assign _GEN_8015 = 6'hd == _T_708 ? welem[13] : _GEN_8014; // @[Execute.scala 117:10]
  assign _GEN_8016 = 6'he == _T_708 ? welem[14] : _GEN_8015; // @[Execute.scala 117:10]
  assign _GEN_8017 = 6'hf == _T_708 ? welem[15] : _GEN_8016; // @[Execute.scala 117:10]
  assign _GEN_8018 = 6'h10 == _T_708 ? welem[16] : _GEN_8017; // @[Execute.scala 117:10]
  assign _GEN_8019 = 6'h11 == _T_708 ? welem[17] : _GEN_8018; // @[Execute.scala 117:10]
  assign _GEN_8020 = 6'h12 == _T_708 ? welem[18] : _GEN_8019; // @[Execute.scala 117:10]
  assign _GEN_8021 = 6'h13 == _T_708 ? welem[19] : _GEN_8020; // @[Execute.scala 117:10]
  assign _GEN_8022 = 6'h14 == _T_708 ? welem[20] : _GEN_8021; // @[Execute.scala 117:10]
  assign _GEN_8023 = 6'h15 == _T_708 ? welem[21] : _GEN_8022; // @[Execute.scala 117:10]
  assign _GEN_8024 = 6'h16 == _T_708 ? welem[22] : _GEN_8023; // @[Execute.scala 117:10]
  assign _GEN_8025 = 6'h17 == _T_708 ? welem[23] : _GEN_8024; // @[Execute.scala 117:10]
  assign _GEN_8026 = 6'h18 == _T_708 ? welem[24] : _GEN_8025; // @[Execute.scala 117:10]
  assign _GEN_8027 = 6'h19 == _T_708 ? welem[25] : _GEN_8026; // @[Execute.scala 117:10]
  assign _GEN_8028 = 6'h1a == _T_708 ? welem[26] : _GEN_8027; // @[Execute.scala 117:10]
  assign _GEN_8029 = 6'h1b == _T_708 ? welem[27] : _GEN_8028; // @[Execute.scala 117:10]
  assign _GEN_8030 = 6'h1c == _T_708 ? welem[28] : _GEN_8029; // @[Execute.scala 117:10]
  assign _GEN_8031 = 6'h1d == _T_708 ? welem[29] : _GEN_8030; // @[Execute.scala 117:10]
  assign _GEN_8032 = 6'h1e == _T_708 ? welem[30] : _GEN_8031; // @[Execute.scala 117:10]
  assign _GEN_8033 = 6'h1f == _T_708 ? welem[31] : _GEN_8032; // @[Execute.scala 117:10]
  assign _GEN_8034 = 6'h20 == _T_708 ? welem[32] : _GEN_8033; // @[Execute.scala 117:10]
  assign _GEN_8035 = 6'h21 == _T_708 ? welem[33] : _GEN_8034; // @[Execute.scala 117:10]
  assign _GEN_8036 = 6'h22 == _T_708 ? welem[34] : _GEN_8035; // @[Execute.scala 117:10]
  assign _GEN_8037 = 6'h23 == _T_708 ? welem[35] : _GEN_8036; // @[Execute.scala 117:10]
  assign _GEN_8038 = 6'h24 == _T_708 ? welem[36] : _GEN_8037; // @[Execute.scala 117:10]
  assign _GEN_8039 = 6'h25 == _T_708 ? welem[37] : _GEN_8038; // @[Execute.scala 117:10]
  assign _GEN_8040 = 6'h26 == _T_708 ? welem[38] : _GEN_8039; // @[Execute.scala 117:10]
  assign _GEN_8041 = 6'h27 == _T_708 ? welem[39] : _GEN_8040; // @[Execute.scala 117:10]
  assign _GEN_8042 = 6'h28 == _T_708 ? welem[40] : _GEN_8041; // @[Execute.scala 117:10]
  assign _GEN_8043 = 6'h29 == _T_708 ? welem[41] : _GEN_8042; // @[Execute.scala 117:10]
  assign _GEN_8044 = 6'h2a == _T_708 ? welem[42] : _GEN_8043; // @[Execute.scala 117:10]
  assign _GEN_8045 = 6'h2b == _T_708 ? welem[43] : _GEN_8044; // @[Execute.scala 117:10]
  assign _GEN_8046 = 6'h2c == _T_708 ? welem[44] : _GEN_8045; // @[Execute.scala 117:10]
  assign _GEN_8047 = 6'h2d == _T_708 ? welem[45] : _GEN_8046; // @[Execute.scala 117:10]
  assign _GEN_8048 = 6'h2e == _T_708 ? welem[46] : _GEN_8047; // @[Execute.scala 117:10]
  assign _GEN_8049 = 6'h2f == _T_708 ? welem[47] : _GEN_8048; // @[Execute.scala 117:10]
  assign _GEN_8050 = 6'h30 == _T_708 ? welem[48] : _GEN_8049; // @[Execute.scala 117:10]
  assign _GEN_8051 = 6'h31 == _T_708 ? welem[49] : _GEN_8050; // @[Execute.scala 117:10]
  assign _GEN_8052 = 6'h32 == _T_708 ? welem[50] : _GEN_8051; // @[Execute.scala 117:10]
  assign _GEN_8053 = 6'h33 == _T_708 ? welem[51] : _GEN_8052; // @[Execute.scala 117:10]
  assign _GEN_8054 = 6'h34 == _T_708 ? welem[52] : _GEN_8053; // @[Execute.scala 117:10]
  assign _GEN_8055 = 6'h35 == _T_708 ? welem[53] : _GEN_8054; // @[Execute.scala 117:10]
  assign _GEN_8056 = 6'h36 == _T_708 ? welem[54] : _GEN_8055; // @[Execute.scala 117:10]
  assign _GEN_8057 = 6'h37 == _T_708 ? welem[55] : _GEN_8056; // @[Execute.scala 117:10]
  assign _GEN_8058 = 6'h38 == _T_708 ? welem[56] : _GEN_8057; // @[Execute.scala 117:10]
  assign _GEN_8059 = 6'h39 == _T_708 ? welem[57] : _GEN_8058; // @[Execute.scala 117:10]
  assign _GEN_8060 = 6'h3a == _T_708 ? welem[58] : _GEN_8059; // @[Execute.scala 117:10]
  assign _GEN_8061 = 6'h3b == _T_708 ? welem[59] : _GEN_8060; // @[Execute.scala 117:10]
  assign _GEN_8062 = 6'h3c == _T_708 ? welem[60] : _GEN_8061; // @[Execute.scala 117:10]
  assign _GEN_8063 = 6'h3d == _T_708 ? welem[61] : _GEN_8062; // @[Execute.scala 117:10]
  assign _GEN_8064 = 6'h3e == _T_708 ? welem[62] : _GEN_8063; // @[Execute.scala 117:10]
  assign _GEN_8065 = 6'h3f == _T_708 ? welem[63] : _GEN_8064; // @[Execute.scala 117:10]
  assign _T_711 = _T_702 ? _GEN_8001 : _GEN_8065; // @[Execute.scala 117:10]
  assign _T_712 = r < 6'h2; // @[Execute.scala 117:15]
  assign _T_714 = r - 6'h2; // @[Execute.scala 117:37]
  assign _T_718 = 6'h3e + r; // @[Execute.scala 117:60]
  assign _GEN_8067 = 6'h1 == _T_714 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8068 = 6'h2 == _T_714 ? welem[2] : _GEN_8067; // @[Execute.scala 117:10]
  assign _GEN_8069 = 6'h3 == _T_714 ? welem[3] : _GEN_8068; // @[Execute.scala 117:10]
  assign _GEN_8070 = 6'h4 == _T_714 ? welem[4] : _GEN_8069; // @[Execute.scala 117:10]
  assign _GEN_8071 = 6'h5 == _T_714 ? welem[5] : _GEN_8070; // @[Execute.scala 117:10]
  assign _GEN_8072 = 6'h6 == _T_714 ? welem[6] : _GEN_8071; // @[Execute.scala 117:10]
  assign _GEN_8073 = 6'h7 == _T_714 ? welem[7] : _GEN_8072; // @[Execute.scala 117:10]
  assign _GEN_8074 = 6'h8 == _T_714 ? welem[8] : _GEN_8073; // @[Execute.scala 117:10]
  assign _GEN_8075 = 6'h9 == _T_714 ? welem[9] : _GEN_8074; // @[Execute.scala 117:10]
  assign _GEN_8076 = 6'ha == _T_714 ? welem[10] : _GEN_8075; // @[Execute.scala 117:10]
  assign _GEN_8077 = 6'hb == _T_714 ? welem[11] : _GEN_8076; // @[Execute.scala 117:10]
  assign _GEN_8078 = 6'hc == _T_714 ? welem[12] : _GEN_8077; // @[Execute.scala 117:10]
  assign _GEN_8079 = 6'hd == _T_714 ? welem[13] : _GEN_8078; // @[Execute.scala 117:10]
  assign _GEN_8080 = 6'he == _T_714 ? welem[14] : _GEN_8079; // @[Execute.scala 117:10]
  assign _GEN_8081 = 6'hf == _T_714 ? welem[15] : _GEN_8080; // @[Execute.scala 117:10]
  assign _GEN_8082 = 6'h10 == _T_714 ? welem[16] : _GEN_8081; // @[Execute.scala 117:10]
  assign _GEN_8083 = 6'h11 == _T_714 ? welem[17] : _GEN_8082; // @[Execute.scala 117:10]
  assign _GEN_8084 = 6'h12 == _T_714 ? welem[18] : _GEN_8083; // @[Execute.scala 117:10]
  assign _GEN_8085 = 6'h13 == _T_714 ? welem[19] : _GEN_8084; // @[Execute.scala 117:10]
  assign _GEN_8086 = 6'h14 == _T_714 ? welem[20] : _GEN_8085; // @[Execute.scala 117:10]
  assign _GEN_8087 = 6'h15 == _T_714 ? welem[21] : _GEN_8086; // @[Execute.scala 117:10]
  assign _GEN_8088 = 6'h16 == _T_714 ? welem[22] : _GEN_8087; // @[Execute.scala 117:10]
  assign _GEN_8089 = 6'h17 == _T_714 ? welem[23] : _GEN_8088; // @[Execute.scala 117:10]
  assign _GEN_8090 = 6'h18 == _T_714 ? welem[24] : _GEN_8089; // @[Execute.scala 117:10]
  assign _GEN_8091 = 6'h19 == _T_714 ? welem[25] : _GEN_8090; // @[Execute.scala 117:10]
  assign _GEN_8092 = 6'h1a == _T_714 ? welem[26] : _GEN_8091; // @[Execute.scala 117:10]
  assign _GEN_8093 = 6'h1b == _T_714 ? welem[27] : _GEN_8092; // @[Execute.scala 117:10]
  assign _GEN_8094 = 6'h1c == _T_714 ? welem[28] : _GEN_8093; // @[Execute.scala 117:10]
  assign _GEN_8095 = 6'h1d == _T_714 ? welem[29] : _GEN_8094; // @[Execute.scala 117:10]
  assign _GEN_8096 = 6'h1e == _T_714 ? welem[30] : _GEN_8095; // @[Execute.scala 117:10]
  assign _GEN_8097 = 6'h1f == _T_714 ? welem[31] : _GEN_8096; // @[Execute.scala 117:10]
  assign _GEN_8098 = 6'h20 == _T_714 ? welem[32] : _GEN_8097; // @[Execute.scala 117:10]
  assign _GEN_8099 = 6'h21 == _T_714 ? welem[33] : _GEN_8098; // @[Execute.scala 117:10]
  assign _GEN_8100 = 6'h22 == _T_714 ? welem[34] : _GEN_8099; // @[Execute.scala 117:10]
  assign _GEN_8101 = 6'h23 == _T_714 ? welem[35] : _GEN_8100; // @[Execute.scala 117:10]
  assign _GEN_8102 = 6'h24 == _T_714 ? welem[36] : _GEN_8101; // @[Execute.scala 117:10]
  assign _GEN_8103 = 6'h25 == _T_714 ? welem[37] : _GEN_8102; // @[Execute.scala 117:10]
  assign _GEN_8104 = 6'h26 == _T_714 ? welem[38] : _GEN_8103; // @[Execute.scala 117:10]
  assign _GEN_8105 = 6'h27 == _T_714 ? welem[39] : _GEN_8104; // @[Execute.scala 117:10]
  assign _GEN_8106 = 6'h28 == _T_714 ? welem[40] : _GEN_8105; // @[Execute.scala 117:10]
  assign _GEN_8107 = 6'h29 == _T_714 ? welem[41] : _GEN_8106; // @[Execute.scala 117:10]
  assign _GEN_8108 = 6'h2a == _T_714 ? welem[42] : _GEN_8107; // @[Execute.scala 117:10]
  assign _GEN_8109 = 6'h2b == _T_714 ? welem[43] : _GEN_8108; // @[Execute.scala 117:10]
  assign _GEN_8110 = 6'h2c == _T_714 ? welem[44] : _GEN_8109; // @[Execute.scala 117:10]
  assign _GEN_8111 = 6'h2d == _T_714 ? welem[45] : _GEN_8110; // @[Execute.scala 117:10]
  assign _GEN_8112 = 6'h2e == _T_714 ? welem[46] : _GEN_8111; // @[Execute.scala 117:10]
  assign _GEN_8113 = 6'h2f == _T_714 ? welem[47] : _GEN_8112; // @[Execute.scala 117:10]
  assign _GEN_8114 = 6'h30 == _T_714 ? welem[48] : _GEN_8113; // @[Execute.scala 117:10]
  assign _GEN_8115 = 6'h31 == _T_714 ? welem[49] : _GEN_8114; // @[Execute.scala 117:10]
  assign _GEN_8116 = 6'h32 == _T_714 ? welem[50] : _GEN_8115; // @[Execute.scala 117:10]
  assign _GEN_8117 = 6'h33 == _T_714 ? welem[51] : _GEN_8116; // @[Execute.scala 117:10]
  assign _GEN_8118 = 6'h34 == _T_714 ? welem[52] : _GEN_8117; // @[Execute.scala 117:10]
  assign _GEN_8119 = 6'h35 == _T_714 ? welem[53] : _GEN_8118; // @[Execute.scala 117:10]
  assign _GEN_8120 = 6'h36 == _T_714 ? welem[54] : _GEN_8119; // @[Execute.scala 117:10]
  assign _GEN_8121 = 6'h37 == _T_714 ? welem[55] : _GEN_8120; // @[Execute.scala 117:10]
  assign _GEN_8122 = 6'h38 == _T_714 ? welem[56] : _GEN_8121; // @[Execute.scala 117:10]
  assign _GEN_8123 = 6'h39 == _T_714 ? welem[57] : _GEN_8122; // @[Execute.scala 117:10]
  assign _GEN_8124 = 6'h3a == _T_714 ? welem[58] : _GEN_8123; // @[Execute.scala 117:10]
  assign _GEN_8125 = 6'h3b == _T_714 ? welem[59] : _GEN_8124; // @[Execute.scala 117:10]
  assign _GEN_8126 = 6'h3c == _T_714 ? welem[60] : _GEN_8125; // @[Execute.scala 117:10]
  assign _GEN_8127 = 6'h3d == _T_714 ? welem[61] : _GEN_8126; // @[Execute.scala 117:10]
  assign _GEN_8128 = 6'h3e == _T_714 ? welem[62] : _GEN_8127; // @[Execute.scala 117:10]
  assign _GEN_8129 = 6'h3f == _T_714 ? welem[63] : _GEN_8128; // @[Execute.scala 117:10]
  assign _GEN_8131 = 6'h1 == _T_718 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8132 = 6'h2 == _T_718 ? welem[2] : _GEN_8131; // @[Execute.scala 117:10]
  assign _GEN_8133 = 6'h3 == _T_718 ? welem[3] : _GEN_8132; // @[Execute.scala 117:10]
  assign _GEN_8134 = 6'h4 == _T_718 ? welem[4] : _GEN_8133; // @[Execute.scala 117:10]
  assign _GEN_8135 = 6'h5 == _T_718 ? welem[5] : _GEN_8134; // @[Execute.scala 117:10]
  assign _GEN_8136 = 6'h6 == _T_718 ? welem[6] : _GEN_8135; // @[Execute.scala 117:10]
  assign _GEN_8137 = 6'h7 == _T_718 ? welem[7] : _GEN_8136; // @[Execute.scala 117:10]
  assign _GEN_8138 = 6'h8 == _T_718 ? welem[8] : _GEN_8137; // @[Execute.scala 117:10]
  assign _GEN_8139 = 6'h9 == _T_718 ? welem[9] : _GEN_8138; // @[Execute.scala 117:10]
  assign _GEN_8140 = 6'ha == _T_718 ? welem[10] : _GEN_8139; // @[Execute.scala 117:10]
  assign _GEN_8141 = 6'hb == _T_718 ? welem[11] : _GEN_8140; // @[Execute.scala 117:10]
  assign _GEN_8142 = 6'hc == _T_718 ? welem[12] : _GEN_8141; // @[Execute.scala 117:10]
  assign _GEN_8143 = 6'hd == _T_718 ? welem[13] : _GEN_8142; // @[Execute.scala 117:10]
  assign _GEN_8144 = 6'he == _T_718 ? welem[14] : _GEN_8143; // @[Execute.scala 117:10]
  assign _GEN_8145 = 6'hf == _T_718 ? welem[15] : _GEN_8144; // @[Execute.scala 117:10]
  assign _GEN_8146 = 6'h10 == _T_718 ? welem[16] : _GEN_8145; // @[Execute.scala 117:10]
  assign _GEN_8147 = 6'h11 == _T_718 ? welem[17] : _GEN_8146; // @[Execute.scala 117:10]
  assign _GEN_8148 = 6'h12 == _T_718 ? welem[18] : _GEN_8147; // @[Execute.scala 117:10]
  assign _GEN_8149 = 6'h13 == _T_718 ? welem[19] : _GEN_8148; // @[Execute.scala 117:10]
  assign _GEN_8150 = 6'h14 == _T_718 ? welem[20] : _GEN_8149; // @[Execute.scala 117:10]
  assign _GEN_8151 = 6'h15 == _T_718 ? welem[21] : _GEN_8150; // @[Execute.scala 117:10]
  assign _GEN_8152 = 6'h16 == _T_718 ? welem[22] : _GEN_8151; // @[Execute.scala 117:10]
  assign _GEN_8153 = 6'h17 == _T_718 ? welem[23] : _GEN_8152; // @[Execute.scala 117:10]
  assign _GEN_8154 = 6'h18 == _T_718 ? welem[24] : _GEN_8153; // @[Execute.scala 117:10]
  assign _GEN_8155 = 6'h19 == _T_718 ? welem[25] : _GEN_8154; // @[Execute.scala 117:10]
  assign _GEN_8156 = 6'h1a == _T_718 ? welem[26] : _GEN_8155; // @[Execute.scala 117:10]
  assign _GEN_8157 = 6'h1b == _T_718 ? welem[27] : _GEN_8156; // @[Execute.scala 117:10]
  assign _GEN_8158 = 6'h1c == _T_718 ? welem[28] : _GEN_8157; // @[Execute.scala 117:10]
  assign _GEN_8159 = 6'h1d == _T_718 ? welem[29] : _GEN_8158; // @[Execute.scala 117:10]
  assign _GEN_8160 = 6'h1e == _T_718 ? welem[30] : _GEN_8159; // @[Execute.scala 117:10]
  assign _GEN_8161 = 6'h1f == _T_718 ? welem[31] : _GEN_8160; // @[Execute.scala 117:10]
  assign _GEN_8162 = 6'h20 == _T_718 ? welem[32] : _GEN_8161; // @[Execute.scala 117:10]
  assign _GEN_8163 = 6'h21 == _T_718 ? welem[33] : _GEN_8162; // @[Execute.scala 117:10]
  assign _GEN_8164 = 6'h22 == _T_718 ? welem[34] : _GEN_8163; // @[Execute.scala 117:10]
  assign _GEN_8165 = 6'h23 == _T_718 ? welem[35] : _GEN_8164; // @[Execute.scala 117:10]
  assign _GEN_8166 = 6'h24 == _T_718 ? welem[36] : _GEN_8165; // @[Execute.scala 117:10]
  assign _GEN_8167 = 6'h25 == _T_718 ? welem[37] : _GEN_8166; // @[Execute.scala 117:10]
  assign _GEN_8168 = 6'h26 == _T_718 ? welem[38] : _GEN_8167; // @[Execute.scala 117:10]
  assign _GEN_8169 = 6'h27 == _T_718 ? welem[39] : _GEN_8168; // @[Execute.scala 117:10]
  assign _GEN_8170 = 6'h28 == _T_718 ? welem[40] : _GEN_8169; // @[Execute.scala 117:10]
  assign _GEN_8171 = 6'h29 == _T_718 ? welem[41] : _GEN_8170; // @[Execute.scala 117:10]
  assign _GEN_8172 = 6'h2a == _T_718 ? welem[42] : _GEN_8171; // @[Execute.scala 117:10]
  assign _GEN_8173 = 6'h2b == _T_718 ? welem[43] : _GEN_8172; // @[Execute.scala 117:10]
  assign _GEN_8174 = 6'h2c == _T_718 ? welem[44] : _GEN_8173; // @[Execute.scala 117:10]
  assign _GEN_8175 = 6'h2d == _T_718 ? welem[45] : _GEN_8174; // @[Execute.scala 117:10]
  assign _GEN_8176 = 6'h2e == _T_718 ? welem[46] : _GEN_8175; // @[Execute.scala 117:10]
  assign _GEN_8177 = 6'h2f == _T_718 ? welem[47] : _GEN_8176; // @[Execute.scala 117:10]
  assign _GEN_8178 = 6'h30 == _T_718 ? welem[48] : _GEN_8177; // @[Execute.scala 117:10]
  assign _GEN_8179 = 6'h31 == _T_718 ? welem[49] : _GEN_8178; // @[Execute.scala 117:10]
  assign _GEN_8180 = 6'h32 == _T_718 ? welem[50] : _GEN_8179; // @[Execute.scala 117:10]
  assign _GEN_8181 = 6'h33 == _T_718 ? welem[51] : _GEN_8180; // @[Execute.scala 117:10]
  assign _GEN_8182 = 6'h34 == _T_718 ? welem[52] : _GEN_8181; // @[Execute.scala 117:10]
  assign _GEN_8183 = 6'h35 == _T_718 ? welem[53] : _GEN_8182; // @[Execute.scala 117:10]
  assign _GEN_8184 = 6'h36 == _T_718 ? welem[54] : _GEN_8183; // @[Execute.scala 117:10]
  assign _GEN_8185 = 6'h37 == _T_718 ? welem[55] : _GEN_8184; // @[Execute.scala 117:10]
  assign _GEN_8186 = 6'h38 == _T_718 ? welem[56] : _GEN_8185; // @[Execute.scala 117:10]
  assign _GEN_8187 = 6'h39 == _T_718 ? welem[57] : _GEN_8186; // @[Execute.scala 117:10]
  assign _GEN_8188 = 6'h3a == _T_718 ? welem[58] : _GEN_8187; // @[Execute.scala 117:10]
  assign _GEN_8189 = 6'h3b == _T_718 ? welem[59] : _GEN_8188; // @[Execute.scala 117:10]
  assign _GEN_8190 = 6'h3c == _T_718 ? welem[60] : _GEN_8189; // @[Execute.scala 117:10]
  assign _GEN_8191 = 6'h3d == _T_718 ? welem[61] : _GEN_8190; // @[Execute.scala 117:10]
  assign _GEN_8192 = 6'h3e == _T_718 ? welem[62] : _GEN_8191; // @[Execute.scala 117:10]
  assign _GEN_8193 = 6'h3f == _T_718 ? welem[63] : _GEN_8192; // @[Execute.scala 117:10]
  assign _T_721 = _T_712 ? _GEN_8129 : _GEN_8193; // @[Execute.scala 117:10]
  assign _T_722 = r < 6'h1; // @[Execute.scala 117:15]
  assign _T_724 = r - 6'h1; // @[Execute.scala 117:37]
  assign _T_728 = 6'h3f + r; // @[Execute.scala 117:60]
  assign _GEN_8195 = 6'h1 == _T_724 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8196 = 6'h2 == _T_724 ? welem[2] : _GEN_8195; // @[Execute.scala 117:10]
  assign _GEN_8197 = 6'h3 == _T_724 ? welem[3] : _GEN_8196; // @[Execute.scala 117:10]
  assign _GEN_8198 = 6'h4 == _T_724 ? welem[4] : _GEN_8197; // @[Execute.scala 117:10]
  assign _GEN_8199 = 6'h5 == _T_724 ? welem[5] : _GEN_8198; // @[Execute.scala 117:10]
  assign _GEN_8200 = 6'h6 == _T_724 ? welem[6] : _GEN_8199; // @[Execute.scala 117:10]
  assign _GEN_8201 = 6'h7 == _T_724 ? welem[7] : _GEN_8200; // @[Execute.scala 117:10]
  assign _GEN_8202 = 6'h8 == _T_724 ? welem[8] : _GEN_8201; // @[Execute.scala 117:10]
  assign _GEN_8203 = 6'h9 == _T_724 ? welem[9] : _GEN_8202; // @[Execute.scala 117:10]
  assign _GEN_8204 = 6'ha == _T_724 ? welem[10] : _GEN_8203; // @[Execute.scala 117:10]
  assign _GEN_8205 = 6'hb == _T_724 ? welem[11] : _GEN_8204; // @[Execute.scala 117:10]
  assign _GEN_8206 = 6'hc == _T_724 ? welem[12] : _GEN_8205; // @[Execute.scala 117:10]
  assign _GEN_8207 = 6'hd == _T_724 ? welem[13] : _GEN_8206; // @[Execute.scala 117:10]
  assign _GEN_8208 = 6'he == _T_724 ? welem[14] : _GEN_8207; // @[Execute.scala 117:10]
  assign _GEN_8209 = 6'hf == _T_724 ? welem[15] : _GEN_8208; // @[Execute.scala 117:10]
  assign _GEN_8210 = 6'h10 == _T_724 ? welem[16] : _GEN_8209; // @[Execute.scala 117:10]
  assign _GEN_8211 = 6'h11 == _T_724 ? welem[17] : _GEN_8210; // @[Execute.scala 117:10]
  assign _GEN_8212 = 6'h12 == _T_724 ? welem[18] : _GEN_8211; // @[Execute.scala 117:10]
  assign _GEN_8213 = 6'h13 == _T_724 ? welem[19] : _GEN_8212; // @[Execute.scala 117:10]
  assign _GEN_8214 = 6'h14 == _T_724 ? welem[20] : _GEN_8213; // @[Execute.scala 117:10]
  assign _GEN_8215 = 6'h15 == _T_724 ? welem[21] : _GEN_8214; // @[Execute.scala 117:10]
  assign _GEN_8216 = 6'h16 == _T_724 ? welem[22] : _GEN_8215; // @[Execute.scala 117:10]
  assign _GEN_8217 = 6'h17 == _T_724 ? welem[23] : _GEN_8216; // @[Execute.scala 117:10]
  assign _GEN_8218 = 6'h18 == _T_724 ? welem[24] : _GEN_8217; // @[Execute.scala 117:10]
  assign _GEN_8219 = 6'h19 == _T_724 ? welem[25] : _GEN_8218; // @[Execute.scala 117:10]
  assign _GEN_8220 = 6'h1a == _T_724 ? welem[26] : _GEN_8219; // @[Execute.scala 117:10]
  assign _GEN_8221 = 6'h1b == _T_724 ? welem[27] : _GEN_8220; // @[Execute.scala 117:10]
  assign _GEN_8222 = 6'h1c == _T_724 ? welem[28] : _GEN_8221; // @[Execute.scala 117:10]
  assign _GEN_8223 = 6'h1d == _T_724 ? welem[29] : _GEN_8222; // @[Execute.scala 117:10]
  assign _GEN_8224 = 6'h1e == _T_724 ? welem[30] : _GEN_8223; // @[Execute.scala 117:10]
  assign _GEN_8225 = 6'h1f == _T_724 ? welem[31] : _GEN_8224; // @[Execute.scala 117:10]
  assign _GEN_8226 = 6'h20 == _T_724 ? welem[32] : _GEN_8225; // @[Execute.scala 117:10]
  assign _GEN_8227 = 6'h21 == _T_724 ? welem[33] : _GEN_8226; // @[Execute.scala 117:10]
  assign _GEN_8228 = 6'h22 == _T_724 ? welem[34] : _GEN_8227; // @[Execute.scala 117:10]
  assign _GEN_8229 = 6'h23 == _T_724 ? welem[35] : _GEN_8228; // @[Execute.scala 117:10]
  assign _GEN_8230 = 6'h24 == _T_724 ? welem[36] : _GEN_8229; // @[Execute.scala 117:10]
  assign _GEN_8231 = 6'h25 == _T_724 ? welem[37] : _GEN_8230; // @[Execute.scala 117:10]
  assign _GEN_8232 = 6'h26 == _T_724 ? welem[38] : _GEN_8231; // @[Execute.scala 117:10]
  assign _GEN_8233 = 6'h27 == _T_724 ? welem[39] : _GEN_8232; // @[Execute.scala 117:10]
  assign _GEN_8234 = 6'h28 == _T_724 ? welem[40] : _GEN_8233; // @[Execute.scala 117:10]
  assign _GEN_8235 = 6'h29 == _T_724 ? welem[41] : _GEN_8234; // @[Execute.scala 117:10]
  assign _GEN_8236 = 6'h2a == _T_724 ? welem[42] : _GEN_8235; // @[Execute.scala 117:10]
  assign _GEN_8237 = 6'h2b == _T_724 ? welem[43] : _GEN_8236; // @[Execute.scala 117:10]
  assign _GEN_8238 = 6'h2c == _T_724 ? welem[44] : _GEN_8237; // @[Execute.scala 117:10]
  assign _GEN_8239 = 6'h2d == _T_724 ? welem[45] : _GEN_8238; // @[Execute.scala 117:10]
  assign _GEN_8240 = 6'h2e == _T_724 ? welem[46] : _GEN_8239; // @[Execute.scala 117:10]
  assign _GEN_8241 = 6'h2f == _T_724 ? welem[47] : _GEN_8240; // @[Execute.scala 117:10]
  assign _GEN_8242 = 6'h30 == _T_724 ? welem[48] : _GEN_8241; // @[Execute.scala 117:10]
  assign _GEN_8243 = 6'h31 == _T_724 ? welem[49] : _GEN_8242; // @[Execute.scala 117:10]
  assign _GEN_8244 = 6'h32 == _T_724 ? welem[50] : _GEN_8243; // @[Execute.scala 117:10]
  assign _GEN_8245 = 6'h33 == _T_724 ? welem[51] : _GEN_8244; // @[Execute.scala 117:10]
  assign _GEN_8246 = 6'h34 == _T_724 ? welem[52] : _GEN_8245; // @[Execute.scala 117:10]
  assign _GEN_8247 = 6'h35 == _T_724 ? welem[53] : _GEN_8246; // @[Execute.scala 117:10]
  assign _GEN_8248 = 6'h36 == _T_724 ? welem[54] : _GEN_8247; // @[Execute.scala 117:10]
  assign _GEN_8249 = 6'h37 == _T_724 ? welem[55] : _GEN_8248; // @[Execute.scala 117:10]
  assign _GEN_8250 = 6'h38 == _T_724 ? welem[56] : _GEN_8249; // @[Execute.scala 117:10]
  assign _GEN_8251 = 6'h39 == _T_724 ? welem[57] : _GEN_8250; // @[Execute.scala 117:10]
  assign _GEN_8252 = 6'h3a == _T_724 ? welem[58] : _GEN_8251; // @[Execute.scala 117:10]
  assign _GEN_8253 = 6'h3b == _T_724 ? welem[59] : _GEN_8252; // @[Execute.scala 117:10]
  assign _GEN_8254 = 6'h3c == _T_724 ? welem[60] : _GEN_8253; // @[Execute.scala 117:10]
  assign _GEN_8255 = 6'h3d == _T_724 ? welem[61] : _GEN_8254; // @[Execute.scala 117:10]
  assign _GEN_8256 = 6'h3e == _T_724 ? welem[62] : _GEN_8255; // @[Execute.scala 117:10]
  assign _GEN_8257 = 6'h3f == _T_724 ? welem[63] : _GEN_8256; // @[Execute.scala 117:10]
  assign _GEN_8259 = 6'h1 == _T_728 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8260 = 6'h2 == _T_728 ? welem[2] : _GEN_8259; // @[Execute.scala 117:10]
  assign _GEN_8261 = 6'h3 == _T_728 ? welem[3] : _GEN_8260; // @[Execute.scala 117:10]
  assign _GEN_8262 = 6'h4 == _T_728 ? welem[4] : _GEN_8261; // @[Execute.scala 117:10]
  assign _GEN_8263 = 6'h5 == _T_728 ? welem[5] : _GEN_8262; // @[Execute.scala 117:10]
  assign _GEN_8264 = 6'h6 == _T_728 ? welem[6] : _GEN_8263; // @[Execute.scala 117:10]
  assign _GEN_8265 = 6'h7 == _T_728 ? welem[7] : _GEN_8264; // @[Execute.scala 117:10]
  assign _GEN_8266 = 6'h8 == _T_728 ? welem[8] : _GEN_8265; // @[Execute.scala 117:10]
  assign _GEN_8267 = 6'h9 == _T_728 ? welem[9] : _GEN_8266; // @[Execute.scala 117:10]
  assign _GEN_8268 = 6'ha == _T_728 ? welem[10] : _GEN_8267; // @[Execute.scala 117:10]
  assign _GEN_8269 = 6'hb == _T_728 ? welem[11] : _GEN_8268; // @[Execute.scala 117:10]
  assign _GEN_8270 = 6'hc == _T_728 ? welem[12] : _GEN_8269; // @[Execute.scala 117:10]
  assign _GEN_8271 = 6'hd == _T_728 ? welem[13] : _GEN_8270; // @[Execute.scala 117:10]
  assign _GEN_8272 = 6'he == _T_728 ? welem[14] : _GEN_8271; // @[Execute.scala 117:10]
  assign _GEN_8273 = 6'hf == _T_728 ? welem[15] : _GEN_8272; // @[Execute.scala 117:10]
  assign _GEN_8274 = 6'h10 == _T_728 ? welem[16] : _GEN_8273; // @[Execute.scala 117:10]
  assign _GEN_8275 = 6'h11 == _T_728 ? welem[17] : _GEN_8274; // @[Execute.scala 117:10]
  assign _GEN_8276 = 6'h12 == _T_728 ? welem[18] : _GEN_8275; // @[Execute.scala 117:10]
  assign _GEN_8277 = 6'h13 == _T_728 ? welem[19] : _GEN_8276; // @[Execute.scala 117:10]
  assign _GEN_8278 = 6'h14 == _T_728 ? welem[20] : _GEN_8277; // @[Execute.scala 117:10]
  assign _GEN_8279 = 6'h15 == _T_728 ? welem[21] : _GEN_8278; // @[Execute.scala 117:10]
  assign _GEN_8280 = 6'h16 == _T_728 ? welem[22] : _GEN_8279; // @[Execute.scala 117:10]
  assign _GEN_8281 = 6'h17 == _T_728 ? welem[23] : _GEN_8280; // @[Execute.scala 117:10]
  assign _GEN_8282 = 6'h18 == _T_728 ? welem[24] : _GEN_8281; // @[Execute.scala 117:10]
  assign _GEN_8283 = 6'h19 == _T_728 ? welem[25] : _GEN_8282; // @[Execute.scala 117:10]
  assign _GEN_8284 = 6'h1a == _T_728 ? welem[26] : _GEN_8283; // @[Execute.scala 117:10]
  assign _GEN_8285 = 6'h1b == _T_728 ? welem[27] : _GEN_8284; // @[Execute.scala 117:10]
  assign _GEN_8286 = 6'h1c == _T_728 ? welem[28] : _GEN_8285; // @[Execute.scala 117:10]
  assign _GEN_8287 = 6'h1d == _T_728 ? welem[29] : _GEN_8286; // @[Execute.scala 117:10]
  assign _GEN_8288 = 6'h1e == _T_728 ? welem[30] : _GEN_8287; // @[Execute.scala 117:10]
  assign _GEN_8289 = 6'h1f == _T_728 ? welem[31] : _GEN_8288; // @[Execute.scala 117:10]
  assign _GEN_8290 = 6'h20 == _T_728 ? welem[32] : _GEN_8289; // @[Execute.scala 117:10]
  assign _GEN_8291 = 6'h21 == _T_728 ? welem[33] : _GEN_8290; // @[Execute.scala 117:10]
  assign _GEN_8292 = 6'h22 == _T_728 ? welem[34] : _GEN_8291; // @[Execute.scala 117:10]
  assign _GEN_8293 = 6'h23 == _T_728 ? welem[35] : _GEN_8292; // @[Execute.scala 117:10]
  assign _GEN_8294 = 6'h24 == _T_728 ? welem[36] : _GEN_8293; // @[Execute.scala 117:10]
  assign _GEN_8295 = 6'h25 == _T_728 ? welem[37] : _GEN_8294; // @[Execute.scala 117:10]
  assign _GEN_8296 = 6'h26 == _T_728 ? welem[38] : _GEN_8295; // @[Execute.scala 117:10]
  assign _GEN_8297 = 6'h27 == _T_728 ? welem[39] : _GEN_8296; // @[Execute.scala 117:10]
  assign _GEN_8298 = 6'h28 == _T_728 ? welem[40] : _GEN_8297; // @[Execute.scala 117:10]
  assign _GEN_8299 = 6'h29 == _T_728 ? welem[41] : _GEN_8298; // @[Execute.scala 117:10]
  assign _GEN_8300 = 6'h2a == _T_728 ? welem[42] : _GEN_8299; // @[Execute.scala 117:10]
  assign _GEN_8301 = 6'h2b == _T_728 ? welem[43] : _GEN_8300; // @[Execute.scala 117:10]
  assign _GEN_8302 = 6'h2c == _T_728 ? welem[44] : _GEN_8301; // @[Execute.scala 117:10]
  assign _GEN_8303 = 6'h2d == _T_728 ? welem[45] : _GEN_8302; // @[Execute.scala 117:10]
  assign _GEN_8304 = 6'h2e == _T_728 ? welem[46] : _GEN_8303; // @[Execute.scala 117:10]
  assign _GEN_8305 = 6'h2f == _T_728 ? welem[47] : _GEN_8304; // @[Execute.scala 117:10]
  assign _GEN_8306 = 6'h30 == _T_728 ? welem[48] : _GEN_8305; // @[Execute.scala 117:10]
  assign _GEN_8307 = 6'h31 == _T_728 ? welem[49] : _GEN_8306; // @[Execute.scala 117:10]
  assign _GEN_8308 = 6'h32 == _T_728 ? welem[50] : _GEN_8307; // @[Execute.scala 117:10]
  assign _GEN_8309 = 6'h33 == _T_728 ? welem[51] : _GEN_8308; // @[Execute.scala 117:10]
  assign _GEN_8310 = 6'h34 == _T_728 ? welem[52] : _GEN_8309; // @[Execute.scala 117:10]
  assign _GEN_8311 = 6'h35 == _T_728 ? welem[53] : _GEN_8310; // @[Execute.scala 117:10]
  assign _GEN_8312 = 6'h36 == _T_728 ? welem[54] : _GEN_8311; // @[Execute.scala 117:10]
  assign _GEN_8313 = 6'h37 == _T_728 ? welem[55] : _GEN_8312; // @[Execute.scala 117:10]
  assign _GEN_8314 = 6'h38 == _T_728 ? welem[56] : _GEN_8313; // @[Execute.scala 117:10]
  assign _GEN_8315 = 6'h39 == _T_728 ? welem[57] : _GEN_8314; // @[Execute.scala 117:10]
  assign _GEN_8316 = 6'h3a == _T_728 ? welem[58] : _GEN_8315; // @[Execute.scala 117:10]
  assign _GEN_8317 = 6'h3b == _T_728 ? welem[59] : _GEN_8316; // @[Execute.scala 117:10]
  assign _GEN_8318 = 6'h3c == _T_728 ? welem[60] : _GEN_8317; // @[Execute.scala 117:10]
  assign _GEN_8319 = 6'h3d == _T_728 ? welem[61] : _GEN_8318; // @[Execute.scala 117:10]
  assign _GEN_8320 = 6'h3e == _T_728 ? welem[62] : _GEN_8319; // @[Execute.scala 117:10]
  assign _GEN_8321 = 6'h3f == _T_728 ? welem[63] : _GEN_8320; // @[Execute.scala 117:10]
  assign _T_731 = _T_722 ? _GEN_8257 : _GEN_8321; // @[Execute.scala 117:10]
  assign _T_739 = {_T_171,_T_161,_T_151,_T_141,_T_131,_T_121,_T_111,_GEN_193}; // @[Execute.scala 302:55]
  assign _T_747 = {_T_251,_T_241,_T_231,_T_221,_T_211,_T_201,_T_191,_T_181,_T_739}; // @[Execute.scala 302:55]
  assign _T_754 = {_T_331,_T_321,_T_311,_T_301,_T_291,_T_281,_T_271,_T_261}; // @[Execute.scala 302:55]
  assign _T_763 = {_T_411,_T_401,_T_391,_T_381,_T_371,_T_361,_T_351,_T_341,_T_754,_T_747}; // @[Execute.scala 302:55]
  assign _T_770 = {_T_491,_T_481,_T_471,_T_461,_T_451,_T_441,_T_431,_T_421}; // @[Execute.scala 302:55]
  assign _T_778 = {_T_571,_T_561,_T_551,_T_541,_T_531,_T_521,_T_511,_T_501,_T_770}; // @[Execute.scala 302:55]
  assign _T_785 = {_T_651,_T_641,_T_631,_T_621,_T_611,_T_601,_T_591,_T_581}; // @[Execute.scala 302:55]
  assign _T_794 = {_T_731,_T_721,_T_711,_T_701,_T_691,_T_681,_T_671,_T_661,_T_785,_T_778}; // @[Execute.scala 302:55]
  assign _T_795 = {_T_794,_T_763}; // @[Execute.scala 302:55]
  assign _GEN_8323 = 7'h1 == onesD[6:0] ? 64'h1 : 64'h0; // @[Execute.scala 304:9]
  assign _GEN_8324 = 7'h2 == onesD[6:0] ? 64'h3 : _GEN_8323; // @[Execute.scala 304:9]
  assign _GEN_8325 = 7'h3 == onesD[6:0] ? 64'h7 : _GEN_8324; // @[Execute.scala 304:9]
  assign _GEN_8326 = 7'h4 == onesD[6:0] ? 64'hf : _GEN_8325; // @[Execute.scala 304:9]
  assign _GEN_8327 = 7'h5 == onesD[6:0] ? 64'h1f : _GEN_8326; // @[Execute.scala 304:9]
  assign _GEN_8328 = 7'h6 == onesD[6:0] ? 64'h3f : _GEN_8327; // @[Execute.scala 304:9]
  assign _GEN_8329 = 7'h7 == onesD[6:0] ? 64'h7f : _GEN_8328; // @[Execute.scala 304:9]
  assign _GEN_8330 = 7'h8 == onesD[6:0] ? 64'hff : _GEN_8329; // @[Execute.scala 304:9]
  assign _GEN_8331 = 7'h9 == onesD[6:0] ? 64'h1ff : _GEN_8330; // @[Execute.scala 304:9]
  assign _GEN_8332 = 7'ha == onesD[6:0] ? 64'h3ff : _GEN_8331; // @[Execute.scala 304:9]
  assign _GEN_8333 = 7'hb == onesD[6:0] ? 64'h7ff : _GEN_8332; // @[Execute.scala 304:9]
  assign _GEN_8334 = 7'hc == onesD[6:0] ? 64'hfff : _GEN_8333; // @[Execute.scala 304:9]
  assign _GEN_8335 = 7'hd == onesD[6:0] ? 64'h1fff : _GEN_8334; // @[Execute.scala 304:9]
  assign _GEN_8336 = 7'he == onesD[6:0] ? 64'h3fff : _GEN_8335; // @[Execute.scala 304:9]
  assign _GEN_8337 = 7'hf == onesD[6:0] ? 64'h7fff : _GEN_8336; // @[Execute.scala 304:9]
  assign _GEN_8338 = 7'h10 == onesD[6:0] ? 64'hffff : _GEN_8337; // @[Execute.scala 304:9]
  assign _GEN_8339 = 7'h11 == onesD[6:0] ? 64'h1ffff : _GEN_8338; // @[Execute.scala 304:9]
  assign _GEN_8340 = 7'h12 == onesD[6:0] ? 64'h3ffff : _GEN_8339; // @[Execute.scala 304:9]
  assign _GEN_8341 = 7'h13 == onesD[6:0] ? 64'h7ffff : _GEN_8340; // @[Execute.scala 304:9]
  assign _GEN_8342 = 7'h14 == onesD[6:0] ? 64'hfffff : _GEN_8341; // @[Execute.scala 304:9]
  assign _GEN_8343 = 7'h15 == onesD[6:0] ? 64'h1fffff : _GEN_8342; // @[Execute.scala 304:9]
  assign _GEN_8344 = 7'h16 == onesD[6:0] ? 64'h3fffff : _GEN_8343; // @[Execute.scala 304:9]
  assign _GEN_8345 = 7'h17 == onesD[6:0] ? 64'h7fffff : _GEN_8344; // @[Execute.scala 304:9]
  assign _GEN_8346 = 7'h18 == onesD[6:0] ? 64'hffffff : _GEN_8345; // @[Execute.scala 304:9]
  assign _GEN_8347 = 7'h19 == onesD[6:0] ? 64'h1ffffff : _GEN_8346; // @[Execute.scala 304:9]
  assign _GEN_8348 = 7'h1a == onesD[6:0] ? 64'h3ffffff : _GEN_8347; // @[Execute.scala 304:9]
  assign _GEN_8349 = 7'h1b == onesD[6:0] ? 64'h7ffffff : _GEN_8348; // @[Execute.scala 304:9]
  assign _GEN_8350 = 7'h1c == onesD[6:0] ? 64'hfffffff : _GEN_8349; // @[Execute.scala 304:9]
  assign _GEN_8351 = 7'h1d == onesD[6:0] ? 64'h1fffffff : _GEN_8350; // @[Execute.scala 304:9]
  assign _GEN_8352 = 7'h1e == onesD[6:0] ? 64'h3fffffff : _GEN_8351; // @[Execute.scala 304:9]
  assign _GEN_8353 = 7'h1f == onesD[6:0] ? 64'h7fffffff : _GEN_8352; // @[Execute.scala 304:9]
  assign _GEN_8354 = 7'h20 == onesD[6:0] ? 64'hffffffff : _GEN_8353; // @[Execute.scala 304:9]
  assign _GEN_8355 = 7'h21 == onesD[6:0] ? 64'h1ffffffff : _GEN_8354; // @[Execute.scala 304:9]
  assign _GEN_8356 = 7'h22 == onesD[6:0] ? 64'h3ffffffff : _GEN_8355; // @[Execute.scala 304:9]
  assign _GEN_8357 = 7'h23 == onesD[6:0] ? 64'h7ffffffff : _GEN_8356; // @[Execute.scala 304:9]
  assign _GEN_8358 = 7'h24 == onesD[6:0] ? 64'hfffffffff : _GEN_8357; // @[Execute.scala 304:9]
  assign _GEN_8359 = 7'h25 == onesD[6:0] ? 64'h1fffffffff : _GEN_8358; // @[Execute.scala 304:9]
  assign _GEN_8360 = 7'h26 == onesD[6:0] ? 64'h3fffffffff : _GEN_8359; // @[Execute.scala 304:9]
  assign _GEN_8361 = 7'h27 == onesD[6:0] ? 64'h7fffffffff : _GEN_8360; // @[Execute.scala 304:9]
  assign _GEN_8362 = 7'h28 == onesD[6:0] ? 64'hffffffffff : _GEN_8361; // @[Execute.scala 304:9]
  assign _GEN_8363 = 7'h29 == onesD[6:0] ? 64'h1ffffffffff : _GEN_8362; // @[Execute.scala 304:9]
  assign _GEN_8364 = 7'h2a == onesD[6:0] ? 64'h3ffffffffff : _GEN_8363; // @[Execute.scala 304:9]
  assign _GEN_8365 = 7'h2b == onesD[6:0] ? 64'h7ffffffffff : _GEN_8364; // @[Execute.scala 304:9]
  assign _GEN_8366 = 7'h2c == onesD[6:0] ? 64'hfffffffffff : _GEN_8365; // @[Execute.scala 304:9]
  assign _GEN_8367 = 7'h2d == onesD[6:0] ? 64'h1fffffffffff : _GEN_8366; // @[Execute.scala 304:9]
  assign _GEN_8368 = 7'h2e == onesD[6:0] ? 64'h3fffffffffff : _GEN_8367; // @[Execute.scala 304:9]
  assign _GEN_8369 = 7'h2f == onesD[6:0] ? 64'h7fffffffffff : _GEN_8368; // @[Execute.scala 304:9]
  assign _GEN_8370 = 7'h30 == onesD[6:0] ? 64'hffffffffffff : _GEN_8369; // @[Execute.scala 304:9]
  assign _GEN_8371 = 7'h31 == onesD[6:0] ? 64'h1ffffffffffff : _GEN_8370; // @[Execute.scala 304:9]
  assign _GEN_8372 = 7'h32 == onesD[6:0] ? 64'h3ffffffffffff : _GEN_8371; // @[Execute.scala 304:9]
  assign _GEN_8373 = 7'h33 == onesD[6:0] ? 64'h7ffffffffffff : _GEN_8372; // @[Execute.scala 304:9]
  assign _GEN_8374 = 7'h34 == onesD[6:0] ? 64'hfffffffffffff : _GEN_8373; // @[Execute.scala 304:9]
  assign _GEN_8375 = 7'h35 == onesD[6:0] ? 64'h1fffffffffffff : _GEN_8374; // @[Execute.scala 304:9]
  assign _GEN_8376 = 7'h36 == onesD[6:0] ? 64'h3fffffffffffff : _GEN_8375; // @[Execute.scala 304:9]
  assign _GEN_8377 = 7'h37 == onesD[6:0] ? 64'h7fffffffffffff : _GEN_8376; // @[Execute.scala 304:9]
  assign _GEN_8378 = 7'h38 == onesD[6:0] ? 64'hffffffffffffff : _GEN_8377; // @[Execute.scala 304:9]
  assign _GEN_8379 = 7'h39 == onesD[6:0] ? 64'h1ffffffffffffff : _GEN_8378; // @[Execute.scala 304:9]
  assign _GEN_8380 = 7'h3a == onesD[6:0] ? 64'h3ffffffffffffff : _GEN_8379; // @[Execute.scala 304:9]
  assign _GEN_8381 = 7'h3b == onesD[6:0] ? 64'h7ffffffffffffff : _GEN_8380; // @[Execute.scala 304:9]
  assign _GEN_8382 = 7'h3c == onesD[6:0] ? 64'hfffffffffffffff : _GEN_8381; // @[Execute.scala 304:9]
  assign _GEN_8383 = 7'h3d == onesD[6:0] ? 64'h1fffffffffffffff : _GEN_8382; // @[Execute.scala 304:9]
  assign _GEN_8384 = 7'h3e == onesD[6:0] ? 64'h3fffffffffffffff : _GEN_8383; // @[Execute.scala 304:9]
  assign _GEN_8385 = 7'h3f == onesD[6:0] ? 64'h7fffffffffffffff : _GEN_8384; // @[Execute.scala 304:9]
  assign _GEN_10438 = {{1'd0}, r[4:0]}; // @[Execute.scala 117:37]
  assign _T_835 = _GEN_10438 - 6'h20; // @[Execute.scala 117:37]
  assign _GEN_8388 = 5'h1 == _T_835[4:0] ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8389 = 5'h2 == _T_835[4:0] ? welem[2] : _GEN_8388; // @[Execute.scala 117:10]
  assign _GEN_8390 = 5'h3 == _T_835[4:0] ? welem[3] : _GEN_8389; // @[Execute.scala 117:10]
  assign _GEN_8391 = 5'h4 == _T_835[4:0] ? welem[4] : _GEN_8390; // @[Execute.scala 117:10]
  assign _GEN_8392 = 5'h5 == _T_835[4:0] ? welem[5] : _GEN_8391; // @[Execute.scala 117:10]
  assign _GEN_8393 = 5'h6 == _T_835[4:0] ? welem[6] : _GEN_8392; // @[Execute.scala 117:10]
  assign _GEN_8394 = 5'h7 == _T_835[4:0] ? welem[7] : _GEN_8393; // @[Execute.scala 117:10]
  assign _GEN_8395 = 5'h8 == _T_835[4:0] ? welem[8] : _GEN_8394; // @[Execute.scala 117:10]
  assign _GEN_8396 = 5'h9 == _T_835[4:0] ? welem[9] : _GEN_8395; // @[Execute.scala 117:10]
  assign _GEN_8397 = 5'ha == _T_835[4:0] ? welem[10] : _GEN_8396; // @[Execute.scala 117:10]
  assign _GEN_8398 = 5'hb == _T_835[4:0] ? welem[11] : _GEN_8397; // @[Execute.scala 117:10]
  assign _GEN_8399 = 5'hc == _T_835[4:0] ? welem[12] : _GEN_8398; // @[Execute.scala 117:10]
  assign _GEN_8400 = 5'hd == _T_835[4:0] ? welem[13] : _GEN_8399; // @[Execute.scala 117:10]
  assign _GEN_8401 = 5'he == _T_835[4:0] ? welem[14] : _GEN_8400; // @[Execute.scala 117:10]
  assign _GEN_8402 = 5'hf == _T_835[4:0] ? welem[15] : _GEN_8401; // @[Execute.scala 117:10]
  assign _GEN_8403 = 5'h10 == _T_835[4:0] ? welem[16] : _GEN_8402; // @[Execute.scala 117:10]
  assign _GEN_8404 = 5'h11 == _T_835[4:0] ? welem[17] : _GEN_8403; // @[Execute.scala 117:10]
  assign _GEN_8405 = 5'h12 == _T_835[4:0] ? welem[18] : _GEN_8404; // @[Execute.scala 117:10]
  assign _GEN_8406 = 5'h13 == _T_835[4:0] ? welem[19] : _GEN_8405; // @[Execute.scala 117:10]
  assign _GEN_8407 = 5'h14 == _T_835[4:0] ? welem[20] : _GEN_8406; // @[Execute.scala 117:10]
  assign _GEN_8408 = 5'h15 == _T_835[4:0] ? welem[21] : _GEN_8407; // @[Execute.scala 117:10]
  assign _GEN_8409 = 5'h16 == _T_835[4:0] ? welem[22] : _GEN_8408; // @[Execute.scala 117:10]
  assign _GEN_8410 = 5'h17 == _T_835[4:0] ? welem[23] : _GEN_8409; // @[Execute.scala 117:10]
  assign _GEN_8411 = 5'h18 == _T_835[4:0] ? welem[24] : _GEN_8410; // @[Execute.scala 117:10]
  assign _GEN_8412 = 5'h19 == _T_835[4:0] ? welem[25] : _GEN_8411; // @[Execute.scala 117:10]
  assign _GEN_8413 = 5'h1a == _T_835[4:0] ? welem[26] : _GEN_8412; // @[Execute.scala 117:10]
  assign _GEN_8414 = 5'h1b == _T_835[4:0] ? welem[27] : _GEN_8413; // @[Execute.scala 117:10]
  assign _GEN_8415 = 5'h1c == _T_835[4:0] ? welem[28] : _GEN_8414; // @[Execute.scala 117:10]
  assign _GEN_8416 = 5'h1d == _T_835[4:0] ? welem[29] : _GEN_8415; // @[Execute.scala 117:10]
  assign _GEN_8417 = 5'h1e == _T_835[4:0] ? welem[30] : _GEN_8416; // @[Execute.scala 117:10]
  assign _GEN_8418 = 5'h1f == _T_835[4:0] ? welem[31] : _GEN_8417; // @[Execute.scala 117:10]
  assign _T_840 = r[4:0] < 5'h1f; // @[Execute.scala 117:15]
  assign _T_842 = r[4:0] - 5'h1f; // @[Execute.scala 117:37]
  assign _T_844 = 5'h1 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_8452 = 5'h1 == _T_842 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8453 = 5'h2 == _T_842 ? welem[2] : _GEN_8452; // @[Execute.scala 117:10]
  assign _GEN_8454 = 5'h3 == _T_842 ? welem[3] : _GEN_8453; // @[Execute.scala 117:10]
  assign _GEN_8455 = 5'h4 == _T_842 ? welem[4] : _GEN_8454; // @[Execute.scala 117:10]
  assign _GEN_8456 = 5'h5 == _T_842 ? welem[5] : _GEN_8455; // @[Execute.scala 117:10]
  assign _GEN_8457 = 5'h6 == _T_842 ? welem[6] : _GEN_8456; // @[Execute.scala 117:10]
  assign _GEN_8458 = 5'h7 == _T_842 ? welem[7] : _GEN_8457; // @[Execute.scala 117:10]
  assign _GEN_8459 = 5'h8 == _T_842 ? welem[8] : _GEN_8458; // @[Execute.scala 117:10]
  assign _GEN_8460 = 5'h9 == _T_842 ? welem[9] : _GEN_8459; // @[Execute.scala 117:10]
  assign _GEN_8461 = 5'ha == _T_842 ? welem[10] : _GEN_8460; // @[Execute.scala 117:10]
  assign _GEN_8462 = 5'hb == _T_842 ? welem[11] : _GEN_8461; // @[Execute.scala 117:10]
  assign _GEN_8463 = 5'hc == _T_842 ? welem[12] : _GEN_8462; // @[Execute.scala 117:10]
  assign _GEN_8464 = 5'hd == _T_842 ? welem[13] : _GEN_8463; // @[Execute.scala 117:10]
  assign _GEN_8465 = 5'he == _T_842 ? welem[14] : _GEN_8464; // @[Execute.scala 117:10]
  assign _GEN_8466 = 5'hf == _T_842 ? welem[15] : _GEN_8465; // @[Execute.scala 117:10]
  assign _GEN_8467 = 5'h10 == _T_842 ? welem[16] : _GEN_8466; // @[Execute.scala 117:10]
  assign _GEN_8468 = 5'h11 == _T_842 ? welem[17] : _GEN_8467; // @[Execute.scala 117:10]
  assign _GEN_8469 = 5'h12 == _T_842 ? welem[18] : _GEN_8468; // @[Execute.scala 117:10]
  assign _GEN_8470 = 5'h13 == _T_842 ? welem[19] : _GEN_8469; // @[Execute.scala 117:10]
  assign _GEN_8471 = 5'h14 == _T_842 ? welem[20] : _GEN_8470; // @[Execute.scala 117:10]
  assign _GEN_8472 = 5'h15 == _T_842 ? welem[21] : _GEN_8471; // @[Execute.scala 117:10]
  assign _GEN_8473 = 5'h16 == _T_842 ? welem[22] : _GEN_8472; // @[Execute.scala 117:10]
  assign _GEN_8474 = 5'h17 == _T_842 ? welem[23] : _GEN_8473; // @[Execute.scala 117:10]
  assign _GEN_8475 = 5'h18 == _T_842 ? welem[24] : _GEN_8474; // @[Execute.scala 117:10]
  assign _GEN_8476 = 5'h19 == _T_842 ? welem[25] : _GEN_8475; // @[Execute.scala 117:10]
  assign _GEN_8477 = 5'h1a == _T_842 ? welem[26] : _GEN_8476; // @[Execute.scala 117:10]
  assign _GEN_8478 = 5'h1b == _T_842 ? welem[27] : _GEN_8477; // @[Execute.scala 117:10]
  assign _GEN_8479 = 5'h1c == _T_842 ? welem[28] : _GEN_8478; // @[Execute.scala 117:10]
  assign _GEN_8480 = 5'h1d == _T_842 ? welem[29] : _GEN_8479; // @[Execute.scala 117:10]
  assign _GEN_8481 = 5'h1e == _T_842 ? welem[30] : _GEN_8480; // @[Execute.scala 117:10]
  assign _GEN_8482 = 5'h1f == _T_842 ? welem[31] : _GEN_8481; // @[Execute.scala 117:10]
  assign _GEN_8484 = 5'h1 == _T_844 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8485 = 5'h2 == _T_844 ? welem[2] : _GEN_8484; // @[Execute.scala 117:10]
  assign _GEN_8486 = 5'h3 == _T_844 ? welem[3] : _GEN_8485; // @[Execute.scala 117:10]
  assign _GEN_8487 = 5'h4 == _T_844 ? welem[4] : _GEN_8486; // @[Execute.scala 117:10]
  assign _GEN_8488 = 5'h5 == _T_844 ? welem[5] : _GEN_8487; // @[Execute.scala 117:10]
  assign _GEN_8489 = 5'h6 == _T_844 ? welem[6] : _GEN_8488; // @[Execute.scala 117:10]
  assign _GEN_8490 = 5'h7 == _T_844 ? welem[7] : _GEN_8489; // @[Execute.scala 117:10]
  assign _GEN_8491 = 5'h8 == _T_844 ? welem[8] : _GEN_8490; // @[Execute.scala 117:10]
  assign _GEN_8492 = 5'h9 == _T_844 ? welem[9] : _GEN_8491; // @[Execute.scala 117:10]
  assign _GEN_8493 = 5'ha == _T_844 ? welem[10] : _GEN_8492; // @[Execute.scala 117:10]
  assign _GEN_8494 = 5'hb == _T_844 ? welem[11] : _GEN_8493; // @[Execute.scala 117:10]
  assign _GEN_8495 = 5'hc == _T_844 ? welem[12] : _GEN_8494; // @[Execute.scala 117:10]
  assign _GEN_8496 = 5'hd == _T_844 ? welem[13] : _GEN_8495; // @[Execute.scala 117:10]
  assign _GEN_8497 = 5'he == _T_844 ? welem[14] : _GEN_8496; // @[Execute.scala 117:10]
  assign _GEN_8498 = 5'hf == _T_844 ? welem[15] : _GEN_8497; // @[Execute.scala 117:10]
  assign _GEN_8499 = 5'h10 == _T_844 ? welem[16] : _GEN_8498; // @[Execute.scala 117:10]
  assign _GEN_8500 = 5'h11 == _T_844 ? welem[17] : _GEN_8499; // @[Execute.scala 117:10]
  assign _GEN_8501 = 5'h12 == _T_844 ? welem[18] : _GEN_8500; // @[Execute.scala 117:10]
  assign _GEN_8502 = 5'h13 == _T_844 ? welem[19] : _GEN_8501; // @[Execute.scala 117:10]
  assign _GEN_8503 = 5'h14 == _T_844 ? welem[20] : _GEN_8502; // @[Execute.scala 117:10]
  assign _GEN_8504 = 5'h15 == _T_844 ? welem[21] : _GEN_8503; // @[Execute.scala 117:10]
  assign _GEN_8505 = 5'h16 == _T_844 ? welem[22] : _GEN_8504; // @[Execute.scala 117:10]
  assign _GEN_8506 = 5'h17 == _T_844 ? welem[23] : _GEN_8505; // @[Execute.scala 117:10]
  assign _GEN_8507 = 5'h18 == _T_844 ? welem[24] : _GEN_8506; // @[Execute.scala 117:10]
  assign _GEN_8508 = 5'h19 == _T_844 ? welem[25] : _GEN_8507; // @[Execute.scala 117:10]
  assign _GEN_8509 = 5'h1a == _T_844 ? welem[26] : _GEN_8508; // @[Execute.scala 117:10]
  assign _GEN_8510 = 5'h1b == _T_844 ? welem[27] : _GEN_8509; // @[Execute.scala 117:10]
  assign _GEN_8511 = 5'h1c == _T_844 ? welem[28] : _GEN_8510; // @[Execute.scala 117:10]
  assign _GEN_8512 = 5'h1d == _T_844 ? welem[29] : _GEN_8511; // @[Execute.scala 117:10]
  assign _GEN_8513 = 5'h1e == _T_844 ? welem[30] : _GEN_8512; // @[Execute.scala 117:10]
  assign _GEN_8514 = 5'h1f == _T_844 ? welem[31] : _GEN_8513; // @[Execute.scala 117:10]
  assign _T_845 = _T_840 ? _GEN_8482 : _GEN_8514; // @[Execute.scala 117:10]
  assign _T_846 = r[4:0] < 5'h1e; // @[Execute.scala 117:15]
  assign _T_848 = r[4:0] - 5'h1e; // @[Execute.scala 117:37]
  assign _T_850 = 5'h2 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_8516 = 5'h1 == _T_848 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8517 = 5'h2 == _T_848 ? welem[2] : _GEN_8516; // @[Execute.scala 117:10]
  assign _GEN_8518 = 5'h3 == _T_848 ? welem[3] : _GEN_8517; // @[Execute.scala 117:10]
  assign _GEN_8519 = 5'h4 == _T_848 ? welem[4] : _GEN_8518; // @[Execute.scala 117:10]
  assign _GEN_8520 = 5'h5 == _T_848 ? welem[5] : _GEN_8519; // @[Execute.scala 117:10]
  assign _GEN_8521 = 5'h6 == _T_848 ? welem[6] : _GEN_8520; // @[Execute.scala 117:10]
  assign _GEN_8522 = 5'h7 == _T_848 ? welem[7] : _GEN_8521; // @[Execute.scala 117:10]
  assign _GEN_8523 = 5'h8 == _T_848 ? welem[8] : _GEN_8522; // @[Execute.scala 117:10]
  assign _GEN_8524 = 5'h9 == _T_848 ? welem[9] : _GEN_8523; // @[Execute.scala 117:10]
  assign _GEN_8525 = 5'ha == _T_848 ? welem[10] : _GEN_8524; // @[Execute.scala 117:10]
  assign _GEN_8526 = 5'hb == _T_848 ? welem[11] : _GEN_8525; // @[Execute.scala 117:10]
  assign _GEN_8527 = 5'hc == _T_848 ? welem[12] : _GEN_8526; // @[Execute.scala 117:10]
  assign _GEN_8528 = 5'hd == _T_848 ? welem[13] : _GEN_8527; // @[Execute.scala 117:10]
  assign _GEN_8529 = 5'he == _T_848 ? welem[14] : _GEN_8528; // @[Execute.scala 117:10]
  assign _GEN_8530 = 5'hf == _T_848 ? welem[15] : _GEN_8529; // @[Execute.scala 117:10]
  assign _GEN_8531 = 5'h10 == _T_848 ? welem[16] : _GEN_8530; // @[Execute.scala 117:10]
  assign _GEN_8532 = 5'h11 == _T_848 ? welem[17] : _GEN_8531; // @[Execute.scala 117:10]
  assign _GEN_8533 = 5'h12 == _T_848 ? welem[18] : _GEN_8532; // @[Execute.scala 117:10]
  assign _GEN_8534 = 5'h13 == _T_848 ? welem[19] : _GEN_8533; // @[Execute.scala 117:10]
  assign _GEN_8535 = 5'h14 == _T_848 ? welem[20] : _GEN_8534; // @[Execute.scala 117:10]
  assign _GEN_8536 = 5'h15 == _T_848 ? welem[21] : _GEN_8535; // @[Execute.scala 117:10]
  assign _GEN_8537 = 5'h16 == _T_848 ? welem[22] : _GEN_8536; // @[Execute.scala 117:10]
  assign _GEN_8538 = 5'h17 == _T_848 ? welem[23] : _GEN_8537; // @[Execute.scala 117:10]
  assign _GEN_8539 = 5'h18 == _T_848 ? welem[24] : _GEN_8538; // @[Execute.scala 117:10]
  assign _GEN_8540 = 5'h19 == _T_848 ? welem[25] : _GEN_8539; // @[Execute.scala 117:10]
  assign _GEN_8541 = 5'h1a == _T_848 ? welem[26] : _GEN_8540; // @[Execute.scala 117:10]
  assign _GEN_8542 = 5'h1b == _T_848 ? welem[27] : _GEN_8541; // @[Execute.scala 117:10]
  assign _GEN_8543 = 5'h1c == _T_848 ? welem[28] : _GEN_8542; // @[Execute.scala 117:10]
  assign _GEN_8544 = 5'h1d == _T_848 ? welem[29] : _GEN_8543; // @[Execute.scala 117:10]
  assign _GEN_8545 = 5'h1e == _T_848 ? welem[30] : _GEN_8544; // @[Execute.scala 117:10]
  assign _GEN_8546 = 5'h1f == _T_848 ? welem[31] : _GEN_8545; // @[Execute.scala 117:10]
  assign _GEN_8548 = 5'h1 == _T_850 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8549 = 5'h2 == _T_850 ? welem[2] : _GEN_8548; // @[Execute.scala 117:10]
  assign _GEN_8550 = 5'h3 == _T_850 ? welem[3] : _GEN_8549; // @[Execute.scala 117:10]
  assign _GEN_8551 = 5'h4 == _T_850 ? welem[4] : _GEN_8550; // @[Execute.scala 117:10]
  assign _GEN_8552 = 5'h5 == _T_850 ? welem[5] : _GEN_8551; // @[Execute.scala 117:10]
  assign _GEN_8553 = 5'h6 == _T_850 ? welem[6] : _GEN_8552; // @[Execute.scala 117:10]
  assign _GEN_8554 = 5'h7 == _T_850 ? welem[7] : _GEN_8553; // @[Execute.scala 117:10]
  assign _GEN_8555 = 5'h8 == _T_850 ? welem[8] : _GEN_8554; // @[Execute.scala 117:10]
  assign _GEN_8556 = 5'h9 == _T_850 ? welem[9] : _GEN_8555; // @[Execute.scala 117:10]
  assign _GEN_8557 = 5'ha == _T_850 ? welem[10] : _GEN_8556; // @[Execute.scala 117:10]
  assign _GEN_8558 = 5'hb == _T_850 ? welem[11] : _GEN_8557; // @[Execute.scala 117:10]
  assign _GEN_8559 = 5'hc == _T_850 ? welem[12] : _GEN_8558; // @[Execute.scala 117:10]
  assign _GEN_8560 = 5'hd == _T_850 ? welem[13] : _GEN_8559; // @[Execute.scala 117:10]
  assign _GEN_8561 = 5'he == _T_850 ? welem[14] : _GEN_8560; // @[Execute.scala 117:10]
  assign _GEN_8562 = 5'hf == _T_850 ? welem[15] : _GEN_8561; // @[Execute.scala 117:10]
  assign _GEN_8563 = 5'h10 == _T_850 ? welem[16] : _GEN_8562; // @[Execute.scala 117:10]
  assign _GEN_8564 = 5'h11 == _T_850 ? welem[17] : _GEN_8563; // @[Execute.scala 117:10]
  assign _GEN_8565 = 5'h12 == _T_850 ? welem[18] : _GEN_8564; // @[Execute.scala 117:10]
  assign _GEN_8566 = 5'h13 == _T_850 ? welem[19] : _GEN_8565; // @[Execute.scala 117:10]
  assign _GEN_8567 = 5'h14 == _T_850 ? welem[20] : _GEN_8566; // @[Execute.scala 117:10]
  assign _GEN_8568 = 5'h15 == _T_850 ? welem[21] : _GEN_8567; // @[Execute.scala 117:10]
  assign _GEN_8569 = 5'h16 == _T_850 ? welem[22] : _GEN_8568; // @[Execute.scala 117:10]
  assign _GEN_8570 = 5'h17 == _T_850 ? welem[23] : _GEN_8569; // @[Execute.scala 117:10]
  assign _GEN_8571 = 5'h18 == _T_850 ? welem[24] : _GEN_8570; // @[Execute.scala 117:10]
  assign _GEN_8572 = 5'h19 == _T_850 ? welem[25] : _GEN_8571; // @[Execute.scala 117:10]
  assign _GEN_8573 = 5'h1a == _T_850 ? welem[26] : _GEN_8572; // @[Execute.scala 117:10]
  assign _GEN_8574 = 5'h1b == _T_850 ? welem[27] : _GEN_8573; // @[Execute.scala 117:10]
  assign _GEN_8575 = 5'h1c == _T_850 ? welem[28] : _GEN_8574; // @[Execute.scala 117:10]
  assign _GEN_8576 = 5'h1d == _T_850 ? welem[29] : _GEN_8575; // @[Execute.scala 117:10]
  assign _GEN_8577 = 5'h1e == _T_850 ? welem[30] : _GEN_8576; // @[Execute.scala 117:10]
  assign _GEN_8578 = 5'h1f == _T_850 ? welem[31] : _GEN_8577; // @[Execute.scala 117:10]
  assign _T_851 = _T_846 ? _GEN_8546 : _GEN_8578; // @[Execute.scala 117:10]
  assign _T_852 = r[4:0] < 5'h1d; // @[Execute.scala 117:15]
  assign _T_854 = r[4:0] - 5'h1d; // @[Execute.scala 117:37]
  assign _T_856 = 5'h3 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_8580 = 5'h1 == _T_854 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8581 = 5'h2 == _T_854 ? welem[2] : _GEN_8580; // @[Execute.scala 117:10]
  assign _GEN_8582 = 5'h3 == _T_854 ? welem[3] : _GEN_8581; // @[Execute.scala 117:10]
  assign _GEN_8583 = 5'h4 == _T_854 ? welem[4] : _GEN_8582; // @[Execute.scala 117:10]
  assign _GEN_8584 = 5'h5 == _T_854 ? welem[5] : _GEN_8583; // @[Execute.scala 117:10]
  assign _GEN_8585 = 5'h6 == _T_854 ? welem[6] : _GEN_8584; // @[Execute.scala 117:10]
  assign _GEN_8586 = 5'h7 == _T_854 ? welem[7] : _GEN_8585; // @[Execute.scala 117:10]
  assign _GEN_8587 = 5'h8 == _T_854 ? welem[8] : _GEN_8586; // @[Execute.scala 117:10]
  assign _GEN_8588 = 5'h9 == _T_854 ? welem[9] : _GEN_8587; // @[Execute.scala 117:10]
  assign _GEN_8589 = 5'ha == _T_854 ? welem[10] : _GEN_8588; // @[Execute.scala 117:10]
  assign _GEN_8590 = 5'hb == _T_854 ? welem[11] : _GEN_8589; // @[Execute.scala 117:10]
  assign _GEN_8591 = 5'hc == _T_854 ? welem[12] : _GEN_8590; // @[Execute.scala 117:10]
  assign _GEN_8592 = 5'hd == _T_854 ? welem[13] : _GEN_8591; // @[Execute.scala 117:10]
  assign _GEN_8593 = 5'he == _T_854 ? welem[14] : _GEN_8592; // @[Execute.scala 117:10]
  assign _GEN_8594 = 5'hf == _T_854 ? welem[15] : _GEN_8593; // @[Execute.scala 117:10]
  assign _GEN_8595 = 5'h10 == _T_854 ? welem[16] : _GEN_8594; // @[Execute.scala 117:10]
  assign _GEN_8596 = 5'h11 == _T_854 ? welem[17] : _GEN_8595; // @[Execute.scala 117:10]
  assign _GEN_8597 = 5'h12 == _T_854 ? welem[18] : _GEN_8596; // @[Execute.scala 117:10]
  assign _GEN_8598 = 5'h13 == _T_854 ? welem[19] : _GEN_8597; // @[Execute.scala 117:10]
  assign _GEN_8599 = 5'h14 == _T_854 ? welem[20] : _GEN_8598; // @[Execute.scala 117:10]
  assign _GEN_8600 = 5'h15 == _T_854 ? welem[21] : _GEN_8599; // @[Execute.scala 117:10]
  assign _GEN_8601 = 5'h16 == _T_854 ? welem[22] : _GEN_8600; // @[Execute.scala 117:10]
  assign _GEN_8602 = 5'h17 == _T_854 ? welem[23] : _GEN_8601; // @[Execute.scala 117:10]
  assign _GEN_8603 = 5'h18 == _T_854 ? welem[24] : _GEN_8602; // @[Execute.scala 117:10]
  assign _GEN_8604 = 5'h19 == _T_854 ? welem[25] : _GEN_8603; // @[Execute.scala 117:10]
  assign _GEN_8605 = 5'h1a == _T_854 ? welem[26] : _GEN_8604; // @[Execute.scala 117:10]
  assign _GEN_8606 = 5'h1b == _T_854 ? welem[27] : _GEN_8605; // @[Execute.scala 117:10]
  assign _GEN_8607 = 5'h1c == _T_854 ? welem[28] : _GEN_8606; // @[Execute.scala 117:10]
  assign _GEN_8608 = 5'h1d == _T_854 ? welem[29] : _GEN_8607; // @[Execute.scala 117:10]
  assign _GEN_8609 = 5'h1e == _T_854 ? welem[30] : _GEN_8608; // @[Execute.scala 117:10]
  assign _GEN_8610 = 5'h1f == _T_854 ? welem[31] : _GEN_8609; // @[Execute.scala 117:10]
  assign _GEN_8612 = 5'h1 == _T_856 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8613 = 5'h2 == _T_856 ? welem[2] : _GEN_8612; // @[Execute.scala 117:10]
  assign _GEN_8614 = 5'h3 == _T_856 ? welem[3] : _GEN_8613; // @[Execute.scala 117:10]
  assign _GEN_8615 = 5'h4 == _T_856 ? welem[4] : _GEN_8614; // @[Execute.scala 117:10]
  assign _GEN_8616 = 5'h5 == _T_856 ? welem[5] : _GEN_8615; // @[Execute.scala 117:10]
  assign _GEN_8617 = 5'h6 == _T_856 ? welem[6] : _GEN_8616; // @[Execute.scala 117:10]
  assign _GEN_8618 = 5'h7 == _T_856 ? welem[7] : _GEN_8617; // @[Execute.scala 117:10]
  assign _GEN_8619 = 5'h8 == _T_856 ? welem[8] : _GEN_8618; // @[Execute.scala 117:10]
  assign _GEN_8620 = 5'h9 == _T_856 ? welem[9] : _GEN_8619; // @[Execute.scala 117:10]
  assign _GEN_8621 = 5'ha == _T_856 ? welem[10] : _GEN_8620; // @[Execute.scala 117:10]
  assign _GEN_8622 = 5'hb == _T_856 ? welem[11] : _GEN_8621; // @[Execute.scala 117:10]
  assign _GEN_8623 = 5'hc == _T_856 ? welem[12] : _GEN_8622; // @[Execute.scala 117:10]
  assign _GEN_8624 = 5'hd == _T_856 ? welem[13] : _GEN_8623; // @[Execute.scala 117:10]
  assign _GEN_8625 = 5'he == _T_856 ? welem[14] : _GEN_8624; // @[Execute.scala 117:10]
  assign _GEN_8626 = 5'hf == _T_856 ? welem[15] : _GEN_8625; // @[Execute.scala 117:10]
  assign _GEN_8627 = 5'h10 == _T_856 ? welem[16] : _GEN_8626; // @[Execute.scala 117:10]
  assign _GEN_8628 = 5'h11 == _T_856 ? welem[17] : _GEN_8627; // @[Execute.scala 117:10]
  assign _GEN_8629 = 5'h12 == _T_856 ? welem[18] : _GEN_8628; // @[Execute.scala 117:10]
  assign _GEN_8630 = 5'h13 == _T_856 ? welem[19] : _GEN_8629; // @[Execute.scala 117:10]
  assign _GEN_8631 = 5'h14 == _T_856 ? welem[20] : _GEN_8630; // @[Execute.scala 117:10]
  assign _GEN_8632 = 5'h15 == _T_856 ? welem[21] : _GEN_8631; // @[Execute.scala 117:10]
  assign _GEN_8633 = 5'h16 == _T_856 ? welem[22] : _GEN_8632; // @[Execute.scala 117:10]
  assign _GEN_8634 = 5'h17 == _T_856 ? welem[23] : _GEN_8633; // @[Execute.scala 117:10]
  assign _GEN_8635 = 5'h18 == _T_856 ? welem[24] : _GEN_8634; // @[Execute.scala 117:10]
  assign _GEN_8636 = 5'h19 == _T_856 ? welem[25] : _GEN_8635; // @[Execute.scala 117:10]
  assign _GEN_8637 = 5'h1a == _T_856 ? welem[26] : _GEN_8636; // @[Execute.scala 117:10]
  assign _GEN_8638 = 5'h1b == _T_856 ? welem[27] : _GEN_8637; // @[Execute.scala 117:10]
  assign _GEN_8639 = 5'h1c == _T_856 ? welem[28] : _GEN_8638; // @[Execute.scala 117:10]
  assign _GEN_8640 = 5'h1d == _T_856 ? welem[29] : _GEN_8639; // @[Execute.scala 117:10]
  assign _GEN_8641 = 5'h1e == _T_856 ? welem[30] : _GEN_8640; // @[Execute.scala 117:10]
  assign _GEN_8642 = 5'h1f == _T_856 ? welem[31] : _GEN_8641; // @[Execute.scala 117:10]
  assign _T_857 = _T_852 ? _GEN_8610 : _GEN_8642; // @[Execute.scala 117:10]
  assign _T_858 = r[4:0] < 5'h1c; // @[Execute.scala 117:15]
  assign _T_860 = r[4:0] - 5'h1c; // @[Execute.scala 117:37]
  assign _T_862 = 5'h4 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_8644 = 5'h1 == _T_860 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8645 = 5'h2 == _T_860 ? welem[2] : _GEN_8644; // @[Execute.scala 117:10]
  assign _GEN_8646 = 5'h3 == _T_860 ? welem[3] : _GEN_8645; // @[Execute.scala 117:10]
  assign _GEN_8647 = 5'h4 == _T_860 ? welem[4] : _GEN_8646; // @[Execute.scala 117:10]
  assign _GEN_8648 = 5'h5 == _T_860 ? welem[5] : _GEN_8647; // @[Execute.scala 117:10]
  assign _GEN_8649 = 5'h6 == _T_860 ? welem[6] : _GEN_8648; // @[Execute.scala 117:10]
  assign _GEN_8650 = 5'h7 == _T_860 ? welem[7] : _GEN_8649; // @[Execute.scala 117:10]
  assign _GEN_8651 = 5'h8 == _T_860 ? welem[8] : _GEN_8650; // @[Execute.scala 117:10]
  assign _GEN_8652 = 5'h9 == _T_860 ? welem[9] : _GEN_8651; // @[Execute.scala 117:10]
  assign _GEN_8653 = 5'ha == _T_860 ? welem[10] : _GEN_8652; // @[Execute.scala 117:10]
  assign _GEN_8654 = 5'hb == _T_860 ? welem[11] : _GEN_8653; // @[Execute.scala 117:10]
  assign _GEN_8655 = 5'hc == _T_860 ? welem[12] : _GEN_8654; // @[Execute.scala 117:10]
  assign _GEN_8656 = 5'hd == _T_860 ? welem[13] : _GEN_8655; // @[Execute.scala 117:10]
  assign _GEN_8657 = 5'he == _T_860 ? welem[14] : _GEN_8656; // @[Execute.scala 117:10]
  assign _GEN_8658 = 5'hf == _T_860 ? welem[15] : _GEN_8657; // @[Execute.scala 117:10]
  assign _GEN_8659 = 5'h10 == _T_860 ? welem[16] : _GEN_8658; // @[Execute.scala 117:10]
  assign _GEN_8660 = 5'h11 == _T_860 ? welem[17] : _GEN_8659; // @[Execute.scala 117:10]
  assign _GEN_8661 = 5'h12 == _T_860 ? welem[18] : _GEN_8660; // @[Execute.scala 117:10]
  assign _GEN_8662 = 5'h13 == _T_860 ? welem[19] : _GEN_8661; // @[Execute.scala 117:10]
  assign _GEN_8663 = 5'h14 == _T_860 ? welem[20] : _GEN_8662; // @[Execute.scala 117:10]
  assign _GEN_8664 = 5'h15 == _T_860 ? welem[21] : _GEN_8663; // @[Execute.scala 117:10]
  assign _GEN_8665 = 5'h16 == _T_860 ? welem[22] : _GEN_8664; // @[Execute.scala 117:10]
  assign _GEN_8666 = 5'h17 == _T_860 ? welem[23] : _GEN_8665; // @[Execute.scala 117:10]
  assign _GEN_8667 = 5'h18 == _T_860 ? welem[24] : _GEN_8666; // @[Execute.scala 117:10]
  assign _GEN_8668 = 5'h19 == _T_860 ? welem[25] : _GEN_8667; // @[Execute.scala 117:10]
  assign _GEN_8669 = 5'h1a == _T_860 ? welem[26] : _GEN_8668; // @[Execute.scala 117:10]
  assign _GEN_8670 = 5'h1b == _T_860 ? welem[27] : _GEN_8669; // @[Execute.scala 117:10]
  assign _GEN_8671 = 5'h1c == _T_860 ? welem[28] : _GEN_8670; // @[Execute.scala 117:10]
  assign _GEN_8672 = 5'h1d == _T_860 ? welem[29] : _GEN_8671; // @[Execute.scala 117:10]
  assign _GEN_8673 = 5'h1e == _T_860 ? welem[30] : _GEN_8672; // @[Execute.scala 117:10]
  assign _GEN_8674 = 5'h1f == _T_860 ? welem[31] : _GEN_8673; // @[Execute.scala 117:10]
  assign _GEN_8676 = 5'h1 == _T_862 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8677 = 5'h2 == _T_862 ? welem[2] : _GEN_8676; // @[Execute.scala 117:10]
  assign _GEN_8678 = 5'h3 == _T_862 ? welem[3] : _GEN_8677; // @[Execute.scala 117:10]
  assign _GEN_8679 = 5'h4 == _T_862 ? welem[4] : _GEN_8678; // @[Execute.scala 117:10]
  assign _GEN_8680 = 5'h5 == _T_862 ? welem[5] : _GEN_8679; // @[Execute.scala 117:10]
  assign _GEN_8681 = 5'h6 == _T_862 ? welem[6] : _GEN_8680; // @[Execute.scala 117:10]
  assign _GEN_8682 = 5'h7 == _T_862 ? welem[7] : _GEN_8681; // @[Execute.scala 117:10]
  assign _GEN_8683 = 5'h8 == _T_862 ? welem[8] : _GEN_8682; // @[Execute.scala 117:10]
  assign _GEN_8684 = 5'h9 == _T_862 ? welem[9] : _GEN_8683; // @[Execute.scala 117:10]
  assign _GEN_8685 = 5'ha == _T_862 ? welem[10] : _GEN_8684; // @[Execute.scala 117:10]
  assign _GEN_8686 = 5'hb == _T_862 ? welem[11] : _GEN_8685; // @[Execute.scala 117:10]
  assign _GEN_8687 = 5'hc == _T_862 ? welem[12] : _GEN_8686; // @[Execute.scala 117:10]
  assign _GEN_8688 = 5'hd == _T_862 ? welem[13] : _GEN_8687; // @[Execute.scala 117:10]
  assign _GEN_8689 = 5'he == _T_862 ? welem[14] : _GEN_8688; // @[Execute.scala 117:10]
  assign _GEN_8690 = 5'hf == _T_862 ? welem[15] : _GEN_8689; // @[Execute.scala 117:10]
  assign _GEN_8691 = 5'h10 == _T_862 ? welem[16] : _GEN_8690; // @[Execute.scala 117:10]
  assign _GEN_8692 = 5'h11 == _T_862 ? welem[17] : _GEN_8691; // @[Execute.scala 117:10]
  assign _GEN_8693 = 5'h12 == _T_862 ? welem[18] : _GEN_8692; // @[Execute.scala 117:10]
  assign _GEN_8694 = 5'h13 == _T_862 ? welem[19] : _GEN_8693; // @[Execute.scala 117:10]
  assign _GEN_8695 = 5'h14 == _T_862 ? welem[20] : _GEN_8694; // @[Execute.scala 117:10]
  assign _GEN_8696 = 5'h15 == _T_862 ? welem[21] : _GEN_8695; // @[Execute.scala 117:10]
  assign _GEN_8697 = 5'h16 == _T_862 ? welem[22] : _GEN_8696; // @[Execute.scala 117:10]
  assign _GEN_8698 = 5'h17 == _T_862 ? welem[23] : _GEN_8697; // @[Execute.scala 117:10]
  assign _GEN_8699 = 5'h18 == _T_862 ? welem[24] : _GEN_8698; // @[Execute.scala 117:10]
  assign _GEN_8700 = 5'h19 == _T_862 ? welem[25] : _GEN_8699; // @[Execute.scala 117:10]
  assign _GEN_8701 = 5'h1a == _T_862 ? welem[26] : _GEN_8700; // @[Execute.scala 117:10]
  assign _GEN_8702 = 5'h1b == _T_862 ? welem[27] : _GEN_8701; // @[Execute.scala 117:10]
  assign _GEN_8703 = 5'h1c == _T_862 ? welem[28] : _GEN_8702; // @[Execute.scala 117:10]
  assign _GEN_8704 = 5'h1d == _T_862 ? welem[29] : _GEN_8703; // @[Execute.scala 117:10]
  assign _GEN_8705 = 5'h1e == _T_862 ? welem[30] : _GEN_8704; // @[Execute.scala 117:10]
  assign _GEN_8706 = 5'h1f == _T_862 ? welem[31] : _GEN_8705; // @[Execute.scala 117:10]
  assign _T_863 = _T_858 ? _GEN_8674 : _GEN_8706; // @[Execute.scala 117:10]
  assign _T_864 = r[4:0] < 5'h1b; // @[Execute.scala 117:15]
  assign _T_866 = r[4:0] - 5'h1b; // @[Execute.scala 117:37]
  assign _T_868 = 5'h5 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_8708 = 5'h1 == _T_866 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8709 = 5'h2 == _T_866 ? welem[2] : _GEN_8708; // @[Execute.scala 117:10]
  assign _GEN_8710 = 5'h3 == _T_866 ? welem[3] : _GEN_8709; // @[Execute.scala 117:10]
  assign _GEN_8711 = 5'h4 == _T_866 ? welem[4] : _GEN_8710; // @[Execute.scala 117:10]
  assign _GEN_8712 = 5'h5 == _T_866 ? welem[5] : _GEN_8711; // @[Execute.scala 117:10]
  assign _GEN_8713 = 5'h6 == _T_866 ? welem[6] : _GEN_8712; // @[Execute.scala 117:10]
  assign _GEN_8714 = 5'h7 == _T_866 ? welem[7] : _GEN_8713; // @[Execute.scala 117:10]
  assign _GEN_8715 = 5'h8 == _T_866 ? welem[8] : _GEN_8714; // @[Execute.scala 117:10]
  assign _GEN_8716 = 5'h9 == _T_866 ? welem[9] : _GEN_8715; // @[Execute.scala 117:10]
  assign _GEN_8717 = 5'ha == _T_866 ? welem[10] : _GEN_8716; // @[Execute.scala 117:10]
  assign _GEN_8718 = 5'hb == _T_866 ? welem[11] : _GEN_8717; // @[Execute.scala 117:10]
  assign _GEN_8719 = 5'hc == _T_866 ? welem[12] : _GEN_8718; // @[Execute.scala 117:10]
  assign _GEN_8720 = 5'hd == _T_866 ? welem[13] : _GEN_8719; // @[Execute.scala 117:10]
  assign _GEN_8721 = 5'he == _T_866 ? welem[14] : _GEN_8720; // @[Execute.scala 117:10]
  assign _GEN_8722 = 5'hf == _T_866 ? welem[15] : _GEN_8721; // @[Execute.scala 117:10]
  assign _GEN_8723 = 5'h10 == _T_866 ? welem[16] : _GEN_8722; // @[Execute.scala 117:10]
  assign _GEN_8724 = 5'h11 == _T_866 ? welem[17] : _GEN_8723; // @[Execute.scala 117:10]
  assign _GEN_8725 = 5'h12 == _T_866 ? welem[18] : _GEN_8724; // @[Execute.scala 117:10]
  assign _GEN_8726 = 5'h13 == _T_866 ? welem[19] : _GEN_8725; // @[Execute.scala 117:10]
  assign _GEN_8727 = 5'h14 == _T_866 ? welem[20] : _GEN_8726; // @[Execute.scala 117:10]
  assign _GEN_8728 = 5'h15 == _T_866 ? welem[21] : _GEN_8727; // @[Execute.scala 117:10]
  assign _GEN_8729 = 5'h16 == _T_866 ? welem[22] : _GEN_8728; // @[Execute.scala 117:10]
  assign _GEN_8730 = 5'h17 == _T_866 ? welem[23] : _GEN_8729; // @[Execute.scala 117:10]
  assign _GEN_8731 = 5'h18 == _T_866 ? welem[24] : _GEN_8730; // @[Execute.scala 117:10]
  assign _GEN_8732 = 5'h19 == _T_866 ? welem[25] : _GEN_8731; // @[Execute.scala 117:10]
  assign _GEN_8733 = 5'h1a == _T_866 ? welem[26] : _GEN_8732; // @[Execute.scala 117:10]
  assign _GEN_8734 = 5'h1b == _T_866 ? welem[27] : _GEN_8733; // @[Execute.scala 117:10]
  assign _GEN_8735 = 5'h1c == _T_866 ? welem[28] : _GEN_8734; // @[Execute.scala 117:10]
  assign _GEN_8736 = 5'h1d == _T_866 ? welem[29] : _GEN_8735; // @[Execute.scala 117:10]
  assign _GEN_8737 = 5'h1e == _T_866 ? welem[30] : _GEN_8736; // @[Execute.scala 117:10]
  assign _GEN_8738 = 5'h1f == _T_866 ? welem[31] : _GEN_8737; // @[Execute.scala 117:10]
  assign _GEN_8740 = 5'h1 == _T_868 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8741 = 5'h2 == _T_868 ? welem[2] : _GEN_8740; // @[Execute.scala 117:10]
  assign _GEN_8742 = 5'h3 == _T_868 ? welem[3] : _GEN_8741; // @[Execute.scala 117:10]
  assign _GEN_8743 = 5'h4 == _T_868 ? welem[4] : _GEN_8742; // @[Execute.scala 117:10]
  assign _GEN_8744 = 5'h5 == _T_868 ? welem[5] : _GEN_8743; // @[Execute.scala 117:10]
  assign _GEN_8745 = 5'h6 == _T_868 ? welem[6] : _GEN_8744; // @[Execute.scala 117:10]
  assign _GEN_8746 = 5'h7 == _T_868 ? welem[7] : _GEN_8745; // @[Execute.scala 117:10]
  assign _GEN_8747 = 5'h8 == _T_868 ? welem[8] : _GEN_8746; // @[Execute.scala 117:10]
  assign _GEN_8748 = 5'h9 == _T_868 ? welem[9] : _GEN_8747; // @[Execute.scala 117:10]
  assign _GEN_8749 = 5'ha == _T_868 ? welem[10] : _GEN_8748; // @[Execute.scala 117:10]
  assign _GEN_8750 = 5'hb == _T_868 ? welem[11] : _GEN_8749; // @[Execute.scala 117:10]
  assign _GEN_8751 = 5'hc == _T_868 ? welem[12] : _GEN_8750; // @[Execute.scala 117:10]
  assign _GEN_8752 = 5'hd == _T_868 ? welem[13] : _GEN_8751; // @[Execute.scala 117:10]
  assign _GEN_8753 = 5'he == _T_868 ? welem[14] : _GEN_8752; // @[Execute.scala 117:10]
  assign _GEN_8754 = 5'hf == _T_868 ? welem[15] : _GEN_8753; // @[Execute.scala 117:10]
  assign _GEN_8755 = 5'h10 == _T_868 ? welem[16] : _GEN_8754; // @[Execute.scala 117:10]
  assign _GEN_8756 = 5'h11 == _T_868 ? welem[17] : _GEN_8755; // @[Execute.scala 117:10]
  assign _GEN_8757 = 5'h12 == _T_868 ? welem[18] : _GEN_8756; // @[Execute.scala 117:10]
  assign _GEN_8758 = 5'h13 == _T_868 ? welem[19] : _GEN_8757; // @[Execute.scala 117:10]
  assign _GEN_8759 = 5'h14 == _T_868 ? welem[20] : _GEN_8758; // @[Execute.scala 117:10]
  assign _GEN_8760 = 5'h15 == _T_868 ? welem[21] : _GEN_8759; // @[Execute.scala 117:10]
  assign _GEN_8761 = 5'h16 == _T_868 ? welem[22] : _GEN_8760; // @[Execute.scala 117:10]
  assign _GEN_8762 = 5'h17 == _T_868 ? welem[23] : _GEN_8761; // @[Execute.scala 117:10]
  assign _GEN_8763 = 5'h18 == _T_868 ? welem[24] : _GEN_8762; // @[Execute.scala 117:10]
  assign _GEN_8764 = 5'h19 == _T_868 ? welem[25] : _GEN_8763; // @[Execute.scala 117:10]
  assign _GEN_8765 = 5'h1a == _T_868 ? welem[26] : _GEN_8764; // @[Execute.scala 117:10]
  assign _GEN_8766 = 5'h1b == _T_868 ? welem[27] : _GEN_8765; // @[Execute.scala 117:10]
  assign _GEN_8767 = 5'h1c == _T_868 ? welem[28] : _GEN_8766; // @[Execute.scala 117:10]
  assign _GEN_8768 = 5'h1d == _T_868 ? welem[29] : _GEN_8767; // @[Execute.scala 117:10]
  assign _GEN_8769 = 5'h1e == _T_868 ? welem[30] : _GEN_8768; // @[Execute.scala 117:10]
  assign _GEN_8770 = 5'h1f == _T_868 ? welem[31] : _GEN_8769; // @[Execute.scala 117:10]
  assign _T_869 = _T_864 ? _GEN_8738 : _GEN_8770; // @[Execute.scala 117:10]
  assign _T_870 = r[4:0] < 5'h1a; // @[Execute.scala 117:15]
  assign _T_872 = r[4:0] - 5'h1a; // @[Execute.scala 117:37]
  assign _T_874 = 5'h6 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_8772 = 5'h1 == _T_872 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8773 = 5'h2 == _T_872 ? welem[2] : _GEN_8772; // @[Execute.scala 117:10]
  assign _GEN_8774 = 5'h3 == _T_872 ? welem[3] : _GEN_8773; // @[Execute.scala 117:10]
  assign _GEN_8775 = 5'h4 == _T_872 ? welem[4] : _GEN_8774; // @[Execute.scala 117:10]
  assign _GEN_8776 = 5'h5 == _T_872 ? welem[5] : _GEN_8775; // @[Execute.scala 117:10]
  assign _GEN_8777 = 5'h6 == _T_872 ? welem[6] : _GEN_8776; // @[Execute.scala 117:10]
  assign _GEN_8778 = 5'h7 == _T_872 ? welem[7] : _GEN_8777; // @[Execute.scala 117:10]
  assign _GEN_8779 = 5'h8 == _T_872 ? welem[8] : _GEN_8778; // @[Execute.scala 117:10]
  assign _GEN_8780 = 5'h9 == _T_872 ? welem[9] : _GEN_8779; // @[Execute.scala 117:10]
  assign _GEN_8781 = 5'ha == _T_872 ? welem[10] : _GEN_8780; // @[Execute.scala 117:10]
  assign _GEN_8782 = 5'hb == _T_872 ? welem[11] : _GEN_8781; // @[Execute.scala 117:10]
  assign _GEN_8783 = 5'hc == _T_872 ? welem[12] : _GEN_8782; // @[Execute.scala 117:10]
  assign _GEN_8784 = 5'hd == _T_872 ? welem[13] : _GEN_8783; // @[Execute.scala 117:10]
  assign _GEN_8785 = 5'he == _T_872 ? welem[14] : _GEN_8784; // @[Execute.scala 117:10]
  assign _GEN_8786 = 5'hf == _T_872 ? welem[15] : _GEN_8785; // @[Execute.scala 117:10]
  assign _GEN_8787 = 5'h10 == _T_872 ? welem[16] : _GEN_8786; // @[Execute.scala 117:10]
  assign _GEN_8788 = 5'h11 == _T_872 ? welem[17] : _GEN_8787; // @[Execute.scala 117:10]
  assign _GEN_8789 = 5'h12 == _T_872 ? welem[18] : _GEN_8788; // @[Execute.scala 117:10]
  assign _GEN_8790 = 5'h13 == _T_872 ? welem[19] : _GEN_8789; // @[Execute.scala 117:10]
  assign _GEN_8791 = 5'h14 == _T_872 ? welem[20] : _GEN_8790; // @[Execute.scala 117:10]
  assign _GEN_8792 = 5'h15 == _T_872 ? welem[21] : _GEN_8791; // @[Execute.scala 117:10]
  assign _GEN_8793 = 5'h16 == _T_872 ? welem[22] : _GEN_8792; // @[Execute.scala 117:10]
  assign _GEN_8794 = 5'h17 == _T_872 ? welem[23] : _GEN_8793; // @[Execute.scala 117:10]
  assign _GEN_8795 = 5'h18 == _T_872 ? welem[24] : _GEN_8794; // @[Execute.scala 117:10]
  assign _GEN_8796 = 5'h19 == _T_872 ? welem[25] : _GEN_8795; // @[Execute.scala 117:10]
  assign _GEN_8797 = 5'h1a == _T_872 ? welem[26] : _GEN_8796; // @[Execute.scala 117:10]
  assign _GEN_8798 = 5'h1b == _T_872 ? welem[27] : _GEN_8797; // @[Execute.scala 117:10]
  assign _GEN_8799 = 5'h1c == _T_872 ? welem[28] : _GEN_8798; // @[Execute.scala 117:10]
  assign _GEN_8800 = 5'h1d == _T_872 ? welem[29] : _GEN_8799; // @[Execute.scala 117:10]
  assign _GEN_8801 = 5'h1e == _T_872 ? welem[30] : _GEN_8800; // @[Execute.scala 117:10]
  assign _GEN_8802 = 5'h1f == _T_872 ? welem[31] : _GEN_8801; // @[Execute.scala 117:10]
  assign _GEN_8804 = 5'h1 == _T_874 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8805 = 5'h2 == _T_874 ? welem[2] : _GEN_8804; // @[Execute.scala 117:10]
  assign _GEN_8806 = 5'h3 == _T_874 ? welem[3] : _GEN_8805; // @[Execute.scala 117:10]
  assign _GEN_8807 = 5'h4 == _T_874 ? welem[4] : _GEN_8806; // @[Execute.scala 117:10]
  assign _GEN_8808 = 5'h5 == _T_874 ? welem[5] : _GEN_8807; // @[Execute.scala 117:10]
  assign _GEN_8809 = 5'h6 == _T_874 ? welem[6] : _GEN_8808; // @[Execute.scala 117:10]
  assign _GEN_8810 = 5'h7 == _T_874 ? welem[7] : _GEN_8809; // @[Execute.scala 117:10]
  assign _GEN_8811 = 5'h8 == _T_874 ? welem[8] : _GEN_8810; // @[Execute.scala 117:10]
  assign _GEN_8812 = 5'h9 == _T_874 ? welem[9] : _GEN_8811; // @[Execute.scala 117:10]
  assign _GEN_8813 = 5'ha == _T_874 ? welem[10] : _GEN_8812; // @[Execute.scala 117:10]
  assign _GEN_8814 = 5'hb == _T_874 ? welem[11] : _GEN_8813; // @[Execute.scala 117:10]
  assign _GEN_8815 = 5'hc == _T_874 ? welem[12] : _GEN_8814; // @[Execute.scala 117:10]
  assign _GEN_8816 = 5'hd == _T_874 ? welem[13] : _GEN_8815; // @[Execute.scala 117:10]
  assign _GEN_8817 = 5'he == _T_874 ? welem[14] : _GEN_8816; // @[Execute.scala 117:10]
  assign _GEN_8818 = 5'hf == _T_874 ? welem[15] : _GEN_8817; // @[Execute.scala 117:10]
  assign _GEN_8819 = 5'h10 == _T_874 ? welem[16] : _GEN_8818; // @[Execute.scala 117:10]
  assign _GEN_8820 = 5'h11 == _T_874 ? welem[17] : _GEN_8819; // @[Execute.scala 117:10]
  assign _GEN_8821 = 5'h12 == _T_874 ? welem[18] : _GEN_8820; // @[Execute.scala 117:10]
  assign _GEN_8822 = 5'h13 == _T_874 ? welem[19] : _GEN_8821; // @[Execute.scala 117:10]
  assign _GEN_8823 = 5'h14 == _T_874 ? welem[20] : _GEN_8822; // @[Execute.scala 117:10]
  assign _GEN_8824 = 5'h15 == _T_874 ? welem[21] : _GEN_8823; // @[Execute.scala 117:10]
  assign _GEN_8825 = 5'h16 == _T_874 ? welem[22] : _GEN_8824; // @[Execute.scala 117:10]
  assign _GEN_8826 = 5'h17 == _T_874 ? welem[23] : _GEN_8825; // @[Execute.scala 117:10]
  assign _GEN_8827 = 5'h18 == _T_874 ? welem[24] : _GEN_8826; // @[Execute.scala 117:10]
  assign _GEN_8828 = 5'h19 == _T_874 ? welem[25] : _GEN_8827; // @[Execute.scala 117:10]
  assign _GEN_8829 = 5'h1a == _T_874 ? welem[26] : _GEN_8828; // @[Execute.scala 117:10]
  assign _GEN_8830 = 5'h1b == _T_874 ? welem[27] : _GEN_8829; // @[Execute.scala 117:10]
  assign _GEN_8831 = 5'h1c == _T_874 ? welem[28] : _GEN_8830; // @[Execute.scala 117:10]
  assign _GEN_8832 = 5'h1d == _T_874 ? welem[29] : _GEN_8831; // @[Execute.scala 117:10]
  assign _GEN_8833 = 5'h1e == _T_874 ? welem[30] : _GEN_8832; // @[Execute.scala 117:10]
  assign _GEN_8834 = 5'h1f == _T_874 ? welem[31] : _GEN_8833; // @[Execute.scala 117:10]
  assign _T_875 = _T_870 ? _GEN_8802 : _GEN_8834; // @[Execute.scala 117:10]
  assign _T_876 = r[4:0] < 5'h19; // @[Execute.scala 117:15]
  assign _T_878 = r[4:0] - 5'h19; // @[Execute.scala 117:37]
  assign _T_880 = 5'h7 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_8836 = 5'h1 == _T_878 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8837 = 5'h2 == _T_878 ? welem[2] : _GEN_8836; // @[Execute.scala 117:10]
  assign _GEN_8838 = 5'h3 == _T_878 ? welem[3] : _GEN_8837; // @[Execute.scala 117:10]
  assign _GEN_8839 = 5'h4 == _T_878 ? welem[4] : _GEN_8838; // @[Execute.scala 117:10]
  assign _GEN_8840 = 5'h5 == _T_878 ? welem[5] : _GEN_8839; // @[Execute.scala 117:10]
  assign _GEN_8841 = 5'h6 == _T_878 ? welem[6] : _GEN_8840; // @[Execute.scala 117:10]
  assign _GEN_8842 = 5'h7 == _T_878 ? welem[7] : _GEN_8841; // @[Execute.scala 117:10]
  assign _GEN_8843 = 5'h8 == _T_878 ? welem[8] : _GEN_8842; // @[Execute.scala 117:10]
  assign _GEN_8844 = 5'h9 == _T_878 ? welem[9] : _GEN_8843; // @[Execute.scala 117:10]
  assign _GEN_8845 = 5'ha == _T_878 ? welem[10] : _GEN_8844; // @[Execute.scala 117:10]
  assign _GEN_8846 = 5'hb == _T_878 ? welem[11] : _GEN_8845; // @[Execute.scala 117:10]
  assign _GEN_8847 = 5'hc == _T_878 ? welem[12] : _GEN_8846; // @[Execute.scala 117:10]
  assign _GEN_8848 = 5'hd == _T_878 ? welem[13] : _GEN_8847; // @[Execute.scala 117:10]
  assign _GEN_8849 = 5'he == _T_878 ? welem[14] : _GEN_8848; // @[Execute.scala 117:10]
  assign _GEN_8850 = 5'hf == _T_878 ? welem[15] : _GEN_8849; // @[Execute.scala 117:10]
  assign _GEN_8851 = 5'h10 == _T_878 ? welem[16] : _GEN_8850; // @[Execute.scala 117:10]
  assign _GEN_8852 = 5'h11 == _T_878 ? welem[17] : _GEN_8851; // @[Execute.scala 117:10]
  assign _GEN_8853 = 5'h12 == _T_878 ? welem[18] : _GEN_8852; // @[Execute.scala 117:10]
  assign _GEN_8854 = 5'h13 == _T_878 ? welem[19] : _GEN_8853; // @[Execute.scala 117:10]
  assign _GEN_8855 = 5'h14 == _T_878 ? welem[20] : _GEN_8854; // @[Execute.scala 117:10]
  assign _GEN_8856 = 5'h15 == _T_878 ? welem[21] : _GEN_8855; // @[Execute.scala 117:10]
  assign _GEN_8857 = 5'h16 == _T_878 ? welem[22] : _GEN_8856; // @[Execute.scala 117:10]
  assign _GEN_8858 = 5'h17 == _T_878 ? welem[23] : _GEN_8857; // @[Execute.scala 117:10]
  assign _GEN_8859 = 5'h18 == _T_878 ? welem[24] : _GEN_8858; // @[Execute.scala 117:10]
  assign _GEN_8860 = 5'h19 == _T_878 ? welem[25] : _GEN_8859; // @[Execute.scala 117:10]
  assign _GEN_8861 = 5'h1a == _T_878 ? welem[26] : _GEN_8860; // @[Execute.scala 117:10]
  assign _GEN_8862 = 5'h1b == _T_878 ? welem[27] : _GEN_8861; // @[Execute.scala 117:10]
  assign _GEN_8863 = 5'h1c == _T_878 ? welem[28] : _GEN_8862; // @[Execute.scala 117:10]
  assign _GEN_8864 = 5'h1d == _T_878 ? welem[29] : _GEN_8863; // @[Execute.scala 117:10]
  assign _GEN_8865 = 5'h1e == _T_878 ? welem[30] : _GEN_8864; // @[Execute.scala 117:10]
  assign _GEN_8866 = 5'h1f == _T_878 ? welem[31] : _GEN_8865; // @[Execute.scala 117:10]
  assign _GEN_8868 = 5'h1 == _T_880 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8869 = 5'h2 == _T_880 ? welem[2] : _GEN_8868; // @[Execute.scala 117:10]
  assign _GEN_8870 = 5'h3 == _T_880 ? welem[3] : _GEN_8869; // @[Execute.scala 117:10]
  assign _GEN_8871 = 5'h4 == _T_880 ? welem[4] : _GEN_8870; // @[Execute.scala 117:10]
  assign _GEN_8872 = 5'h5 == _T_880 ? welem[5] : _GEN_8871; // @[Execute.scala 117:10]
  assign _GEN_8873 = 5'h6 == _T_880 ? welem[6] : _GEN_8872; // @[Execute.scala 117:10]
  assign _GEN_8874 = 5'h7 == _T_880 ? welem[7] : _GEN_8873; // @[Execute.scala 117:10]
  assign _GEN_8875 = 5'h8 == _T_880 ? welem[8] : _GEN_8874; // @[Execute.scala 117:10]
  assign _GEN_8876 = 5'h9 == _T_880 ? welem[9] : _GEN_8875; // @[Execute.scala 117:10]
  assign _GEN_8877 = 5'ha == _T_880 ? welem[10] : _GEN_8876; // @[Execute.scala 117:10]
  assign _GEN_8878 = 5'hb == _T_880 ? welem[11] : _GEN_8877; // @[Execute.scala 117:10]
  assign _GEN_8879 = 5'hc == _T_880 ? welem[12] : _GEN_8878; // @[Execute.scala 117:10]
  assign _GEN_8880 = 5'hd == _T_880 ? welem[13] : _GEN_8879; // @[Execute.scala 117:10]
  assign _GEN_8881 = 5'he == _T_880 ? welem[14] : _GEN_8880; // @[Execute.scala 117:10]
  assign _GEN_8882 = 5'hf == _T_880 ? welem[15] : _GEN_8881; // @[Execute.scala 117:10]
  assign _GEN_8883 = 5'h10 == _T_880 ? welem[16] : _GEN_8882; // @[Execute.scala 117:10]
  assign _GEN_8884 = 5'h11 == _T_880 ? welem[17] : _GEN_8883; // @[Execute.scala 117:10]
  assign _GEN_8885 = 5'h12 == _T_880 ? welem[18] : _GEN_8884; // @[Execute.scala 117:10]
  assign _GEN_8886 = 5'h13 == _T_880 ? welem[19] : _GEN_8885; // @[Execute.scala 117:10]
  assign _GEN_8887 = 5'h14 == _T_880 ? welem[20] : _GEN_8886; // @[Execute.scala 117:10]
  assign _GEN_8888 = 5'h15 == _T_880 ? welem[21] : _GEN_8887; // @[Execute.scala 117:10]
  assign _GEN_8889 = 5'h16 == _T_880 ? welem[22] : _GEN_8888; // @[Execute.scala 117:10]
  assign _GEN_8890 = 5'h17 == _T_880 ? welem[23] : _GEN_8889; // @[Execute.scala 117:10]
  assign _GEN_8891 = 5'h18 == _T_880 ? welem[24] : _GEN_8890; // @[Execute.scala 117:10]
  assign _GEN_8892 = 5'h19 == _T_880 ? welem[25] : _GEN_8891; // @[Execute.scala 117:10]
  assign _GEN_8893 = 5'h1a == _T_880 ? welem[26] : _GEN_8892; // @[Execute.scala 117:10]
  assign _GEN_8894 = 5'h1b == _T_880 ? welem[27] : _GEN_8893; // @[Execute.scala 117:10]
  assign _GEN_8895 = 5'h1c == _T_880 ? welem[28] : _GEN_8894; // @[Execute.scala 117:10]
  assign _GEN_8896 = 5'h1d == _T_880 ? welem[29] : _GEN_8895; // @[Execute.scala 117:10]
  assign _GEN_8897 = 5'h1e == _T_880 ? welem[30] : _GEN_8896; // @[Execute.scala 117:10]
  assign _GEN_8898 = 5'h1f == _T_880 ? welem[31] : _GEN_8897; // @[Execute.scala 117:10]
  assign _T_881 = _T_876 ? _GEN_8866 : _GEN_8898; // @[Execute.scala 117:10]
  assign _T_882 = r[4:0] < 5'h18; // @[Execute.scala 117:15]
  assign _T_884 = r[4:0] - 5'h18; // @[Execute.scala 117:37]
  assign _T_886 = 5'h8 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_8900 = 5'h1 == _T_884 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8901 = 5'h2 == _T_884 ? welem[2] : _GEN_8900; // @[Execute.scala 117:10]
  assign _GEN_8902 = 5'h3 == _T_884 ? welem[3] : _GEN_8901; // @[Execute.scala 117:10]
  assign _GEN_8903 = 5'h4 == _T_884 ? welem[4] : _GEN_8902; // @[Execute.scala 117:10]
  assign _GEN_8904 = 5'h5 == _T_884 ? welem[5] : _GEN_8903; // @[Execute.scala 117:10]
  assign _GEN_8905 = 5'h6 == _T_884 ? welem[6] : _GEN_8904; // @[Execute.scala 117:10]
  assign _GEN_8906 = 5'h7 == _T_884 ? welem[7] : _GEN_8905; // @[Execute.scala 117:10]
  assign _GEN_8907 = 5'h8 == _T_884 ? welem[8] : _GEN_8906; // @[Execute.scala 117:10]
  assign _GEN_8908 = 5'h9 == _T_884 ? welem[9] : _GEN_8907; // @[Execute.scala 117:10]
  assign _GEN_8909 = 5'ha == _T_884 ? welem[10] : _GEN_8908; // @[Execute.scala 117:10]
  assign _GEN_8910 = 5'hb == _T_884 ? welem[11] : _GEN_8909; // @[Execute.scala 117:10]
  assign _GEN_8911 = 5'hc == _T_884 ? welem[12] : _GEN_8910; // @[Execute.scala 117:10]
  assign _GEN_8912 = 5'hd == _T_884 ? welem[13] : _GEN_8911; // @[Execute.scala 117:10]
  assign _GEN_8913 = 5'he == _T_884 ? welem[14] : _GEN_8912; // @[Execute.scala 117:10]
  assign _GEN_8914 = 5'hf == _T_884 ? welem[15] : _GEN_8913; // @[Execute.scala 117:10]
  assign _GEN_8915 = 5'h10 == _T_884 ? welem[16] : _GEN_8914; // @[Execute.scala 117:10]
  assign _GEN_8916 = 5'h11 == _T_884 ? welem[17] : _GEN_8915; // @[Execute.scala 117:10]
  assign _GEN_8917 = 5'h12 == _T_884 ? welem[18] : _GEN_8916; // @[Execute.scala 117:10]
  assign _GEN_8918 = 5'h13 == _T_884 ? welem[19] : _GEN_8917; // @[Execute.scala 117:10]
  assign _GEN_8919 = 5'h14 == _T_884 ? welem[20] : _GEN_8918; // @[Execute.scala 117:10]
  assign _GEN_8920 = 5'h15 == _T_884 ? welem[21] : _GEN_8919; // @[Execute.scala 117:10]
  assign _GEN_8921 = 5'h16 == _T_884 ? welem[22] : _GEN_8920; // @[Execute.scala 117:10]
  assign _GEN_8922 = 5'h17 == _T_884 ? welem[23] : _GEN_8921; // @[Execute.scala 117:10]
  assign _GEN_8923 = 5'h18 == _T_884 ? welem[24] : _GEN_8922; // @[Execute.scala 117:10]
  assign _GEN_8924 = 5'h19 == _T_884 ? welem[25] : _GEN_8923; // @[Execute.scala 117:10]
  assign _GEN_8925 = 5'h1a == _T_884 ? welem[26] : _GEN_8924; // @[Execute.scala 117:10]
  assign _GEN_8926 = 5'h1b == _T_884 ? welem[27] : _GEN_8925; // @[Execute.scala 117:10]
  assign _GEN_8927 = 5'h1c == _T_884 ? welem[28] : _GEN_8926; // @[Execute.scala 117:10]
  assign _GEN_8928 = 5'h1d == _T_884 ? welem[29] : _GEN_8927; // @[Execute.scala 117:10]
  assign _GEN_8929 = 5'h1e == _T_884 ? welem[30] : _GEN_8928; // @[Execute.scala 117:10]
  assign _GEN_8930 = 5'h1f == _T_884 ? welem[31] : _GEN_8929; // @[Execute.scala 117:10]
  assign _GEN_8932 = 5'h1 == _T_886 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8933 = 5'h2 == _T_886 ? welem[2] : _GEN_8932; // @[Execute.scala 117:10]
  assign _GEN_8934 = 5'h3 == _T_886 ? welem[3] : _GEN_8933; // @[Execute.scala 117:10]
  assign _GEN_8935 = 5'h4 == _T_886 ? welem[4] : _GEN_8934; // @[Execute.scala 117:10]
  assign _GEN_8936 = 5'h5 == _T_886 ? welem[5] : _GEN_8935; // @[Execute.scala 117:10]
  assign _GEN_8937 = 5'h6 == _T_886 ? welem[6] : _GEN_8936; // @[Execute.scala 117:10]
  assign _GEN_8938 = 5'h7 == _T_886 ? welem[7] : _GEN_8937; // @[Execute.scala 117:10]
  assign _GEN_8939 = 5'h8 == _T_886 ? welem[8] : _GEN_8938; // @[Execute.scala 117:10]
  assign _GEN_8940 = 5'h9 == _T_886 ? welem[9] : _GEN_8939; // @[Execute.scala 117:10]
  assign _GEN_8941 = 5'ha == _T_886 ? welem[10] : _GEN_8940; // @[Execute.scala 117:10]
  assign _GEN_8942 = 5'hb == _T_886 ? welem[11] : _GEN_8941; // @[Execute.scala 117:10]
  assign _GEN_8943 = 5'hc == _T_886 ? welem[12] : _GEN_8942; // @[Execute.scala 117:10]
  assign _GEN_8944 = 5'hd == _T_886 ? welem[13] : _GEN_8943; // @[Execute.scala 117:10]
  assign _GEN_8945 = 5'he == _T_886 ? welem[14] : _GEN_8944; // @[Execute.scala 117:10]
  assign _GEN_8946 = 5'hf == _T_886 ? welem[15] : _GEN_8945; // @[Execute.scala 117:10]
  assign _GEN_8947 = 5'h10 == _T_886 ? welem[16] : _GEN_8946; // @[Execute.scala 117:10]
  assign _GEN_8948 = 5'h11 == _T_886 ? welem[17] : _GEN_8947; // @[Execute.scala 117:10]
  assign _GEN_8949 = 5'h12 == _T_886 ? welem[18] : _GEN_8948; // @[Execute.scala 117:10]
  assign _GEN_8950 = 5'h13 == _T_886 ? welem[19] : _GEN_8949; // @[Execute.scala 117:10]
  assign _GEN_8951 = 5'h14 == _T_886 ? welem[20] : _GEN_8950; // @[Execute.scala 117:10]
  assign _GEN_8952 = 5'h15 == _T_886 ? welem[21] : _GEN_8951; // @[Execute.scala 117:10]
  assign _GEN_8953 = 5'h16 == _T_886 ? welem[22] : _GEN_8952; // @[Execute.scala 117:10]
  assign _GEN_8954 = 5'h17 == _T_886 ? welem[23] : _GEN_8953; // @[Execute.scala 117:10]
  assign _GEN_8955 = 5'h18 == _T_886 ? welem[24] : _GEN_8954; // @[Execute.scala 117:10]
  assign _GEN_8956 = 5'h19 == _T_886 ? welem[25] : _GEN_8955; // @[Execute.scala 117:10]
  assign _GEN_8957 = 5'h1a == _T_886 ? welem[26] : _GEN_8956; // @[Execute.scala 117:10]
  assign _GEN_8958 = 5'h1b == _T_886 ? welem[27] : _GEN_8957; // @[Execute.scala 117:10]
  assign _GEN_8959 = 5'h1c == _T_886 ? welem[28] : _GEN_8958; // @[Execute.scala 117:10]
  assign _GEN_8960 = 5'h1d == _T_886 ? welem[29] : _GEN_8959; // @[Execute.scala 117:10]
  assign _GEN_8961 = 5'h1e == _T_886 ? welem[30] : _GEN_8960; // @[Execute.scala 117:10]
  assign _GEN_8962 = 5'h1f == _T_886 ? welem[31] : _GEN_8961; // @[Execute.scala 117:10]
  assign _T_887 = _T_882 ? _GEN_8930 : _GEN_8962; // @[Execute.scala 117:10]
  assign _T_888 = r[4:0] < 5'h17; // @[Execute.scala 117:15]
  assign _T_890 = r[4:0] - 5'h17; // @[Execute.scala 117:37]
  assign _T_892 = 5'h9 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_8964 = 5'h1 == _T_890 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8965 = 5'h2 == _T_890 ? welem[2] : _GEN_8964; // @[Execute.scala 117:10]
  assign _GEN_8966 = 5'h3 == _T_890 ? welem[3] : _GEN_8965; // @[Execute.scala 117:10]
  assign _GEN_8967 = 5'h4 == _T_890 ? welem[4] : _GEN_8966; // @[Execute.scala 117:10]
  assign _GEN_8968 = 5'h5 == _T_890 ? welem[5] : _GEN_8967; // @[Execute.scala 117:10]
  assign _GEN_8969 = 5'h6 == _T_890 ? welem[6] : _GEN_8968; // @[Execute.scala 117:10]
  assign _GEN_8970 = 5'h7 == _T_890 ? welem[7] : _GEN_8969; // @[Execute.scala 117:10]
  assign _GEN_8971 = 5'h8 == _T_890 ? welem[8] : _GEN_8970; // @[Execute.scala 117:10]
  assign _GEN_8972 = 5'h9 == _T_890 ? welem[9] : _GEN_8971; // @[Execute.scala 117:10]
  assign _GEN_8973 = 5'ha == _T_890 ? welem[10] : _GEN_8972; // @[Execute.scala 117:10]
  assign _GEN_8974 = 5'hb == _T_890 ? welem[11] : _GEN_8973; // @[Execute.scala 117:10]
  assign _GEN_8975 = 5'hc == _T_890 ? welem[12] : _GEN_8974; // @[Execute.scala 117:10]
  assign _GEN_8976 = 5'hd == _T_890 ? welem[13] : _GEN_8975; // @[Execute.scala 117:10]
  assign _GEN_8977 = 5'he == _T_890 ? welem[14] : _GEN_8976; // @[Execute.scala 117:10]
  assign _GEN_8978 = 5'hf == _T_890 ? welem[15] : _GEN_8977; // @[Execute.scala 117:10]
  assign _GEN_8979 = 5'h10 == _T_890 ? welem[16] : _GEN_8978; // @[Execute.scala 117:10]
  assign _GEN_8980 = 5'h11 == _T_890 ? welem[17] : _GEN_8979; // @[Execute.scala 117:10]
  assign _GEN_8981 = 5'h12 == _T_890 ? welem[18] : _GEN_8980; // @[Execute.scala 117:10]
  assign _GEN_8982 = 5'h13 == _T_890 ? welem[19] : _GEN_8981; // @[Execute.scala 117:10]
  assign _GEN_8983 = 5'h14 == _T_890 ? welem[20] : _GEN_8982; // @[Execute.scala 117:10]
  assign _GEN_8984 = 5'h15 == _T_890 ? welem[21] : _GEN_8983; // @[Execute.scala 117:10]
  assign _GEN_8985 = 5'h16 == _T_890 ? welem[22] : _GEN_8984; // @[Execute.scala 117:10]
  assign _GEN_8986 = 5'h17 == _T_890 ? welem[23] : _GEN_8985; // @[Execute.scala 117:10]
  assign _GEN_8987 = 5'h18 == _T_890 ? welem[24] : _GEN_8986; // @[Execute.scala 117:10]
  assign _GEN_8988 = 5'h19 == _T_890 ? welem[25] : _GEN_8987; // @[Execute.scala 117:10]
  assign _GEN_8989 = 5'h1a == _T_890 ? welem[26] : _GEN_8988; // @[Execute.scala 117:10]
  assign _GEN_8990 = 5'h1b == _T_890 ? welem[27] : _GEN_8989; // @[Execute.scala 117:10]
  assign _GEN_8991 = 5'h1c == _T_890 ? welem[28] : _GEN_8990; // @[Execute.scala 117:10]
  assign _GEN_8992 = 5'h1d == _T_890 ? welem[29] : _GEN_8991; // @[Execute.scala 117:10]
  assign _GEN_8993 = 5'h1e == _T_890 ? welem[30] : _GEN_8992; // @[Execute.scala 117:10]
  assign _GEN_8994 = 5'h1f == _T_890 ? welem[31] : _GEN_8993; // @[Execute.scala 117:10]
  assign _GEN_8996 = 5'h1 == _T_892 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_8997 = 5'h2 == _T_892 ? welem[2] : _GEN_8996; // @[Execute.scala 117:10]
  assign _GEN_8998 = 5'h3 == _T_892 ? welem[3] : _GEN_8997; // @[Execute.scala 117:10]
  assign _GEN_8999 = 5'h4 == _T_892 ? welem[4] : _GEN_8998; // @[Execute.scala 117:10]
  assign _GEN_9000 = 5'h5 == _T_892 ? welem[5] : _GEN_8999; // @[Execute.scala 117:10]
  assign _GEN_9001 = 5'h6 == _T_892 ? welem[6] : _GEN_9000; // @[Execute.scala 117:10]
  assign _GEN_9002 = 5'h7 == _T_892 ? welem[7] : _GEN_9001; // @[Execute.scala 117:10]
  assign _GEN_9003 = 5'h8 == _T_892 ? welem[8] : _GEN_9002; // @[Execute.scala 117:10]
  assign _GEN_9004 = 5'h9 == _T_892 ? welem[9] : _GEN_9003; // @[Execute.scala 117:10]
  assign _GEN_9005 = 5'ha == _T_892 ? welem[10] : _GEN_9004; // @[Execute.scala 117:10]
  assign _GEN_9006 = 5'hb == _T_892 ? welem[11] : _GEN_9005; // @[Execute.scala 117:10]
  assign _GEN_9007 = 5'hc == _T_892 ? welem[12] : _GEN_9006; // @[Execute.scala 117:10]
  assign _GEN_9008 = 5'hd == _T_892 ? welem[13] : _GEN_9007; // @[Execute.scala 117:10]
  assign _GEN_9009 = 5'he == _T_892 ? welem[14] : _GEN_9008; // @[Execute.scala 117:10]
  assign _GEN_9010 = 5'hf == _T_892 ? welem[15] : _GEN_9009; // @[Execute.scala 117:10]
  assign _GEN_9011 = 5'h10 == _T_892 ? welem[16] : _GEN_9010; // @[Execute.scala 117:10]
  assign _GEN_9012 = 5'h11 == _T_892 ? welem[17] : _GEN_9011; // @[Execute.scala 117:10]
  assign _GEN_9013 = 5'h12 == _T_892 ? welem[18] : _GEN_9012; // @[Execute.scala 117:10]
  assign _GEN_9014 = 5'h13 == _T_892 ? welem[19] : _GEN_9013; // @[Execute.scala 117:10]
  assign _GEN_9015 = 5'h14 == _T_892 ? welem[20] : _GEN_9014; // @[Execute.scala 117:10]
  assign _GEN_9016 = 5'h15 == _T_892 ? welem[21] : _GEN_9015; // @[Execute.scala 117:10]
  assign _GEN_9017 = 5'h16 == _T_892 ? welem[22] : _GEN_9016; // @[Execute.scala 117:10]
  assign _GEN_9018 = 5'h17 == _T_892 ? welem[23] : _GEN_9017; // @[Execute.scala 117:10]
  assign _GEN_9019 = 5'h18 == _T_892 ? welem[24] : _GEN_9018; // @[Execute.scala 117:10]
  assign _GEN_9020 = 5'h19 == _T_892 ? welem[25] : _GEN_9019; // @[Execute.scala 117:10]
  assign _GEN_9021 = 5'h1a == _T_892 ? welem[26] : _GEN_9020; // @[Execute.scala 117:10]
  assign _GEN_9022 = 5'h1b == _T_892 ? welem[27] : _GEN_9021; // @[Execute.scala 117:10]
  assign _GEN_9023 = 5'h1c == _T_892 ? welem[28] : _GEN_9022; // @[Execute.scala 117:10]
  assign _GEN_9024 = 5'h1d == _T_892 ? welem[29] : _GEN_9023; // @[Execute.scala 117:10]
  assign _GEN_9025 = 5'h1e == _T_892 ? welem[30] : _GEN_9024; // @[Execute.scala 117:10]
  assign _GEN_9026 = 5'h1f == _T_892 ? welem[31] : _GEN_9025; // @[Execute.scala 117:10]
  assign _T_893 = _T_888 ? _GEN_8994 : _GEN_9026; // @[Execute.scala 117:10]
  assign _T_894 = r[4:0] < 5'h16; // @[Execute.scala 117:15]
  assign _T_896 = r[4:0] - 5'h16; // @[Execute.scala 117:37]
  assign _T_898 = 5'ha + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9028 = 5'h1 == _T_896 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9029 = 5'h2 == _T_896 ? welem[2] : _GEN_9028; // @[Execute.scala 117:10]
  assign _GEN_9030 = 5'h3 == _T_896 ? welem[3] : _GEN_9029; // @[Execute.scala 117:10]
  assign _GEN_9031 = 5'h4 == _T_896 ? welem[4] : _GEN_9030; // @[Execute.scala 117:10]
  assign _GEN_9032 = 5'h5 == _T_896 ? welem[5] : _GEN_9031; // @[Execute.scala 117:10]
  assign _GEN_9033 = 5'h6 == _T_896 ? welem[6] : _GEN_9032; // @[Execute.scala 117:10]
  assign _GEN_9034 = 5'h7 == _T_896 ? welem[7] : _GEN_9033; // @[Execute.scala 117:10]
  assign _GEN_9035 = 5'h8 == _T_896 ? welem[8] : _GEN_9034; // @[Execute.scala 117:10]
  assign _GEN_9036 = 5'h9 == _T_896 ? welem[9] : _GEN_9035; // @[Execute.scala 117:10]
  assign _GEN_9037 = 5'ha == _T_896 ? welem[10] : _GEN_9036; // @[Execute.scala 117:10]
  assign _GEN_9038 = 5'hb == _T_896 ? welem[11] : _GEN_9037; // @[Execute.scala 117:10]
  assign _GEN_9039 = 5'hc == _T_896 ? welem[12] : _GEN_9038; // @[Execute.scala 117:10]
  assign _GEN_9040 = 5'hd == _T_896 ? welem[13] : _GEN_9039; // @[Execute.scala 117:10]
  assign _GEN_9041 = 5'he == _T_896 ? welem[14] : _GEN_9040; // @[Execute.scala 117:10]
  assign _GEN_9042 = 5'hf == _T_896 ? welem[15] : _GEN_9041; // @[Execute.scala 117:10]
  assign _GEN_9043 = 5'h10 == _T_896 ? welem[16] : _GEN_9042; // @[Execute.scala 117:10]
  assign _GEN_9044 = 5'h11 == _T_896 ? welem[17] : _GEN_9043; // @[Execute.scala 117:10]
  assign _GEN_9045 = 5'h12 == _T_896 ? welem[18] : _GEN_9044; // @[Execute.scala 117:10]
  assign _GEN_9046 = 5'h13 == _T_896 ? welem[19] : _GEN_9045; // @[Execute.scala 117:10]
  assign _GEN_9047 = 5'h14 == _T_896 ? welem[20] : _GEN_9046; // @[Execute.scala 117:10]
  assign _GEN_9048 = 5'h15 == _T_896 ? welem[21] : _GEN_9047; // @[Execute.scala 117:10]
  assign _GEN_9049 = 5'h16 == _T_896 ? welem[22] : _GEN_9048; // @[Execute.scala 117:10]
  assign _GEN_9050 = 5'h17 == _T_896 ? welem[23] : _GEN_9049; // @[Execute.scala 117:10]
  assign _GEN_9051 = 5'h18 == _T_896 ? welem[24] : _GEN_9050; // @[Execute.scala 117:10]
  assign _GEN_9052 = 5'h19 == _T_896 ? welem[25] : _GEN_9051; // @[Execute.scala 117:10]
  assign _GEN_9053 = 5'h1a == _T_896 ? welem[26] : _GEN_9052; // @[Execute.scala 117:10]
  assign _GEN_9054 = 5'h1b == _T_896 ? welem[27] : _GEN_9053; // @[Execute.scala 117:10]
  assign _GEN_9055 = 5'h1c == _T_896 ? welem[28] : _GEN_9054; // @[Execute.scala 117:10]
  assign _GEN_9056 = 5'h1d == _T_896 ? welem[29] : _GEN_9055; // @[Execute.scala 117:10]
  assign _GEN_9057 = 5'h1e == _T_896 ? welem[30] : _GEN_9056; // @[Execute.scala 117:10]
  assign _GEN_9058 = 5'h1f == _T_896 ? welem[31] : _GEN_9057; // @[Execute.scala 117:10]
  assign _GEN_9060 = 5'h1 == _T_898 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9061 = 5'h2 == _T_898 ? welem[2] : _GEN_9060; // @[Execute.scala 117:10]
  assign _GEN_9062 = 5'h3 == _T_898 ? welem[3] : _GEN_9061; // @[Execute.scala 117:10]
  assign _GEN_9063 = 5'h4 == _T_898 ? welem[4] : _GEN_9062; // @[Execute.scala 117:10]
  assign _GEN_9064 = 5'h5 == _T_898 ? welem[5] : _GEN_9063; // @[Execute.scala 117:10]
  assign _GEN_9065 = 5'h6 == _T_898 ? welem[6] : _GEN_9064; // @[Execute.scala 117:10]
  assign _GEN_9066 = 5'h7 == _T_898 ? welem[7] : _GEN_9065; // @[Execute.scala 117:10]
  assign _GEN_9067 = 5'h8 == _T_898 ? welem[8] : _GEN_9066; // @[Execute.scala 117:10]
  assign _GEN_9068 = 5'h9 == _T_898 ? welem[9] : _GEN_9067; // @[Execute.scala 117:10]
  assign _GEN_9069 = 5'ha == _T_898 ? welem[10] : _GEN_9068; // @[Execute.scala 117:10]
  assign _GEN_9070 = 5'hb == _T_898 ? welem[11] : _GEN_9069; // @[Execute.scala 117:10]
  assign _GEN_9071 = 5'hc == _T_898 ? welem[12] : _GEN_9070; // @[Execute.scala 117:10]
  assign _GEN_9072 = 5'hd == _T_898 ? welem[13] : _GEN_9071; // @[Execute.scala 117:10]
  assign _GEN_9073 = 5'he == _T_898 ? welem[14] : _GEN_9072; // @[Execute.scala 117:10]
  assign _GEN_9074 = 5'hf == _T_898 ? welem[15] : _GEN_9073; // @[Execute.scala 117:10]
  assign _GEN_9075 = 5'h10 == _T_898 ? welem[16] : _GEN_9074; // @[Execute.scala 117:10]
  assign _GEN_9076 = 5'h11 == _T_898 ? welem[17] : _GEN_9075; // @[Execute.scala 117:10]
  assign _GEN_9077 = 5'h12 == _T_898 ? welem[18] : _GEN_9076; // @[Execute.scala 117:10]
  assign _GEN_9078 = 5'h13 == _T_898 ? welem[19] : _GEN_9077; // @[Execute.scala 117:10]
  assign _GEN_9079 = 5'h14 == _T_898 ? welem[20] : _GEN_9078; // @[Execute.scala 117:10]
  assign _GEN_9080 = 5'h15 == _T_898 ? welem[21] : _GEN_9079; // @[Execute.scala 117:10]
  assign _GEN_9081 = 5'h16 == _T_898 ? welem[22] : _GEN_9080; // @[Execute.scala 117:10]
  assign _GEN_9082 = 5'h17 == _T_898 ? welem[23] : _GEN_9081; // @[Execute.scala 117:10]
  assign _GEN_9083 = 5'h18 == _T_898 ? welem[24] : _GEN_9082; // @[Execute.scala 117:10]
  assign _GEN_9084 = 5'h19 == _T_898 ? welem[25] : _GEN_9083; // @[Execute.scala 117:10]
  assign _GEN_9085 = 5'h1a == _T_898 ? welem[26] : _GEN_9084; // @[Execute.scala 117:10]
  assign _GEN_9086 = 5'h1b == _T_898 ? welem[27] : _GEN_9085; // @[Execute.scala 117:10]
  assign _GEN_9087 = 5'h1c == _T_898 ? welem[28] : _GEN_9086; // @[Execute.scala 117:10]
  assign _GEN_9088 = 5'h1d == _T_898 ? welem[29] : _GEN_9087; // @[Execute.scala 117:10]
  assign _GEN_9089 = 5'h1e == _T_898 ? welem[30] : _GEN_9088; // @[Execute.scala 117:10]
  assign _GEN_9090 = 5'h1f == _T_898 ? welem[31] : _GEN_9089; // @[Execute.scala 117:10]
  assign _T_899 = _T_894 ? _GEN_9058 : _GEN_9090; // @[Execute.scala 117:10]
  assign _T_900 = r[4:0] < 5'h15; // @[Execute.scala 117:15]
  assign _T_902 = r[4:0] - 5'h15; // @[Execute.scala 117:37]
  assign _T_904 = 5'hb + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9092 = 5'h1 == _T_902 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9093 = 5'h2 == _T_902 ? welem[2] : _GEN_9092; // @[Execute.scala 117:10]
  assign _GEN_9094 = 5'h3 == _T_902 ? welem[3] : _GEN_9093; // @[Execute.scala 117:10]
  assign _GEN_9095 = 5'h4 == _T_902 ? welem[4] : _GEN_9094; // @[Execute.scala 117:10]
  assign _GEN_9096 = 5'h5 == _T_902 ? welem[5] : _GEN_9095; // @[Execute.scala 117:10]
  assign _GEN_9097 = 5'h6 == _T_902 ? welem[6] : _GEN_9096; // @[Execute.scala 117:10]
  assign _GEN_9098 = 5'h7 == _T_902 ? welem[7] : _GEN_9097; // @[Execute.scala 117:10]
  assign _GEN_9099 = 5'h8 == _T_902 ? welem[8] : _GEN_9098; // @[Execute.scala 117:10]
  assign _GEN_9100 = 5'h9 == _T_902 ? welem[9] : _GEN_9099; // @[Execute.scala 117:10]
  assign _GEN_9101 = 5'ha == _T_902 ? welem[10] : _GEN_9100; // @[Execute.scala 117:10]
  assign _GEN_9102 = 5'hb == _T_902 ? welem[11] : _GEN_9101; // @[Execute.scala 117:10]
  assign _GEN_9103 = 5'hc == _T_902 ? welem[12] : _GEN_9102; // @[Execute.scala 117:10]
  assign _GEN_9104 = 5'hd == _T_902 ? welem[13] : _GEN_9103; // @[Execute.scala 117:10]
  assign _GEN_9105 = 5'he == _T_902 ? welem[14] : _GEN_9104; // @[Execute.scala 117:10]
  assign _GEN_9106 = 5'hf == _T_902 ? welem[15] : _GEN_9105; // @[Execute.scala 117:10]
  assign _GEN_9107 = 5'h10 == _T_902 ? welem[16] : _GEN_9106; // @[Execute.scala 117:10]
  assign _GEN_9108 = 5'h11 == _T_902 ? welem[17] : _GEN_9107; // @[Execute.scala 117:10]
  assign _GEN_9109 = 5'h12 == _T_902 ? welem[18] : _GEN_9108; // @[Execute.scala 117:10]
  assign _GEN_9110 = 5'h13 == _T_902 ? welem[19] : _GEN_9109; // @[Execute.scala 117:10]
  assign _GEN_9111 = 5'h14 == _T_902 ? welem[20] : _GEN_9110; // @[Execute.scala 117:10]
  assign _GEN_9112 = 5'h15 == _T_902 ? welem[21] : _GEN_9111; // @[Execute.scala 117:10]
  assign _GEN_9113 = 5'h16 == _T_902 ? welem[22] : _GEN_9112; // @[Execute.scala 117:10]
  assign _GEN_9114 = 5'h17 == _T_902 ? welem[23] : _GEN_9113; // @[Execute.scala 117:10]
  assign _GEN_9115 = 5'h18 == _T_902 ? welem[24] : _GEN_9114; // @[Execute.scala 117:10]
  assign _GEN_9116 = 5'h19 == _T_902 ? welem[25] : _GEN_9115; // @[Execute.scala 117:10]
  assign _GEN_9117 = 5'h1a == _T_902 ? welem[26] : _GEN_9116; // @[Execute.scala 117:10]
  assign _GEN_9118 = 5'h1b == _T_902 ? welem[27] : _GEN_9117; // @[Execute.scala 117:10]
  assign _GEN_9119 = 5'h1c == _T_902 ? welem[28] : _GEN_9118; // @[Execute.scala 117:10]
  assign _GEN_9120 = 5'h1d == _T_902 ? welem[29] : _GEN_9119; // @[Execute.scala 117:10]
  assign _GEN_9121 = 5'h1e == _T_902 ? welem[30] : _GEN_9120; // @[Execute.scala 117:10]
  assign _GEN_9122 = 5'h1f == _T_902 ? welem[31] : _GEN_9121; // @[Execute.scala 117:10]
  assign _GEN_9124 = 5'h1 == _T_904 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9125 = 5'h2 == _T_904 ? welem[2] : _GEN_9124; // @[Execute.scala 117:10]
  assign _GEN_9126 = 5'h3 == _T_904 ? welem[3] : _GEN_9125; // @[Execute.scala 117:10]
  assign _GEN_9127 = 5'h4 == _T_904 ? welem[4] : _GEN_9126; // @[Execute.scala 117:10]
  assign _GEN_9128 = 5'h5 == _T_904 ? welem[5] : _GEN_9127; // @[Execute.scala 117:10]
  assign _GEN_9129 = 5'h6 == _T_904 ? welem[6] : _GEN_9128; // @[Execute.scala 117:10]
  assign _GEN_9130 = 5'h7 == _T_904 ? welem[7] : _GEN_9129; // @[Execute.scala 117:10]
  assign _GEN_9131 = 5'h8 == _T_904 ? welem[8] : _GEN_9130; // @[Execute.scala 117:10]
  assign _GEN_9132 = 5'h9 == _T_904 ? welem[9] : _GEN_9131; // @[Execute.scala 117:10]
  assign _GEN_9133 = 5'ha == _T_904 ? welem[10] : _GEN_9132; // @[Execute.scala 117:10]
  assign _GEN_9134 = 5'hb == _T_904 ? welem[11] : _GEN_9133; // @[Execute.scala 117:10]
  assign _GEN_9135 = 5'hc == _T_904 ? welem[12] : _GEN_9134; // @[Execute.scala 117:10]
  assign _GEN_9136 = 5'hd == _T_904 ? welem[13] : _GEN_9135; // @[Execute.scala 117:10]
  assign _GEN_9137 = 5'he == _T_904 ? welem[14] : _GEN_9136; // @[Execute.scala 117:10]
  assign _GEN_9138 = 5'hf == _T_904 ? welem[15] : _GEN_9137; // @[Execute.scala 117:10]
  assign _GEN_9139 = 5'h10 == _T_904 ? welem[16] : _GEN_9138; // @[Execute.scala 117:10]
  assign _GEN_9140 = 5'h11 == _T_904 ? welem[17] : _GEN_9139; // @[Execute.scala 117:10]
  assign _GEN_9141 = 5'h12 == _T_904 ? welem[18] : _GEN_9140; // @[Execute.scala 117:10]
  assign _GEN_9142 = 5'h13 == _T_904 ? welem[19] : _GEN_9141; // @[Execute.scala 117:10]
  assign _GEN_9143 = 5'h14 == _T_904 ? welem[20] : _GEN_9142; // @[Execute.scala 117:10]
  assign _GEN_9144 = 5'h15 == _T_904 ? welem[21] : _GEN_9143; // @[Execute.scala 117:10]
  assign _GEN_9145 = 5'h16 == _T_904 ? welem[22] : _GEN_9144; // @[Execute.scala 117:10]
  assign _GEN_9146 = 5'h17 == _T_904 ? welem[23] : _GEN_9145; // @[Execute.scala 117:10]
  assign _GEN_9147 = 5'h18 == _T_904 ? welem[24] : _GEN_9146; // @[Execute.scala 117:10]
  assign _GEN_9148 = 5'h19 == _T_904 ? welem[25] : _GEN_9147; // @[Execute.scala 117:10]
  assign _GEN_9149 = 5'h1a == _T_904 ? welem[26] : _GEN_9148; // @[Execute.scala 117:10]
  assign _GEN_9150 = 5'h1b == _T_904 ? welem[27] : _GEN_9149; // @[Execute.scala 117:10]
  assign _GEN_9151 = 5'h1c == _T_904 ? welem[28] : _GEN_9150; // @[Execute.scala 117:10]
  assign _GEN_9152 = 5'h1d == _T_904 ? welem[29] : _GEN_9151; // @[Execute.scala 117:10]
  assign _GEN_9153 = 5'h1e == _T_904 ? welem[30] : _GEN_9152; // @[Execute.scala 117:10]
  assign _GEN_9154 = 5'h1f == _T_904 ? welem[31] : _GEN_9153; // @[Execute.scala 117:10]
  assign _T_905 = _T_900 ? _GEN_9122 : _GEN_9154; // @[Execute.scala 117:10]
  assign _T_906 = r[4:0] < 5'h14; // @[Execute.scala 117:15]
  assign _T_908 = r[4:0] - 5'h14; // @[Execute.scala 117:37]
  assign _T_910 = 5'hc + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9156 = 5'h1 == _T_908 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9157 = 5'h2 == _T_908 ? welem[2] : _GEN_9156; // @[Execute.scala 117:10]
  assign _GEN_9158 = 5'h3 == _T_908 ? welem[3] : _GEN_9157; // @[Execute.scala 117:10]
  assign _GEN_9159 = 5'h4 == _T_908 ? welem[4] : _GEN_9158; // @[Execute.scala 117:10]
  assign _GEN_9160 = 5'h5 == _T_908 ? welem[5] : _GEN_9159; // @[Execute.scala 117:10]
  assign _GEN_9161 = 5'h6 == _T_908 ? welem[6] : _GEN_9160; // @[Execute.scala 117:10]
  assign _GEN_9162 = 5'h7 == _T_908 ? welem[7] : _GEN_9161; // @[Execute.scala 117:10]
  assign _GEN_9163 = 5'h8 == _T_908 ? welem[8] : _GEN_9162; // @[Execute.scala 117:10]
  assign _GEN_9164 = 5'h9 == _T_908 ? welem[9] : _GEN_9163; // @[Execute.scala 117:10]
  assign _GEN_9165 = 5'ha == _T_908 ? welem[10] : _GEN_9164; // @[Execute.scala 117:10]
  assign _GEN_9166 = 5'hb == _T_908 ? welem[11] : _GEN_9165; // @[Execute.scala 117:10]
  assign _GEN_9167 = 5'hc == _T_908 ? welem[12] : _GEN_9166; // @[Execute.scala 117:10]
  assign _GEN_9168 = 5'hd == _T_908 ? welem[13] : _GEN_9167; // @[Execute.scala 117:10]
  assign _GEN_9169 = 5'he == _T_908 ? welem[14] : _GEN_9168; // @[Execute.scala 117:10]
  assign _GEN_9170 = 5'hf == _T_908 ? welem[15] : _GEN_9169; // @[Execute.scala 117:10]
  assign _GEN_9171 = 5'h10 == _T_908 ? welem[16] : _GEN_9170; // @[Execute.scala 117:10]
  assign _GEN_9172 = 5'h11 == _T_908 ? welem[17] : _GEN_9171; // @[Execute.scala 117:10]
  assign _GEN_9173 = 5'h12 == _T_908 ? welem[18] : _GEN_9172; // @[Execute.scala 117:10]
  assign _GEN_9174 = 5'h13 == _T_908 ? welem[19] : _GEN_9173; // @[Execute.scala 117:10]
  assign _GEN_9175 = 5'h14 == _T_908 ? welem[20] : _GEN_9174; // @[Execute.scala 117:10]
  assign _GEN_9176 = 5'h15 == _T_908 ? welem[21] : _GEN_9175; // @[Execute.scala 117:10]
  assign _GEN_9177 = 5'h16 == _T_908 ? welem[22] : _GEN_9176; // @[Execute.scala 117:10]
  assign _GEN_9178 = 5'h17 == _T_908 ? welem[23] : _GEN_9177; // @[Execute.scala 117:10]
  assign _GEN_9179 = 5'h18 == _T_908 ? welem[24] : _GEN_9178; // @[Execute.scala 117:10]
  assign _GEN_9180 = 5'h19 == _T_908 ? welem[25] : _GEN_9179; // @[Execute.scala 117:10]
  assign _GEN_9181 = 5'h1a == _T_908 ? welem[26] : _GEN_9180; // @[Execute.scala 117:10]
  assign _GEN_9182 = 5'h1b == _T_908 ? welem[27] : _GEN_9181; // @[Execute.scala 117:10]
  assign _GEN_9183 = 5'h1c == _T_908 ? welem[28] : _GEN_9182; // @[Execute.scala 117:10]
  assign _GEN_9184 = 5'h1d == _T_908 ? welem[29] : _GEN_9183; // @[Execute.scala 117:10]
  assign _GEN_9185 = 5'h1e == _T_908 ? welem[30] : _GEN_9184; // @[Execute.scala 117:10]
  assign _GEN_9186 = 5'h1f == _T_908 ? welem[31] : _GEN_9185; // @[Execute.scala 117:10]
  assign _GEN_9188 = 5'h1 == _T_910 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9189 = 5'h2 == _T_910 ? welem[2] : _GEN_9188; // @[Execute.scala 117:10]
  assign _GEN_9190 = 5'h3 == _T_910 ? welem[3] : _GEN_9189; // @[Execute.scala 117:10]
  assign _GEN_9191 = 5'h4 == _T_910 ? welem[4] : _GEN_9190; // @[Execute.scala 117:10]
  assign _GEN_9192 = 5'h5 == _T_910 ? welem[5] : _GEN_9191; // @[Execute.scala 117:10]
  assign _GEN_9193 = 5'h6 == _T_910 ? welem[6] : _GEN_9192; // @[Execute.scala 117:10]
  assign _GEN_9194 = 5'h7 == _T_910 ? welem[7] : _GEN_9193; // @[Execute.scala 117:10]
  assign _GEN_9195 = 5'h8 == _T_910 ? welem[8] : _GEN_9194; // @[Execute.scala 117:10]
  assign _GEN_9196 = 5'h9 == _T_910 ? welem[9] : _GEN_9195; // @[Execute.scala 117:10]
  assign _GEN_9197 = 5'ha == _T_910 ? welem[10] : _GEN_9196; // @[Execute.scala 117:10]
  assign _GEN_9198 = 5'hb == _T_910 ? welem[11] : _GEN_9197; // @[Execute.scala 117:10]
  assign _GEN_9199 = 5'hc == _T_910 ? welem[12] : _GEN_9198; // @[Execute.scala 117:10]
  assign _GEN_9200 = 5'hd == _T_910 ? welem[13] : _GEN_9199; // @[Execute.scala 117:10]
  assign _GEN_9201 = 5'he == _T_910 ? welem[14] : _GEN_9200; // @[Execute.scala 117:10]
  assign _GEN_9202 = 5'hf == _T_910 ? welem[15] : _GEN_9201; // @[Execute.scala 117:10]
  assign _GEN_9203 = 5'h10 == _T_910 ? welem[16] : _GEN_9202; // @[Execute.scala 117:10]
  assign _GEN_9204 = 5'h11 == _T_910 ? welem[17] : _GEN_9203; // @[Execute.scala 117:10]
  assign _GEN_9205 = 5'h12 == _T_910 ? welem[18] : _GEN_9204; // @[Execute.scala 117:10]
  assign _GEN_9206 = 5'h13 == _T_910 ? welem[19] : _GEN_9205; // @[Execute.scala 117:10]
  assign _GEN_9207 = 5'h14 == _T_910 ? welem[20] : _GEN_9206; // @[Execute.scala 117:10]
  assign _GEN_9208 = 5'h15 == _T_910 ? welem[21] : _GEN_9207; // @[Execute.scala 117:10]
  assign _GEN_9209 = 5'h16 == _T_910 ? welem[22] : _GEN_9208; // @[Execute.scala 117:10]
  assign _GEN_9210 = 5'h17 == _T_910 ? welem[23] : _GEN_9209; // @[Execute.scala 117:10]
  assign _GEN_9211 = 5'h18 == _T_910 ? welem[24] : _GEN_9210; // @[Execute.scala 117:10]
  assign _GEN_9212 = 5'h19 == _T_910 ? welem[25] : _GEN_9211; // @[Execute.scala 117:10]
  assign _GEN_9213 = 5'h1a == _T_910 ? welem[26] : _GEN_9212; // @[Execute.scala 117:10]
  assign _GEN_9214 = 5'h1b == _T_910 ? welem[27] : _GEN_9213; // @[Execute.scala 117:10]
  assign _GEN_9215 = 5'h1c == _T_910 ? welem[28] : _GEN_9214; // @[Execute.scala 117:10]
  assign _GEN_9216 = 5'h1d == _T_910 ? welem[29] : _GEN_9215; // @[Execute.scala 117:10]
  assign _GEN_9217 = 5'h1e == _T_910 ? welem[30] : _GEN_9216; // @[Execute.scala 117:10]
  assign _GEN_9218 = 5'h1f == _T_910 ? welem[31] : _GEN_9217; // @[Execute.scala 117:10]
  assign _T_911 = _T_906 ? _GEN_9186 : _GEN_9218; // @[Execute.scala 117:10]
  assign _T_912 = r[4:0] < 5'h13; // @[Execute.scala 117:15]
  assign _T_914 = r[4:0] - 5'h13; // @[Execute.scala 117:37]
  assign _T_916 = 5'hd + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9220 = 5'h1 == _T_914 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9221 = 5'h2 == _T_914 ? welem[2] : _GEN_9220; // @[Execute.scala 117:10]
  assign _GEN_9222 = 5'h3 == _T_914 ? welem[3] : _GEN_9221; // @[Execute.scala 117:10]
  assign _GEN_9223 = 5'h4 == _T_914 ? welem[4] : _GEN_9222; // @[Execute.scala 117:10]
  assign _GEN_9224 = 5'h5 == _T_914 ? welem[5] : _GEN_9223; // @[Execute.scala 117:10]
  assign _GEN_9225 = 5'h6 == _T_914 ? welem[6] : _GEN_9224; // @[Execute.scala 117:10]
  assign _GEN_9226 = 5'h7 == _T_914 ? welem[7] : _GEN_9225; // @[Execute.scala 117:10]
  assign _GEN_9227 = 5'h8 == _T_914 ? welem[8] : _GEN_9226; // @[Execute.scala 117:10]
  assign _GEN_9228 = 5'h9 == _T_914 ? welem[9] : _GEN_9227; // @[Execute.scala 117:10]
  assign _GEN_9229 = 5'ha == _T_914 ? welem[10] : _GEN_9228; // @[Execute.scala 117:10]
  assign _GEN_9230 = 5'hb == _T_914 ? welem[11] : _GEN_9229; // @[Execute.scala 117:10]
  assign _GEN_9231 = 5'hc == _T_914 ? welem[12] : _GEN_9230; // @[Execute.scala 117:10]
  assign _GEN_9232 = 5'hd == _T_914 ? welem[13] : _GEN_9231; // @[Execute.scala 117:10]
  assign _GEN_9233 = 5'he == _T_914 ? welem[14] : _GEN_9232; // @[Execute.scala 117:10]
  assign _GEN_9234 = 5'hf == _T_914 ? welem[15] : _GEN_9233; // @[Execute.scala 117:10]
  assign _GEN_9235 = 5'h10 == _T_914 ? welem[16] : _GEN_9234; // @[Execute.scala 117:10]
  assign _GEN_9236 = 5'h11 == _T_914 ? welem[17] : _GEN_9235; // @[Execute.scala 117:10]
  assign _GEN_9237 = 5'h12 == _T_914 ? welem[18] : _GEN_9236; // @[Execute.scala 117:10]
  assign _GEN_9238 = 5'h13 == _T_914 ? welem[19] : _GEN_9237; // @[Execute.scala 117:10]
  assign _GEN_9239 = 5'h14 == _T_914 ? welem[20] : _GEN_9238; // @[Execute.scala 117:10]
  assign _GEN_9240 = 5'h15 == _T_914 ? welem[21] : _GEN_9239; // @[Execute.scala 117:10]
  assign _GEN_9241 = 5'h16 == _T_914 ? welem[22] : _GEN_9240; // @[Execute.scala 117:10]
  assign _GEN_9242 = 5'h17 == _T_914 ? welem[23] : _GEN_9241; // @[Execute.scala 117:10]
  assign _GEN_9243 = 5'h18 == _T_914 ? welem[24] : _GEN_9242; // @[Execute.scala 117:10]
  assign _GEN_9244 = 5'h19 == _T_914 ? welem[25] : _GEN_9243; // @[Execute.scala 117:10]
  assign _GEN_9245 = 5'h1a == _T_914 ? welem[26] : _GEN_9244; // @[Execute.scala 117:10]
  assign _GEN_9246 = 5'h1b == _T_914 ? welem[27] : _GEN_9245; // @[Execute.scala 117:10]
  assign _GEN_9247 = 5'h1c == _T_914 ? welem[28] : _GEN_9246; // @[Execute.scala 117:10]
  assign _GEN_9248 = 5'h1d == _T_914 ? welem[29] : _GEN_9247; // @[Execute.scala 117:10]
  assign _GEN_9249 = 5'h1e == _T_914 ? welem[30] : _GEN_9248; // @[Execute.scala 117:10]
  assign _GEN_9250 = 5'h1f == _T_914 ? welem[31] : _GEN_9249; // @[Execute.scala 117:10]
  assign _GEN_9252 = 5'h1 == _T_916 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9253 = 5'h2 == _T_916 ? welem[2] : _GEN_9252; // @[Execute.scala 117:10]
  assign _GEN_9254 = 5'h3 == _T_916 ? welem[3] : _GEN_9253; // @[Execute.scala 117:10]
  assign _GEN_9255 = 5'h4 == _T_916 ? welem[4] : _GEN_9254; // @[Execute.scala 117:10]
  assign _GEN_9256 = 5'h5 == _T_916 ? welem[5] : _GEN_9255; // @[Execute.scala 117:10]
  assign _GEN_9257 = 5'h6 == _T_916 ? welem[6] : _GEN_9256; // @[Execute.scala 117:10]
  assign _GEN_9258 = 5'h7 == _T_916 ? welem[7] : _GEN_9257; // @[Execute.scala 117:10]
  assign _GEN_9259 = 5'h8 == _T_916 ? welem[8] : _GEN_9258; // @[Execute.scala 117:10]
  assign _GEN_9260 = 5'h9 == _T_916 ? welem[9] : _GEN_9259; // @[Execute.scala 117:10]
  assign _GEN_9261 = 5'ha == _T_916 ? welem[10] : _GEN_9260; // @[Execute.scala 117:10]
  assign _GEN_9262 = 5'hb == _T_916 ? welem[11] : _GEN_9261; // @[Execute.scala 117:10]
  assign _GEN_9263 = 5'hc == _T_916 ? welem[12] : _GEN_9262; // @[Execute.scala 117:10]
  assign _GEN_9264 = 5'hd == _T_916 ? welem[13] : _GEN_9263; // @[Execute.scala 117:10]
  assign _GEN_9265 = 5'he == _T_916 ? welem[14] : _GEN_9264; // @[Execute.scala 117:10]
  assign _GEN_9266 = 5'hf == _T_916 ? welem[15] : _GEN_9265; // @[Execute.scala 117:10]
  assign _GEN_9267 = 5'h10 == _T_916 ? welem[16] : _GEN_9266; // @[Execute.scala 117:10]
  assign _GEN_9268 = 5'h11 == _T_916 ? welem[17] : _GEN_9267; // @[Execute.scala 117:10]
  assign _GEN_9269 = 5'h12 == _T_916 ? welem[18] : _GEN_9268; // @[Execute.scala 117:10]
  assign _GEN_9270 = 5'h13 == _T_916 ? welem[19] : _GEN_9269; // @[Execute.scala 117:10]
  assign _GEN_9271 = 5'h14 == _T_916 ? welem[20] : _GEN_9270; // @[Execute.scala 117:10]
  assign _GEN_9272 = 5'h15 == _T_916 ? welem[21] : _GEN_9271; // @[Execute.scala 117:10]
  assign _GEN_9273 = 5'h16 == _T_916 ? welem[22] : _GEN_9272; // @[Execute.scala 117:10]
  assign _GEN_9274 = 5'h17 == _T_916 ? welem[23] : _GEN_9273; // @[Execute.scala 117:10]
  assign _GEN_9275 = 5'h18 == _T_916 ? welem[24] : _GEN_9274; // @[Execute.scala 117:10]
  assign _GEN_9276 = 5'h19 == _T_916 ? welem[25] : _GEN_9275; // @[Execute.scala 117:10]
  assign _GEN_9277 = 5'h1a == _T_916 ? welem[26] : _GEN_9276; // @[Execute.scala 117:10]
  assign _GEN_9278 = 5'h1b == _T_916 ? welem[27] : _GEN_9277; // @[Execute.scala 117:10]
  assign _GEN_9279 = 5'h1c == _T_916 ? welem[28] : _GEN_9278; // @[Execute.scala 117:10]
  assign _GEN_9280 = 5'h1d == _T_916 ? welem[29] : _GEN_9279; // @[Execute.scala 117:10]
  assign _GEN_9281 = 5'h1e == _T_916 ? welem[30] : _GEN_9280; // @[Execute.scala 117:10]
  assign _GEN_9282 = 5'h1f == _T_916 ? welem[31] : _GEN_9281; // @[Execute.scala 117:10]
  assign _T_917 = _T_912 ? _GEN_9250 : _GEN_9282; // @[Execute.scala 117:10]
  assign _T_918 = r[4:0] < 5'h12; // @[Execute.scala 117:15]
  assign _T_920 = r[4:0] - 5'h12; // @[Execute.scala 117:37]
  assign _T_922 = 5'he + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9284 = 5'h1 == _T_920 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9285 = 5'h2 == _T_920 ? welem[2] : _GEN_9284; // @[Execute.scala 117:10]
  assign _GEN_9286 = 5'h3 == _T_920 ? welem[3] : _GEN_9285; // @[Execute.scala 117:10]
  assign _GEN_9287 = 5'h4 == _T_920 ? welem[4] : _GEN_9286; // @[Execute.scala 117:10]
  assign _GEN_9288 = 5'h5 == _T_920 ? welem[5] : _GEN_9287; // @[Execute.scala 117:10]
  assign _GEN_9289 = 5'h6 == _T_920 ? welem[6] : _GEN_9288; // @[Execute.scala 117:10]
  assign _GEN_9290 = 5'h7 == _T_920 ? welem[7] : _GEN_9289; // @[Execute.scala 117:10]
  assign _GEN_9291 = 5'h8 == _T_920 ? welem[8] : _GEN_9290; // @[Execute.scala 117:10]
  assign _GEN_9292 = 5'h9 == _T_920 ? welem[9] : _GEN_9291; // @[Execute.scala 117:10]
  assign _GEN_9293 = 5'ha == _T_920 ? welem[10] : _GEN_9292; // @[Execute.scala 117:10]
  assign _GEN_9294 = 5'hb == _T_920 ? welem[11] : _GEN_9293; // @[Execute.scala 117:10]
  assign _GEN_9295 = 5'hc == _T_920 ? welem[12] : _GEN_9294; // @[Execute.scala 117:10]
  assign _GEN_9296 = 5'hd == _T_920 ? welem[13] : _GEN_9295; // @[Execute.scala 117:10]
  assign _GEN_9297 = 5'he == _T_920 ? welem[14] : _GEN_9296; // @[Execute.scala 117:10]
  assign _GEN_9298 = 5'hf == _T_920 ? welem[15] : _GEN_9297; // @[Execute.scala 117:10]
  assign _GEN_9299 = 5'h10 == _T_920 ? welem[16] : _GEN_9298; // @[Execute.scala 117:10]
  assign _GEN_9300 = 5'h11 == _T_920 ? welem[17] : _GEN_9299; // @[Execute.scala 117:10]
  assign _GEN_9301 = 5'h12 == _T_920 ? welem[18] : _GEN_9300; // @[Execute.scala 117:10]
  assign _GEN_9302 = 5'h13 == _T_920 ? welem[19] : _GEN_9301; // @[Execute.scala 117:10]
  assign _GEN_9303 = 5'h14 == _T_920 ? welem[20] : _GEN_9302; // @[Execute.scala 117:10]
  assign _GEN_9304 = 5'h15 == _T_920 ? welem[21] : _GEN_9303; // @[Execute.scala 117:10]
  assign _GEN_9305 = 5'h16 == _T_920 ? welem[22] : _GEN_9304; // @[Execute.scala 117:10]
  assign _GEN_9306 = 5'h17 == _T_920 ? welem[23] : _GEN_9305; // @[Execute.scala 117:10]
  assign _GEN_9307 = 5'h18 == _T_920 ? welem[24] : _GEN_9306; // @[Execute.scala 117:10]
  assign _GEN_9308 = 5'h19 == _T_920 ? welem[25] : _GEN_9307; // @[Execute.scala 117:10]
  assign _GEN_9309 = 5'h1a == _T_920 ? welem[26] : _GEN_9308; // @[Execute.scala 117:10]
  assign _GEN_9310 = 5'h1b == _T_920 ? welem[27] : _GEN_9309; // @[Execute.scala 117:10]
  assign _GEN_9311 = 5'h1c == _T_920 ? welem[28] : _GEN_9310; // @[Execute.scala 117:10]
  assign _GEN_9312 = 5'h1d == _T_920 ? welem[29] : _GEN_9311; // @[Execute.scala 117:10]
  assign _GEN_9313 = 5'h1e == _T_920 ? welem[30] : _GEN_9312; // @[Execute.scala 117:10]
  assign _GEN_9314 = 5'h1f == _T_920 ? welem[31] : _GEN_9313; // @[Execute.scala 117:10]
  assign _GEN_9316 = 5'h1 == _T_922 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9317 = 5'h2 == _T_922 ? welem[2] : _GEN_9316; // @[Execute.scala 117:10]
  assign _GEN_9318 = 5'h3 == _T_922 ? welem[3] : _GEN_9317; // @[Execute.scala 117:10]
  assign _GEN_9319 = 5'h4 == _T_922 ? welem[4] : _GEN_9318; // @[Execute.scala 117:10]
  assign _GEN_9320 = 5'h5 == _T_922 ? welem[5] : _GEN_9319; // @[Execute.scala 117:10]
  assign _GEN_9321 = 5'h6 == _T_922 ? welem[6] : _GEN_9320; // @[Execute.scala 117:10]
  assign _GEN_9322 = 5'h7 == _T_922 ? welem[7] : _GEN_9321; // @[Execute.scala 117:10]
  assign _GEN_9323 = 5'h8 == _T_922 ? welem[8] : _GEN_9322; // @[Execute.scala 117:10]
  assign _GEN_9324 = 5'h9 == _T_922 ? welem[9] : _GEN_9323; // @[Execute.scala 117:10]
  assign _GEN_9325 = 5'ha == _T_922 ? welem[10] : _GEN_9324; // @[Execute.scala 117:10]
  assign _GEN_9326 = 5'hb == _T_922 ? welem[11] : _GEN_9325; // @[Execute.scala 117:10]
  assign _GEN_9327 = 5'hc == _T_922 ? welem[12] : _GEN_9326; // @[Execute.scala 117:10]
  assign _GEN_9328 = 5'hd == _T_922 ? welem[13] : _GEN_9327; // @[Execute.scala 117:10]
  assign _GEN_9329 = 5'he == _T_922 ? welem[14] : _GEN_9328; // @[Execute.scala 117:10]
  assign _GEN_9330 = 5'hf == _T_922 ? welem[15] : _GEN_9329; // @[Execute.scala 117:10]
  assign _GEN_9331 = 5'h10 == _T_922 ? welem[16] : _GEN_9330; // @[Execute.scala 117:10]
  assign _GEN_9332 = 5'h11 == _T_922 ? welem[17] : _GEN_9331; // @[Execute.scala 117:10]
  assign _GEN_9333 = 5'h12 == _T_922 ? welem[18] : _GEN_9332; // @[Execute.scala 117:10]
  assign _GEN_9334 = 5'h13 == _T_922 ? welem[19] : _GEN_9333; // @[Execute.scala 117:10]
  assign _GEN_9335 = 5'h14 == _T_922 ? welem[20] : _GEN_9334; // @[Execute.scala 117:10]
  assign _GEN_9336 = 5'h15 == _T_922 ? welem[21] : _GEN_9335; // @[Execute.scala 117:10]
  assign _GEN_9337 = 5'h16 == _T_922 ? welem[22] : _GEN_9336; // @[Execute.scala 117:10]
  assign _GEN_9338 = 5'h17 == _T_922 ? welem[23] : _GEN_9337; // @[Execute.scala 117:10]
  assign _GEN_9339 = 5'h18 == _T_922 ? welem[24] : _GEN_9338; // @[Execute.scala 117:10]
  assign _GEN_9340 = 5'h19 == _T_922 ? welem[25] : _GEN_9339; // @[Execute.scala 117:10]
  assign _GEN_9341 = 5'h1a == _T_922 ? welem[26] : _GEN_9340; // @[Execute.scala 117:10]
  assign _GEN_9342 = 5'h1b == _T_922 ? welem[27] : _GEN_9341; // @[Execute.scala 117:10]
  assign _GEN_9343 = 5'h1c == _T_922 ? welem[28] : _GEN_9342; // @[Execute.scala 117:10]
  assign _GEN_9344 = 5'h1d == _T_922 ? welem[29] : _GEN_9343; // @[Execute.scala 117:10]
  assign _GEN_9345 = 5'h1e == _T_922 ? welem[30] : _GEN_9344; // @[Execute.scala 117:10]
  assign _GEN_9346 = 5'h1f == _T_922 ? welem[31] : _GEN_9345; // @[Execute.scala 117:10]
  assign _T_923 = _T_918 ? _GEN_9314 : _GEN_9346; // @[Execute.scala 117:10]
  assign _T_924 = r[4:0] < 5'h11; // @[Execute.scala 117:15]
  assign _T_926 = r[4:0] - 5'h11; // @[Execute.scala 117:37]
  assign _T_928 = 5'hf + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9348 = 5'h1 == _T_926 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9349 = 5'h2 == _T_926 ? welem[2] : _GEN_9348; // @[Execute.scala 117:10]
  assign _GEN_9350 = 5'h3 == _T_926 ? welem[3] : _GEN_9349; // @[Execute.scala 117:10]
  assign _GEN_9351 = 5'h4 == _T_926 ? welem[4] : _GEN_9350; // @[Execute.scala 117:10]
  assign _GEN_9352 = 5'h5 == _T_926 ? welem[5] : _GEN_9351; // @[Execute.scala 117:10]
  assign _GEN_9353 = 5'h6 == _T_926 ? welem[6] : _GEN_9352; // @[Execute.scala 117:10]
  assign _GEN_9354 = 5'h7 == _T_926 ? welem[7] : _GEN_9353; // @[Execute.scala 117:10]
  assign _GEN_9355 = 5'h8 == _T_926 ? welem[8] : _GEN_9354; // @[Execute.scala 117:10]
  assign _GEN_9356 = 5'h9 == _T_926 ? welem[9] : _GEN_9355; // @[Execute.scala 117:10]
  assign _GEN_9357 = 5'ha == _T_926 ? welem[10] : _GEN_9356; // @[Execute.scala 117:10]
  assign _GEN_9358 = 5'hb == _T_926 ? welem[11] : _GEN_9357; // @[Execute.scala 117:10]
  assign _GEN_9359 = 5'hc == _T_926 ? welem[12] : _GEN_9358; // @[Execute.scala 117:10]
  assign _GEN_9360 = 5'hd == _T_926 ? welem[13] : _GEN_9359; // @[Execute.scala 117:10]
  assign _GEN_9361 = 5'he == _T_926 ? welem[14] : _GEN_9360; // @[Execute.scala 117:10]
  assign _GEN_9362 = 5'hf == _T_926 ? welem[15] : _GEN_9361; // @[Execute.scala 117:10]
  assign _GEN_9363 = 5'h10 == _T_926 ? welem[16] : _GEN_9362; // @[Execute.scala 117:10]
  assign _GEN_9364 = 5'h11 == _T_926 ? welem[17] : _GEN_9363; // @[Execute.scala 117:10]
  assign _GEN_9365 = 5'h12 == _T_926 ? welem[18] : _GEN_9364; // @[Execute.scala 117:10]
  assign _GEN_9366 = 5'h13 == _T_926 ? welem[19] : _GEN_9365; // @[Execute.scala 117:10]
  assign _GEN_9367 = 5'h14 == _T_926 ? welem[20] : _GEN_9366; // @[Execute.scala 117:10]
  assign _GEN_9368 = 5'h15 == _T_926 ? welem[21] : _GEN_9367; // @[Execute.scala 117:10]
  assign _GEN_9369 = 5'h16 == _T_926 ? welem[22] : _GEN_9368; // @[Execute.scala 117:10]
  assign _GEN_9370 = 5'h17 == _T_926 ? welem[23] : _GEN_9369; // @[Execute.scala 117:10]
  assign _GEN_9371 = 5'h18 == _T_926 ? welem[24] : _GEN_9370; // @[Execute.scala 117:10]
  assign _GEN_9372 = 5'h19 == _T_926 ? welem[25] : _GEN_9371; // @[Execute.scala 117:10]
  assign _GEN_9373 = 5'h1a == _T_926 ? welem[26] : _GEN_9372; // @[Execute.scala 117:10]
  assign _GEN_9374 = 5'h1b == _T_926 ? welem[27] : _GEN_9373; // @[Execute.scala 117:10]
  assign _GEN_9375 = 5'h1c == _T_926 ? welem[28] : _GEN_9374; // @[Execute.scala 117:10]
  assign _GEN_9376 = 5'h1d == _T_926 ? welem[29] : _GEN_9375; // @[Execute.scala 117:10]
  assign _GEN_9377 = 5'h1e == _T_926 ? welem[30] : _GEN_9376; // @[Execute.scala 117:10]
  assign _GEN_9378 = 5'h1f == _T_926 ? welem[31] : _GEN_9377; // @[Execute.scala 117:10]
  assign _GEN_9380 = 5'h1 == _T_928 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9381 = 5'h2 == _T_928 ? welem[2] : _GEN_9380; // @[Execute.scala 117:10]
  assign _GEN_9382 = 5'h3 == _T_928 ? welem[3] : _GEN_9381; // @[Execute.scala 117:10]
  assign _GEN_9383 = 5'h4 == _T_928 ? welem[4] : _GEN_9382; // @[Execute.scala 117:10]
  assign _GEN_9384 = 5'h5 == _T_928 ? welem[5] : _GEN_9383; // @[Execute.scala 117:10]
  assign _GEN_9385 = 5'h6 == _T_928 ? welem[6] : _GEN_9384; // @[Execute.scala 117:10]
  assign _GEN_9386 = 5'h7 == _T_928 ? welem[7] : _GEN_9385; // @[Execute.scala 117:10]
  assign _GEN_9387 = 5'h8 == _T_928 ? welem[8] : _GEN_9386; // @[Execute.scala 117:10]
  assign _GEN_9388 = 5'h9 == _T_928 ? welem[9] : _GEN_9387; // @[Execute.scala 117:10]
  assign _GEN_9389 = 5'ha == _T_928 ? welem[10] : _GEN_9388; // @[Execute.scala 117:10]
  assign _GEN_9390 = 5'hb == _T_928 ? welem[11] : _GEN_9389; // @[Execute.scala 117:10]
  assign _GEN_9391 = 5'hc == _T_928 ? welem[12] : _GEN_9390; // @[Execute.scala 117:10]
  assign _GEN_9392 = 5'hd == _T_928 ? welem[13] : _GEN_9391; // @[Execute.scala 117:10]
  assign _GEN_9393 = 5'he == _T_928 ? welem[14] : _GEN_9392; // @[Execute.scala 117:10]
  assign _GEN_9394 = 5'hf == _T_928 ? welem[15] : _GEN_9393; // @[Execute.scala 117:10]
  assign _GEN_9395 = 5'h10 == _T_928 ? welem[16] : _GEN_9394; // @[Execute.scala 117:10]
  assign _GEN_9396 = 5'h11 == _T_928 ? welem[17] : _GEN_9395; // @[Execute.scala 117:10]
  assign _GEN_9397 = 5'h12 == _T_928 ? welem[18] : _GEN_9396; // @[Execute.scala 117:10]
  assign _GEN_9398 = 5'h13 == _T_928 ? welem[19] : _GEN_9397; // @[Execute.scala 117:10]
  assign _GEN_9399 = 5'h14 == _T_928 ? welem[20] : _GEN_9398; // @[Execute.scala 117:10]
  assign _GEN_9400 = 5'h15 == _T_928 ? welem[21] : _GEN_9399; // @[Execute.scala 117:10]
  assign _GEN_9401 = 5'h16 == _T_928 ? welem[22] : _GEN_9400; // @[Execute.scala 117:10]
  assign _GEN_9402 = 5'h17 == _T_928 ? welem[23] : _GEN_9401; // @[Execute.scala 117:10]
  assign _GEN_9403 = 5'h18 == _T_928 ? welem[24] : _GEN_9402; // @[Execute.scala 117:10]
  assign _GEN_9404 = 5'h19 == _T_928 ? welem[25] : _GEN_9403; // @[Execute.scala 117:10]
  assign _GEN_9405 = 5'h1a == _T_928 ? welem[26] : _GEN_9404; // @[Execute.scala 117:10]
  assign _GEN_9406 = 5'h1b == _T_928 ? welem[27] : _GEN_9405; // @[Execute.scala 117:10]
  assign _GEN_9407 = 5'h1c == _T_928 ? welem[28] : _GEN_9406; // @[Execute.scala 117:10]
  assign _GEN_9408 = 5'h1d == _T_928 ? welem[29] : _GEN_9407; // @[Execute.scala 117:10]
  assign _GEN_9409 = 5'h1e == _T_928 ? welem[30] : _GEN_9408; // @[Execute.scala 117:10]
  assign _GEN_9410 = 5'h1f == _T_928 ? welem[31] : _GEN_9409; // @[Execute.scala 117:10]
  assign _T_929 = _T_924 ? _GEN_9378 : _GEN_9410; // @[Execute.scala 117:10]
  assign _T_930 = r[4:0] < 5'h10; // @[Execute.scala 117:15]
  assign _T_932 = r[4:0] - 5'h10; // @[Execute.scala 117:37]
  assign _T_934 = 5'h10 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9412 = 5'h1 == _T_932 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9413 = 5'h2 == _T_932 ? welem[2] : _GEN_9412; // @[Execute.scala 117:10]
  assign _GEN_9414 = 5'h3 == _T_932 ? welem[3] : _GEN_9413; // @[Execute.scala 117:10]
  assign _GEN_9415 = 5'h4 == _T_932 ? welem[4] : _GEN_9414; // @[Execute.scala 117:10]
  assign _GEN_9416 = 5'h5 == _T_932 ? welem[5] : _GEN_9415; // @[Execute.scala 117:10]
  assign _GEN_9417 = 5'h6 == _T_932 ? welem[6] : _GEN_9416; // @[Execute.scala 117:10]
  assign _GEN_9418 = 5'h7 == _T_932 ? welem[7] : _GEN_9417; // @[Execute.scala 117:10]
  assign _GEN_9419 = 5'h8 == _T_932 ? welem[8] : _GEN_9418; // @[Execute.scala 117:10]
  assign _GEN_9420 = 5'h9 == _T_932 ? welem[9] : _GEN_9419; // @[Execute.scala 117:10]
  assign _GEN_9421 = 5'ha == _T_932 ? welem[10] : _GEN_9420; // @[Execute.scala 117:10]
  assign _GEN_9422 = 5'hb == _T_932 ? welem[11] : _GEN_9421; // @[Execute.scala 117:10]
  assign _GEN_9423 = 5'hc == _T_932 ? welem[12] : _GEN_9422; // @[Execute.scala 117:10]
  assign _GEN_9424 = 5'hd == _T_932 ? welem[13] : _GEN_9423; // @[Execute.scala 117:10]
  assign _GEN_9425 = 5'he == _T_932 ? welem[14] : _GEN_9424; // @[Execute.scala 117:10]
  assign _GEN_9426 = 5'hf == _T_932 ? welem[15] : _GEN_9425; // @[Execute.scala 117:10]
  assign _GEN_9427 = 5'h10 == _T_932 ? welem[16] : _GEN_9426; // @[Execute.scala 117:10]
  assign _GEN_9428 = 5'h11 == _T_932 ? welem[17] : _GEN_9427; // @[Execute.scala 117:10]
  assign _GEN_9429 = 5'h12 == _T_932 ? welem[18] : _GEN_9428; // @[Execute.scala 117:10]
  assign _GEN_9430 = 5'h13 == _T_932 ? welem[19] : _GEN_9429; // @[Execute.scala 117:10]
  assign _GEN_9431 = 5'h14 == _T_932 ? welem[20] : _GEN_9430; // @[Execute.scala 117:10]
  assign _GEN_9432 = 5'h15 == _T_932 ? welem[21] : _GEN_9431; // @[Execute.scala 117:10]
  assign _GEN_9433 = 5'h16 == _T_932 ? welem[22] : _GEN_9432; // @[Execute.scala 117:10]
  assign _GEN_9434 = 5'h17 == _T_932 ? welem[23] : _GEN_9433; // @[Execute.scala 117:10]
  assign _GEN_9435 = 5'h18 == _T_932 ? welem[24] : _GEN_9434; // @[Execute.scala 117:10]
  assign _GEN_9436 = 5'h19 == _T_932 ? welem[25] : _GEN_9435; // @[Execute.scala 117:10]
  assign _GEN_9437 = 5'h1a == _T_932 ? welem[26] : _GEN_9436; // @[Execute.scala 117:10]
  assign _GEN_9438 = 5'h1b == _T_932 ? welem[27] : _GEN_9437; // @[Execute.scala 117:10]
  assign _GEN_9439 = 5'h1c == _T_932 ? welem[28] : _GEN_9438; // @[Execute.scala 117:10]
  assign _GEN_9440 = 5'h1d == _T_932 ? welem[29] : _GEN_9439; // @[Execute.scala 117:10]
  assign _GEN_9441 = 5'h1e == _T_932 ? welem[30] : _GEN_9440; // @[Execute.scala 117:10]
  assign _GEN_9442 = 5'h1f == _T_932 ? welem[31] : _GEN_9441; // @[Execute.scala 117:10]
  assign _GEN_9444 = 5'h1 == _T_934 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9445 = 5'h2 == _T_934 ? welem[2] : _GEN_9444; // @[Execute.scala 117:10]
  assign _GEN_9446 = 5'h3 == _T_934 ? welem[3] : _GEN_9445; // @[Execute.scala 117:10]
  assign _GEN_9447 = 5'h4 == _T_934 ? welem[4] : _GEN_9446; // @[Execute.scala 117:10]
  assign _GEN_9448 = 5'h5 == _T_934 ? welem[5] : _GEN_9447; // @[Execute.scala 117:10]
  assign _GEN_9449 = 5'h6 == _T_934 ? welem[6] : _GEN_9448; // @[Execute.scala 117:10]
  assign _GEN_9450 = 5'h7 == _T_934 ? welem[7] : _GEN_9449; // @[Execute.scala 117:10]
  assign _GEN_9451 = 5'h8 == _T_934 ? welem[8] : _GEN_9450; // @[Execute.scala 117:10]
  assign _GEN_9452 = 5'h9 == _T_934 ? welem[9] : _GEN_9451; // @[Execute.scala 117:10]
  assign _GEN_9453 = 5'ha == _T_934 ? welem[10] : _GEN_9452; // @[Execute.scala 117:10]
  assign _GEN_9454 = 5'hb == _T_934 ? welem[11] : _GEN_9453; // @[Execute.scala 117:10]
  assign _GEN_9455 = 5'hc == _T_934 ? welem[12] : _GEN_9454; // @[Execute.scala 117:10]
  assign _GEN_9456 = 5'hd == _T_934 ? welem[13] : _GEN_9455; // @[Execute.scala 117:10]
  assign _GEN_9457 = 5'he == _T_934 ? welem[14] : _GEN_9456; // @[Execute.scala 117:10]
  assign _GEN_9458 = 5'hf == _T_934 ? welem[15] : _GEN_9457; // @[Execute.scala 117:10]
  assign _GEN_9459 = 5'h10 == _T_934 ? welem[16] : _GEN_9458; // @[Execute.scala 117:10]
  assign _GEN_9460 = 5'h11 == _T_934 ? welem[17] : _GEN_9459; // @[Execute.scala 117:10]
  assign _GEN_9461 = 5'h12 == _T_934 ? welem[18] : _GEN_9460; // @[Execute.scala 117:10]
  assign _GEN_9462 = 5'h13 == _T_934 ? welem[19] : _GEN_9461; // @[Execute.scala 117:10]
  assign _GEN_9463 = 5'h14 == _T_934 ? welem[20] : _GEN_9462; // @[Execute.scala 117:10]
  assign _GEN_9464 = 5'h15 == _T_934 ? welem[21] : _GEN_9463; // @[Execute.scala 117:10]
  assign _GEN_9465 = 5'h16 == _T_934 ? welem[22] : _GEN_9464; // @[Execute.scala 117:10]
  assign _GEN_9466 = 5'h17 == _T_934 ? welem[23] : _GEN_9465; // @[Execute.scala 117:10]
  assign _GEN_9467 = 5'h18 == _T_934 ? welem[24] : _GEN_9466; // @[Execute.scala 117:10]
  assign _GEN_9468 = 5'h19 == _T_934 ? welem[25] : _GEN_9467; // @[Execute.scala 117:10]
  assign _GEN_9469 = 5'h1a == _T_934 ? welem[26] : _GEN_9468; // @[Execute.scala 117:10]
  assign _GEN_9470 = 5'h1b == _T_934 ? welem[27] : _GEN_9469; // @[Execute.scala 117:10]
  assign _GEN_9471 = 5'h1c == _T_934 ? welem[28] : _GEN_9470; // @[Execute.scala 117:10]
  assign _GEN_9472 = 5'h1d == _T_934 ? welem[29] : _GEN_9471; // @[Execute.scala 117:10]
  assign _GEN_9473 = 5'h1e == _T_934 ? welem[30] : _GEN_9472; // @[Execute.scala 117:10]
  assign _GEN_9474 = 5'h1f == _T_934 ? welem[31] : _GEN_9473; // @[Execute.scala 117:10]
  assign _T_935 = _T_930 ? _GEN_9442 : _GEN_9474; // @[Execute.scala 117:10]
  assign _T_936 = r[4:0] < 5'hf; // @[Execute.scala 117:15]
  assign _T_938 = r[4:0] - 5'hf; // @[Execute.scala 117:37]
  assign _T_940 = 5'h11 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9476 = 5'h1 == _T_938 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9477 = 5'h2 == _T_938 ? welem[2] : _GEN_9476; // @[Execute.scala 117:10]
  assign _GEN_9478 = 5'h3 == _T_938 ? welem[3] : _GEN_9477; // @[Execute.scala 117:10]
  assign _GEN_9479 = 5'h4 == _T_938 ? welem[4] : _GEN_9478; // @[Execute.scala 117:10]
  assign _GEN_9480 = 5'h5 == _T_938 ? welem[5] : _GEN_9479; // @[Execute.scala 117:10]
  assign _GEN_9481 = 5'h6 == _T_938 ? welem[6] : _GEN_9480; // @[Execute.scala 117:10]
  assign _GEN_9482 = 5'h7 == _T_938 ? welem[7] : _GEN_9481; // @[Execute.scala 117:10]
  assign _GEN_9483 = 5'h8 == _T_938 ? welem[8] : _GEN_9482; // @[Execute.scala 117:10]
  assign _GEN_9484 = 5'h9 == _T_938 ? welem[9] : _GEN_9483; // @[Execute.scala 117:10]
  assign _GEN_9485 = 5'ha == _T_938 ? welem[10] : _GEN_9484; // @[Execute.scala 117:10]
  assign _GEN_9486 = 5'hb == _T_938 ? welem[11] : _GEN_9485; // @[Execute.scala 117:10]
  assign _GEN_9487 = 5'hc == _T_938 ? welem[12] : _GEN_9486; // @[Execute.scala 117:10]
  assign _GEN_9488 = 5'hd == _T_938 ? welem[13] : _GEN_9487; // @[Execute.scala 117:10]
  assign _GEN_9489 = 5'he == _T_938 ? welem[14] : _GEN_9488; // @[Execute.scala 117:10]
  assign _GEN_9490 = 5'hf == _T_938 ? welem[15] : _GEN_9489; // @[Execute.scala 117:10]
  assign _GEN_9491 = 5'h10 == _T_938 ? welem[16] : _GEN_9490; // @[Execute.scala 117:10]
  assign _GEN_9492 = 5'h11 == _T_938 ? welem[17] : _GEN_9491; // @[Execute.scala 117:10]
  assign _GEN_9493 = 5'h12 == _T_938 ? welem[18] : _GEN_9492; // @[Execute.scala 117:10]
  assign _GEN_9494 = 5'h13 == _T_938 ? welem[19] : _GEN_9493; // @[Execute.scala 117:10]
  assign _GEN_9495 = 5'h14 == _T_938 ? welem[20] : _GEN_9494; // @[Execute.scala 117:10]
  assign _GEN_9496 = 5'h15 == _T_938 ? welem[21] : _GEN_9495; // @[Execute.scala 117:10]
  assign _GEN_9497 = 5'h16 == _T_938 ? welem[22] : _GEN_9496; // @[Execute.scala 117:10]
  assign _GEN_9498 = 5'h17 == _T_938 ? welem[23] : _GEN_9497; // @[Execute.scala 117:10]
  assign _GEN_9499 = 5'h18 == _T_938 ? welem[24] : _GEN_9498; // @[Execute.scala 117:10]
  assign _GEN_9500 = 5'h19 == _T_938 ? welem[25] : _GEN_9499; // @[Execute.scala 117:10]
  assign _GEN_9501 = 5'h1a == _T_938 ? welem[26] : _GEN_9500; // @[Execute.scala 117:10]
  assign _GEN_9502 = 5'h1b == _T_938 ? welem[27] : _GEN_9501; // @[Execute.scala 117:10]
  assign _GEN_9503 = 5'h1c == _T_938 ? welem[28] : _GEN_9502; // @[Execute.scala 117:10]
  assign _GEN_9504 = 5'h1d == _T_938 ? welem[29] : _GEN_9503; // @[Execute.scala 117:10]
  assign _GEN_9505 = 5'h1e == _T_938 ? welem[30] : _GEN_9504; // @[Execute.scala 117:10]
  assign _GEN_9506 = 5'h1f == _T_938 ? welem[31] : _GEN_9505; // @[Execute.scala 117:10]
  assign _GEN_9508 = 5'h1 == _T_940 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9509 = 5'h2 == _T_940 ? welem[2] : _GEN_9508; // @[Execute.scala 117:10]
  assign _GEN_9510 = 5'h3 == _T_940 ? welem[3] : _GEN_9509; // @[Execute.scala 117:10]
  assign _GEN_9511 = 5'h4 == _T_940 ? welem[4] : _GEN_9510; // @[Execute.scala 117:10]
  assign _GEN_9512 = 5'h5 == _T_940 ? welem[5] : _GEN_9511; // @[Execute.scala 117:10]
  assign _GEN_9513 = 5'h6 == _T_940 ? welem[6] : _GEN_9512; // @[Execute.scala 117:10]
  assign _GEN_9514 = 5'h7 == _T_940 ? welem[7] : _GEN_9513; // @[Execute.scala 117:10]
  assign _GEN_9515 = 5'h8 == _T_940 ? welem[8] : _GEN_9514; // @[Execute.scala 117:10]
  assign _GEN_9516 = 5'h9 == _T_940 ? welem[9] : _GEN_9515; // @[Execute.scala 117:10]
  assign _GEN_9517 = 5'ha == _T_940 ? welem[10] : _GEN_9516; // @[Execute.scala 117:10]
  assign _GEN_9518 = 5'hb == _T_940 ? welem[11] : _GEN_9517; // @[Execute.scala 117:10]
  assign _GEN_9519 = 5'hc == _T_940 ? welem[12] : _GEN_9518; // @[Execute.scala 117:10]
  assign _GEN_9520 = 5'hd == _T_940 ? welem[13] : _GEN_9519; // @[Execute.scala 117:10]
  assign _GEN_9521 = 5'he == _T_940 ? welem[14] : _GEN_9520; // @[Execute.scala 117:10]
  assign _GEN_9522 = 5'hf == _T_940 ? welem[15] : _GEN_9521; // @[Execute.scala 117:10]
  assign _GEN_9523 = 5'h10 == _T_940 ? welem[16] : _GEN_9522; // @[Execute.scala 117:10]
  assign _GEN_9524 = 5'h11 == _T_940 ? welem[17] : _GEN_9523; // @[Execute.scala 117:10]
  assign _GEN_9525 = 5'h12 == _T_940 ? welem[18] : _GEN_9524; // @[Execute.scala 117:10]
  assign _GEN_9526 = 5'h13 == _T_940 ? welem[19] : _GEN_9525; // @[Execute.scala 117:10]
  assign _GEN_9527 = 5'h14 == _T_940 ? welem[20] : _GEN_9526; // @[Execute.scala 117:10]
  assign _GEN_9528 = 5'h15 == _T_940 ? welem[21] : _GEN_9527; // @[Execute.scala 117:10]
  assign _GEN_9529 = 5'h16 == _T_940 ? welem[22] : _GEN_9528; // @[Execute.scala 117:10]
  assign _GEN_9530 = 5'h17 == _T_940 ? welem[23] : _GEN_9529; // @[Execute.scala 117:10]
  assign _GEN_9531 = 5'h18 == _T_940 ? welem[24] : _GEN_9530; // @[Execute.scala 117:10]
  assign _GEN_9532 = 5'h19 == _T_940 ? welem[25] : _GEN_9531; // @[Execute.scala 117:10]
  assign _GEN_9533 = 5'h1a == _T_940 ? welem[26] : _GEN_9532; // @[Execute.scala 117:10]
  assign _GEN_9534 = 5'h1b == _T_940 ? welem[27] : _GEN_9533; // @[Execute.scala 117:10]
  assign _GEN_9535 = 5'h1c == _T_940 ? welem[28] : _GEN_9534; // @[Execute.scala 117:10]
  assign _GEN_9536 = 5'h1d == _T_940 ? welem[29] : _GEN_9535; // @[Execute.scala 117:10]
  assign _GEN_9537 = 5'h1e == _T_940 ? welem[30] : _GEN_9536; // @[Execute.scala 117:10]
  assign _GEN_9538 = 5'h1f == _T_940 ? welem[31] : _GEN_9537; // @[Execute.scala 117:10]
  assign _T_941 = _T_936 ? _GEN_9506 : _GEN_9538; // @[Execute.scala 117:10]
  assign _T_942 = r[4:0] < 5'he; // @[Execute.scala 117:15]
  assign _T_944 = r[4:0] - 5'he; // @[Execute.scala 117:37]
  assign _T_946 = 5'h12 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9540 = 5'h1 == _T_944 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9541 = 5'h2 == _T_944 ? welem[2] : _GEN_9540; // @[Execute.scala 117:10]
  assign _GEN_9542 = 5'h3 == _T_944 ? welem[3] : _GEN_9541; // @[Execute.scala 117:10]
  assign _GEN_9543 = 5'h4 == _T_944 ? welem[4] : _GEN_9542; // @[Execute.scala 117:10]
  assign _GEN_9544 = 5'h5 == _T_944 ? welem[5] : _GEN_9543; // @[Execute.scala 117:10]
  assign _GEN_9545 = 5'h6 == _T_944 ? welem[6] : _GEN_9544; // @[Execute.scala 117:10]
  assign _GEN_9546 = 5'h7 == _T_944 ? welem[7] : _GEN_9545; // @[Execute.scala 117:10]
  assign _GEN_9547 = 5'h8 == _T_944 ? welem[8] : _GEN_9546; // @[Execute.scala 117:10]
  assign _GEN_9548 = 5'h9 == _T_944 ? welem[9] : _GEN_9547; // @[Execute.scala 117:10]
  assign _GEN_9549 = 5'ha == _T_944 ? welem[10] : _GEN_9548; // @[Execute.scala 117:10]
  assign _GEN_9550 = 5'hb == _T_944 ? welem[11] : _GEN_9549; // @[Execute.scala 117:10]
  assign _GEN_9551 = 5'hc == _T_944 ? welem[12] : _GEN_9550; // @[Execute.scala 117:10]
  assign _GEN_9552 = 5'hd == _T_944 ? welem[13] : _GEN_9551; // @[Execute.scala 117:10]
  assign _GEN_9553 = 5'he == _T_944 ? welem[14] : _GEN_9552; // @[Execute.scala 117:10]
  assign _GEN_9554 = 5'hf == _T_944 ? welem[15] : _GEN_9553; // @[Execute.scala 117:10]
  assign _GEN_9555 = 5'h10 == _T_944 ? welem[16] : _GEN_9554; // @[Execute.scala 117:10]
  assign _GEN_9556 = 5'h11 == _T_944 ? welem[17] : _GEN_9555; // @[Execute.scala 117:10]
  assign _GEN_9557 = 5'h12 == _T_944 ? welem[18] : _GEN_9556; // @[Execute.scala 117:10]
  assign _GEN_9558 = 5'h13 == _T_944 ? welem[19] : _GEN_9557; // @[Execute.scala 117:10]
  assign _GEN_9559 = 5'h14 == _T_944 ? welem[20] : _GEN_9558; // @[Execute.scala 117:10]
  assign _GEN_9560 = 5'h15 == _T_944 ? welem[21] : _GEN_9559; // @[Execute.scala 117:10]
  assign _GEN_9561 = 5'h16 == _T_944 ? welem[22] : _GEN_9560; // @[Execute.scala 117:10]
  assign _GEN_9562 = 5'h17 == _T_944 ? welem[23] : _GEN_9561; // @[Execute.scala 117:10]
  assign _GEN_9563 = 5'h18 == _T_944 ? welem[24] : _GEN_9562; // @[Execute.scala 117:10]
  assign _GEN_9564 = 5'h19 == _T_944 ? welem[25] : _GEN_9563; // @[Execute.scala 117:10]
  assign _GEN_9565 = 5'h1a == _T_944 ? welem[26] : _GEN_9564; // @[Execute.scala 117:10]
  assign _GEN_9566 = 5'h1b == _T_944 ? welem[27] : _GEN_9565; // @[Execute.scala 117:10]
  assign _GEN_9567 = 5'h1c == _T_944 ? welem[28] : _GEN_9566; // @[Execute.scala 117:10]
  assign _GEN_9568 = 5'h1d == _T_944 ? welem[29] : _GEN_9567; // @[Execute.scala 117:10]
  assign _GEN_9569 = 5'h1e == _T_944 ? welem[30] : _GEN_9568; // @[Execute.scala 117:10]
  assign _GEN_9570 = 5'h1f == _T_944 ? welem[31] : _GEN_9569; // @[Execute.scala 117:10]
  assign _GEN_9572 = 5'h1 == _T_946 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9573 = 5'h2 == _T_946 ? welem[2] : _GEN_9572; // @[Execute.scala 117:10]
  assign _GEN_9574 = 5'h3 == _T_946 ? welem[3] : _GEN_9573; // @[Execute.scala 117:10]
  assign _GEN_9575 = 5'h4 == _T_946 ? welem[4] : _GEN_9574; // @[Execute.scala 117:10]
  assign _GEN_9576 = 5'h5 == _T_946 ? welem[5] : _GEN_9575; // @[Execute.scala 117:10]
  assign _GEN_9577 = 5'h6 == _T_946 ? welem[6] : _GEN_9576; // @[Execute.scala 117:10]
  assign _GEN_9578 = 5'h7 == _T_946 ? welem[7] : _GEN_9577; // @[Execute.scala 117:10]
  assign _GEN_9579 = 5'h8 == _T_946 ? welem[8] : _GEN_9578; // @[Execute.scala 117:10]
  assign _GEN_9580 = 5'h9 == _T_946 ? welem[9] : _GEN_9579; // @[Execute.scala 117:10]
  assign _GEN_9581 = 5'ha == _T_946 ? welem[10] : _GEN_9580; // @[Execute.scala 117:10]
  assign _GEN_9582 = 5'hb == _T_946 ? welem[11] : _GEN_9581; // @[Execute.scala 117:10]
  assign _GEN_9583 = 5'hc == _T_946 ? welem[12] : _GEN_9582; // @[Execute.scala 117:10]
  assign _GEN_9584 = 5'hd == _T_946 ? welem[13] : _GEN_9583; // @[Execute.scala 117:10]
  assign _GEN_9585 = 5'he == _T_946 ? welem[14] : _GEN_9584; // @[Execute.scala 117:10]
  assign _GEN_9586 = 5'hf == _T_946 ? welem[15] : _GEN_9585; // @[Execute.scala 117:10]
  assign _GEN_9587 = 5'h10 == _T_946 ? welem[16] : _GEN_9586; // @[Execute.scala 117:10]
  assign _GEN_9588 = 5'h11 == _T_946 ? welem[17] : _GEN_9587; // @[Execute.scala 117:10]
  assign _GEN_9589 = 5'h12 == _T_946 ? welem[18] : _GEN_9588; // @[Execute.scala 117:10]
  assign _GEN_9590 = 5'h13 == _T_946 ? welem[19] : _GEN_9589; // @[Execute.scala 117:10]
  assign _GEN_9591 = 5'h14 == _T_946 ? welem[20] : _GEN_9590; // @[Execute.scala 117:10]
  assign _GEN_9592 = 5'h15 == _T_946 ? welem[21] : _GEN_9591; // @[Execute.scala 117:10]
  assign _GEN_9593 = 5'h16 == _T_946 ? welem[22] : _GEN_9592; // @[Execute.scala 117:10]
  assign _GEN_9594 = 5'h17 == _T_946 ? welem[23] : _GEN_9593; // @[Execute.scala 117:10]
  assign _GEN_9595 = 5'h18 == _T_946 ? welem[24] : _GEN_9594; // @[Execute.scala 117:10]
  assign _GEN_9596 = 5'h19 == _T_946 ? welem[25] : _GEN_9595; // @[Execute.scala 117:10]
  assign _GEN_9597 = 5'h1a == _T_946 ? welem[26] : _GEN_9596; // @[Execute.scala 117:10]
  assign _GEN_9598 = 5'h1b == _T_946 ? welem[27] : _GEN_9597; // @[Execute.scala 117:10]
  assign _GEN_9599 = 5'h1c == _T_946 ? welem[28] : _GEN_9598; // @[Execute.scala 117:10]
  assign _GEN_9600 = 5'h1d == _T_946 ? welem[29] : _GEN_9599; // @[Execute.scala 117:10]
  assign _GEN_9601 = 5'h1e == _T_946 ? welem[30] : _GEN_9600; // @[Execute.scala 117:10]
  assign _GEN_9602 = 5'h1f == _T_946 ? welem[31] : _GEN_9601; // @[Execute.scala 117:10]
  assign _T_947 = _T_942 ? _GEN_9570 : _GEN_9602; // @[Execute.scala 117:10]
  assign _T_948 = r[4:0] < 5'hd; // @[Execute.scala 117:15]
  assign _T_950 = r[4:0] - 5'hd; // @[Execute.scala 117:37]
  assign _T_952 = 5'h13 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9604 = 5'h1 == _T_950 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9605 = 5'h2 == _T_950 ? welem[2] : _GEN_9604; // @[Execute.scala 117:10]
  assign _GEN_9606 = 5'h3 == _T_950 ? welem[3] : _GEN_9605; // @[Execute.scala 117:10]
  assign _GEN_9607 = 5'h4 == _T_950 ? welem[4] : _GEN_9606; // @[Execute.scala 117:10]
  assign _GEN_9608 = 5'h5 == _T_950 ? welem[5] : _GEN_9607; // @[Execute.scala 117:10]
  assign _GEN_9609 = 5'h6 == _T_950 ? welem[6] : _GEN_9608; // @[Execute.scala 117:10]
  assign _GEN_9610 = 5'h7 == _T_950 ? welem[7] : _GEN_9609; // @[Execute.scala 117:10]
  assign _GEN_9611 = 5'h8 == _T_950 ? welem[8] : _GEN_9610; // @[Execute.scala 117:10]
  assign _GEN_9612 = 5'h9 == _T_950 ? welem[9] : _GEN_9611; // @[Execute.scala 117:10]
  assign _GEN_9613 = 5'ha == _T_950 ? welem[10] : _GEN_9612; // @[Execute.scala 117:10]
  assign _GEN_9614 = 5'hb == _T_950 ? welem[11] : _GEN_9613; // @[Execute.scala 117:10]
  assign _GEN_9615 = 5'hc == _T_950 ? welem[12] : _GEN_9614; // @[Execute.scala 117:10]
  assign _GEN_9616 = 5'hd == _T_950 ? welem[13] : _GEN_9615; // @[Execute.scala 117:10]
  assign _GEN_9617 = 5'he == _T_950 ? welem[14] : _GEN_9616; // @[Execute.scala 117:10]
  assign _GEN_9618 = 5'hf == _T_950 ? welem[15] : _GEN_9617; // @[Execute.scala 117:10]
  assign _GEN_9619 = 5'h10 == _T_950 ? welem[16] : _GEN_9618; // @[Execute.scala 117:10]
  assign _GEN_9620 = 5'h11 == _T_950 ? welem[17] : _GEN_9619; // @[Execute.scala 117:10]
  assign _GEN_9621 = 5'h12 == _T_950 ? welem[18] : _GEN_9620; // @[Execute.scala 117:10]
  assign _GEN_9622 = 5'h13 == _T_950 ? welem[19] : _GEN_9621; // @[Execute.scala 117:10]
  assign _GEN_9623 = 5'h14 == _T_950 ? welem[20] : _GEN_9622; // @[Execute.scala 117:10]
  assign _GEN_9624 = 5'h15 == _T_950 ? welem[21] : _GEN_9623; // @[Execute.scala 117:10]
  assign _GEN_9625 = 5'h16 == _T_950 ? welem[22] : _GEN_9624; // @[Execute.scala 117:10]
  assign _GEN_9626 = 5'h17 == _T_950 ? welem[23] : _GEN_9625; // @[Execute.scala 117:10]
  assign _GEN_9627 = 5'h18 == _T_950 ? welem[24] : _GEN_9626; // @[Execute.scala 117:10]
  assign _GEN_9628 = 5'h19 == _T_950 ? welem[25] : _GEN_9627; // @[Execute.scala 117:10]
  assign _GEN_9629 = 5'h1a == _T_950 ? welem[26] : _GEN_9628; // @[Execute.scala 117:10]
  assign _GEN_9630 = 5'h1b == _T_950 ? welem[27] : _GEN_9629; // @[Execute.scala 117:10]
  assign _GEN_9631 = 5'h1c == _T_950 ? welem[28] : _GEN_9630; // @[Execute.scala 117:10]
  assign _GEN_9632 = 5'h1d == _T_950 ? welem[29] : _GEN_9631; // @[Execute.scala 117:10]
  assign _GEN_9633 = 5'h1e == _T_950 ? welem[30] : _GEN_9632; // @[Execute.scala 117:10]
  assign _GEN_9634 = 5'h1f == _T_950 ? welem[31] : _GEN_9633; // @[Execute.scala 117:10]
  assign _GEN_9636 = 5'h1 == _T_952 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9637 = 5'h2 == _T_952 ? welem[2] : _GEN_9636; // @[Execute.scala 117:10]
  assign _GEN_9638 = 5'h3 == _T_952 ? welem[3] : _GEN_9637; // @[Execute.scala 117:10]
  assign _GEN_9639 = 5'h4 == _T_952 ? welem[4] : _GEN_9638; // @[Execute.scala 117:10]
  assign _GEN_9640 = 5'h5 == _T_952 ? welem[5] : _GEN_9639; // @[Execute.scala 117:10]
  assign _GEN_9641 = 5'h6 == _T_952 ? welem[6] : _GEN_9640; // @[Execute.scala 117:10]
  assign _GEN_9642 = 5'h7 == _T_952 ? welem[7] : _GEN_9641; // @[Execute.scala 117:10]
  assign _GEN_9643 = 5'h8 == _T_952 ? welem[8] : _GEN_9642; // @[Execute.scala 117:10]
  assign _GEN_9644 = 5'h9 == _T_952 ? welem[9] : _GEN_9643; // @[Execute.scala 117:10]
  assign _GEN_9645 = 5'ha == _T_952 ? welem[10] : _GEN_9644; // @[Execute.scala 117:10]
  assign _GEN_9646 = 5'hb == _T_952 ? welem[11] : _GEN_9645; // @[Execute.scala 117:10]
  assign _GEN_9647 = 5'hc == _T_952 ? welem[12] : _GEN_9646; // @[Execute.scala 117:10]
  assign _GEN_9648 = 5'hd == _T_952 ? welem[13] : _GEN_9647; // @[Execute.scala 117:10]
  assign _GEN_9649 = 5'he == _T_952 ? welem[14] : _GEN_9648; // @[Execute.scala 117:10]
  assign _GEN_9650 = 5'hf == _T_952 ? welem[15] : _GEN_9649; // @[Execute.scala 117:10]
  assign _GEN_9651 = 5'h10 == _T_952 ? welem[16] : _GEN_9650; // @[Execute.scala 117:10]
  assign _GEN_9652 = 5'h11 == _T_952 ? welem[17] : _GEN_9651; // @[Execute.scala 117:10]
  assign _GEN_9653 = 5'h12 == _T_952 ? welem[18] : _GEN_9652; // @[Execute.scala 117:10]
  assign _GEN_9654 = 5'h13 == _T_952 ? welem[19] : _GEN_9653; // @[Execute.scala 117:10]
  assign _GEN_9655 = 5'h14 == _T_952 ? welem[20] : _GEN_9654; // @[Execute.scala 117:10]
  assign _GEN_9656 = 5'h15 == _T_952 ? welem[21] : _GEN_9655; // @[Execute.scala 117:10]
  assign _GEN_9657 = 5'h16 == _T_952 ? welem[22] : _GEN_9656; // @[Execute.scala 117:10]
  assign _GEN_9658 = 5'h17 == _T_952 ? welem[23] : _GEN_9657; // @[Execute.scala 117:10]
  assign _GEN_9659 = 5'h18 == _T_952 ? welem[24] : _GEN_9658; // @[Execute.scala 117:10]
  assign _GEN_9660 = 5'h19 == _T_952 ? welem[25] : _GEN_9659; // @[Execute.scala 117:10]
  assign _GEN_9661 = 5'h1a == _T_952 ? welem[26] : _GEN_9660; // @[Execute.scala 117:10]
  assign _GEN_9662 = 5'h1b == _T_952 ? welem[27] : _GEN_9661; // @[Execute.scala 117:10]
  assign _GEN_9663 = 5'h1c == _T_952 ? welem[28] : _GEN_9662; // @[Execute.scala 117:10]
  assign _GEN_9664 = 5'h1d == _T_952 ? welem[29] : _GEN_9663; // @[Execute.scala 117:10]
  assign _GEN_9665 = 5'h1e == _T_952 ? welem[30] : _GEN_9664; // @[Execute.scala 117:10]
  assign _GEN_9666 = 5'h1f == _T_952 ? welem[31] : _GEN_9665; // @[Execute.scala 117:10]
  assign _T_953 = _T_948 ? _GEN_9634 : _GEN_9666; // @[Execute.scala 117:10]
  assign _T_954 = r[4:0] < 5'hc; // @[Execute.scala 117:15]
  assign _T_956 = r[4:0] - 5'hc; // @[Execute.scala 117:37]
  assign _T_958 = 5'h14 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9668 = 5'h1 == _T_956 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9669 = 5'h2 == _T_956 ? welem[2] : _GEN_9668; // @[Execute.scala 117:10]
  assign _GEN_9670 = 5'h3 == _T_956 ? welem[3] : _GEN_9669; // @[Execute.scala 117:10]
  assign _GEN_9671 = 5'h4 == _T_956 ? welem[4] : _GEN_9670; // @[Execute.scala 117:10]
  assign _GEN_9672 = 5'h5 == _T_956 ? welem[5] : _GEN_9671; // @[Execute.scala 117:10]
  assign _GEN_9673 = 5'h6 == _T_956 ? welem[6] : _GEN_9672; // @[Execute.scala 117:10]
  assign _GEN_9674 = 5'h7 == _T_956 ? welem[7] : _GEN_9673; // @[Execute.scala 117:10]
  assign _GEN_9675 = 5'h8 == _T_956 ? welem[8] : _GEN_9674; // @[Execute.scala 117:10]
  assign _GEN_9676 = 5'h9 == _T_956 ? welem[9] : _GEN_9675; // @[Execute.scala 117:10]
  assign _GEN_9677 = 5'ha == _T_956 ? welem[10] : _GEN_9676; // @[Execute.scala 117:10]
  assign _GEN_9678 = 5'hb == _T_956 ? welem[11] : _GEN_9677; // @[Execute.scala 117:10]
  assign _GEN_9679 = 5'hc == _T_956 ? welem[12] : _GEN_9678; // @[Execute.scala 117:10]
  assign _GEN_9680 = 5'hd == _T_956 ? welem[13] : _GEN_9679; // @[Execute.scala 117:10]
  assign _GEN_9681 = 5'he == _T_956 ? welem[14] : _GEN_9680; // @[Execute.scala 117:10]
  assign _GEN_9682 = 5'hf == _T_956 ? welem[15] : _GEN_9681; // @[Execute.scala 117:10]
  assign _GEN_9683 = 5'h10 == _T_956 ? welem[16] : _GEN_9682; // @[Execute.scala 117:10]
  assign _GEN_9684 = 5'h11 == _T_956 ? welem[17] : _GEN_9683; // @[Execute.scala 117:10]
  assign _GEN_9685 = 5'h12 == _T_956 ? welem[18] : _GEN_9684; // @[Execute.scala 117:10]
  assign _GEN_9686 = 5'h13 == _T_956 ? welem[19] : _GEN_9685; // @[Execute.scala 117:10]
  assign _GEN_9687 = 5'h14 == _T_956 ? welem[20] : _GEN_9686; // @[Execute.scala 117:10]
  assign _GEN_9688 = 5'h15 == _T_956 ? welem[21] : _GEN_9687; // @[Execute.scala 117:10]
  assign _GEN_9689 = 5'h16 == _T_956 ? welem[22] : _GEN_9688; // @[Execute.scala 117:10]
  assign _GEN_9690 = 5'h17 == _T_956 ? welem[23] : _GEN_9689; // @[Execute.scala 117:10]
  assign _GEN_9691 = 5'h18 == _T_956 ? welem[24] : _GEN_9690; // @[Execute.scala 117:10]
  assign _GEN_9692 = 5'h19 == _T_956 ? welem[25] : _GEN_9691; // @[Execute.scala 117:10]
  assign _GEN_9693 = 5'h1a == _T_956 ? welem[26] : _GEN_9692; // @[Execute.scala 117:10]
  assign _GEN_9694 = 5'h1b == _T_956 ? welem[27] : _GEN_9693; // @[Execute.scala 117:10]
  assign _GEN_9695 = 5'h1c == _T_956 ? welem[28] : _GEN_9694; // @[Execute.scala 117:10]
  assign _GEN_9696 = 5'h1d == _T_956 ? welem[29] : _GEN_9695; // @[Execute.scala 117:10]
  assign _GEN_9697 = 5'h1e == _T_956 ? welem[30] : _GEN_9696; // @[Execute.scala 117:10]
  assign _GEN_9698 = 5'h1f == _T_956 ? welem[31] : _GEN_9697; // @[Execute.scala 117:10]
  assign _GEN_9700 = 5'h1 == _T_958 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9701 = 5'h2 == _T_958 ? welem[2] : _GEN_9700; // @[Execute.scala 117:10]
  assign _GEN_9702 = 5'h3 == _T_958 ? welem[3] : _GEN_9701; // @[Execute.scala 117:10]
  assign _GEN_9703 = 5'h4 == _T_958 ? welem[4] : _GEN_9702; // @[Execute.scala 117:10]
  assign _GEN_9704 = 5'h5 == _T_958 ? welem[5] : _GEN_9703; // @[Execute.scala 117:10]
  assign _GEN_9705 = 5'h6 == _T_958 ? welem[6] : _GEN_9704; // @[Execute.scala 117:10]
  assign _GEN_9706 = 5'h7 == _T_958 ? welem[7] : _GEN_9705; // @[Execute.scala 117:10]
  assign _GEN_9707 = 5'h8 == _T_958 ? welem[8] : _GEN_9706; // @[Execute.scala 117:10]
  assign _GEN_9708 = 5'h9 == _T_958 ? welem[9] : _GEN_9707; // @[Execute.scala 117:10]
  assign _GEN_9709 = 5'ha == _T_958 ? welem[10] : _GEN_9708; // @[Execute.scala 117:10]
  assign _GEN_9710 = 5'hb == _T_958 ? welem[11] : _GEN_9709; // @[Execute.scala 117:10]
  assign _GEN_9711 = 5'hc == _T_958 ? welem[12] : _GEN_9710; // @[Execute.scala 117:10]
  assign _GEN_9712 = 5'hd == _T_958 ? welem[13] : _GEN_9711; // @[Execute.scala 117:10]
  assign _GEN_9713 = 5'he == _T_958 ? welem[14] : _GEN_9712; // @[Execute.scala 117:10]
  assign _GEN_9714 = 5'hf == _T_958 ? welem[15] : _GEN_9713; // @[Execute.scala 117:10]
  assign _GEN_9715 = 5'h10 == _T_958 ? welem[16] : _GEN_9714; // @[Execute.scala 117:10]
  assign _GEN_9716 = 5'h11 == _T_958 ? welem[17] : _GEN_9715; // @[Execute.scala 117:10]
  assign _GEN_9717 = 5'h12 == _T_958 ? welem[18] : _GEN_9716; // @[Execute.scala 117:10]
  assign _GEN_9718 = 5'h13 == _T_958 ? welem[19] : _GEN_9717; // @[Execute.scala 117:10]
  assign _GEN_9719 = 5'h14 == _T_958 ? welem[20] : _GEN_9718; // @[Execute.scala 117:10]
  assign _GEN_9720 = 5'h15 == _T_958 ? welem[21] : _GEN_9719; // @[Execute.scala 117:10]
  assign _GEN_9721 = 5'h16 == _T_958 ? welem[22] : _GEN_9720; // @[Execute.scala 117:10]
  assign _GEN_9722 = 5'h17 == _T_958 ? welem[23] : _GEN_9721; // @[Execute.scala 117:10]
  assign _GEN_9723 = 5'h18 == _T_958 ? welem[24] : _GEN_9722; // @[Execute.scala 117:10]
  assign _GEN_9724 = 5'h19 == _T_958 ? welem[25] : _GEN_9723; // @[Execute.scala 117:10]
  assign _GEN_9725 = 5'h1a == _T_958 ? welem[26] : _GEN_9724; // @[Execute.scala 117:10]
  assign _GEN_9726 = 5'h1b == _T_958 ? welem[27] : _GEN_9725; // @[Execute.scala 117:10]
  assign _GEN_9727 = 5'h1c == _T_958 ? welem[28] : _GEN_9726; // @[Execute.scala 117:10]
  assign _GEN_9728 = 5'h1d == _T_958 ? welem[29] : _GEN_9727; // @[Execute.scala 117:10]
  assign _GEN_9729 = 5'h1e == _T_958 ? welem[30] : _GEN_9728; // @[Execute.scala 117:10]
  assign _GEN_9730 = 5'h1f == _T_958 ? welem[31] : _GEN_9729; // @[Execute.scala 117:10]
  assign _T_959 = _T_954 ? _GEN_9698 : _GEN_9730; // @[Execute.scala 117:10]
  assign _T_960 = r[4:0] < 5'hb; // @[Execute.scala 117:15]
  assign _T_962 = r[4:0] - 5'hb; // @[Execute.scala 117:37]
  assign _T_964 = 5'h15 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9732 = 5'h1 == _T_962 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9733 = 5'h2 == _T_962 ? welem[2] : _GEN_9732; // @[Execute.scala 117:10]
  assign _GEN_9734 = 5'h3 == _T_962 ? welem[3] : _GEN_9733; // @[Execute.scala 117:10]
  assign _GEN_9735 = 5'h4 == _T_962 ? welem[4] : _GEN_9734; // @[Execute.scala 117:10]
  assign _GEN_9736 = 5'h5 == _T_962 ? welem[5] : _GEN_9735; // @[Execute.scala 117:10]
  assign _GEN_9737 = 5'h6 == _T_962 ? welem[6] : _GEN_9736; // @[Execute.scala 117:10]
  assign _GEN_9738 = 5'h7 == _T_962 ? welem[7] : _GEN_9737; // @[Execute.scala 117:10]
  assign _GEN_9739 = 5'h8 == _T_962 ? welem[8] : _GEN_9738; // @[Execute.scala 117:10]
  assign _GEN_9740 = 5'h9 == _T_962 ? welem[9] : _GEN_9739; // @[Execute.scala 117:10]
  assign _GEN_9741 = 5'ha == _T_962 ? welem[10] : _GEN_9740; // @[Execute.scala 117:10]
  assign _GEN_9742 = 5'hb == _T_962 ? welem[11] : _GEN_9741; // @[Execute.scala 117:10]
  assign _GEN_9743 = 5'hc == _T_962 ? welem[12] : _GEN_9742; // @[Execute.scala 117:10]
  assign _GEN_9744 = 5'hd == _T_962 ? welem[13] : _GEN_9743; // @[Execute.scala 117:10]
  assign _GEN_9745 = 5'he == _T_962 ? welem[14] : _GEN_9744; // @[Execute.scala 117:10]
  assign _GEN_9746 = 5'hf == _T_962 ? welem[15] : _GEN_9745; // @[Execute.scala 117:10]
  assign _GEN_9747 = 5'h10 == _T_962 ? welem[16] : _GEN_9746; // @[Execute.scala 117:10]
  assign _GEN_9748 = 5'h11 == _T_962 ? welem[17] : _GEN_9747; // @[Execute.scala 117:10]
  assign _GEN_9749 = 5'h12 == _T_962 ? welem[18] : _GEN_9748; // @[Execute.scala 117:10]
  assign _GEN_9750 = 5'h13 == _T_962 ? welem[19] : _GEN_9749; // @[Execute.scala 117:10]
  assign _GEN_9751 = 5'h14 == _T_962 ? welem[20] : _GEN_9750; // @[Execute.scala 117:10]
  assign _GEN_9752 = 5'h15 == _T_962 ? welem[21] : _GEN_9751; // @[Execute.scala 117:10]
  assign _GEN_9753 = 5'h16 == _T_962 ? welem[22] : _GEN_9752; // @[Execute.scala 117:10]
  assign _GEN_9754 = 5'h17 == _T_962 ? welem[23] : _GEN_9753; // @[Execute.scala 117:10]
  assign _GEN_9755 = 5'h18 == _T_962 ? welem[24] : _GEN_9754; // @[Execute.scala 117:10]
  assign _GEN_9756 = 5'h19 == _T_962 ? welem[25] : _GEN_9755; // @[Execute.scala 117:10]
  assign _GEN_9757 = 5'h1a == _T_962 ? welem[26] : _GEN_9756; // @[Execute.scala 117:10]
  assign _GEN_9758 = 5'h1b == _T_962 ? welem[27] : _GEN_9757; // @[Execute.scala 117:10]
  assign _GEN_9759 = 5'h1c == _T_962 ? welem[28] : _GEN_9758; // @[Execute.scala 117:10]
  assign _GEN_9760 = 5'h1d == _T_962 ? welem[29] : _GEN_9759; // @[Execute.scala 117:10]
  assign _GEN_9761 = 5'h1e == _T_962 ? welem[30] : _GEN_9760; // @[Execute.scala 117:10]
  assign _GEN_9762 = 5'h1f == _T_962 ? welem[31] : _GEN_9761; // @[Execute.scala 117:10]
  assign _GEN_9764 = 5'h1 == _T_964 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9765 = 5'h2 == _T_964 ? welem[2] : _GEN_9764; // @[Execute.scala 117:10]
  assign _GEN_9766 = 5'h3 == _T_964 ? welem[3] : _GEN_9765; // @[Execute.scala 117:10]
  assign _GEN_9767 = 5'h4 == _T_964 ? welem[4] : _GEN_9766; // @[Execute.scala 117:10]
  assign _GEN_9768 = 5'h5 == _T_964 ? welem[5] : _GEN_9767; // @[Execute.scala 117:10]
  assign _GEN_9769 = 5'h6 == _T_964 ? welem[6] : _GEN_9768; // @[Execute.scala 117:10]
  assign _GEN_9770 = 5'h7 == _T_964 ? welem[7] : _GEN_9769; // @[Execute.scala 117:10]
  assign _GEN_9771 = 5'h8 == _T_964 ? welem[8] : _GEN_9770; // @[Execute.scala 117:10]
  assign _GEN_9772 = 5'h9 == _T_964 ? welem[9] : _GEN_9771; // @[Execute.scala 117:10]
  assign _GEN_9773 = 5'ha == _T_964 ? welem[10] : _GEN_9772; // @[Execute.scala 117:10]
  assign _GEN_9774 = 5'hb == _T_964 ? welem[11] : _GEN_9773; // @[Execute.scala 117:10]
  assign _GEN_9775 = 5'hc == _T_964 ? welem[12] : _GEN_9774; // @[Execute.scala 117:10]
  assign _GEN_9776 = 5'hd == _T_964 ? welem[13] : _GEN_9775; // @[Execute.scala 117:10]
  assign _GEN_9777 = 5'he == _T_964 ? welem[14] : _GEN_9776; // @[Execute.scala 117:10]
  assign _GEN_9778 = 5'hf == _T_964 ? welem[15] : _GEN_9777; // @[Execute.scala 117:10]
  assign _GEN_9779 = 5'h10 == _T_964 ? welem[16] : _GEN_9778; // @[Execute.scala 117:10]
  assign _GEN_9780 = 5'h11 == _T_964 ? welem[17] : _GEN_9779; // @[Execute.scala 117:10]
  assign _GEN_9781 = 5'h12 == _T_964 ? welem[18] : _GEN_9780; // @[Execute.scala 117:10]
  assign _GEN_9782 = 5'h13 == _T_964 ? welem[19] : _GEN_9781; // @[Execute.scala 117:10]
  assign _GEN_9783 = 5'h14 == _T_964 ? welem[20] : _GEN_9782; // @[Execute.scala 117:10]
  assign _GEN_9784 = 5'h15 == _T_964 ? welem[21] : _GEN_9783; // @[Execute.scala 117:10]
  assign _GEN_9785 = 5'h16 == _T_964 ? welem[22] : _GEN_9784; // @[Execute.scala 117:10]
  assign _GEN_9786 = 5'h17 == _T_964 ? welem[23] : _GEN_9785; // @[Execute.scala 117:10]
  assign _GEN_9787 = 5'h18 == _T_964 ? welem[24] : _GEN_9786; // @[Execute.scala 117:10]
  assign _GEN_9788 = 5'h19 == _T_964 ? welem[25] : _GEN_9787; // @[Execute.scala 117:10]
  assign _GEN_9789 = 5'h1a == _T_964 ? welem[26] : _GEN_9788; // @[Execute.scala 117:10]
  assign _GEN_9790 = 5'h1b == _T_964 ? welem[27] : _GEN_9789; // @[Execute.scala 117:10]
  assign _GEN_9791 = 5'h1c == _T_964 ? welem[28] : _GEN_9790; // @[Execute.scala 117:10]
  assign _GEN_9792 = 5'h1d == _T_964 ? welem[29] : _GEN_9791; // @[Execute.scala 117:10]
  assign _GEN_9793 = 5'h1e == _T_964 ? welem[30] : _GEN_9792; // @[Execute.scala 117:10]
  assign _GEN_9794 = 5'h1f == _T_964 ? welem[31] : _GEN_9793; // @[Execute.scala 117:10]
  assign _T_965 = _T_960 ? _GEN_9762 : _GEN_9794; // @[Execute.scala 117:10]
  assign _T_966 = r[4:0] < 5'ha; // @[Execute.scala 117:15]
  assign _T_968 = r[4:0] - 5'ha; // @[Execute.scala 117:37]
  assign _T_970 = 5'h16 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9796 = 5'h1 == _T_968 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9797 = 5'h2 == _T_968 ? welem[2] : _GEN_9796; // @[Execute.scala 117:10]
  assign _GEN_9798 = 5'h3 == _T_968 ? welem[3] : _GEN_9797; // @[Execute.scala 117:10]
  assign _GEN_9799 = 5'h4 == _T_968 ? welem[4] : _GEN_9798; // @[Execute.scala 117:10]
  assign _GEN_9800 = 5'h5 == _T_968 ? welem[5] : _GEN_9799; // @[Execute.scala 117:10]
  assign _GEN_9801 = 5'h6 == _T_968 ? welem[6] : _GEN_9800; // @[Execute.scala 117:10]
  assign _GEN_9802 = 5'h7 == _T_968 ? welem[7] : _GEN_9801; // @[Execute.scala 117:10]
  assign _GEN_9803 = 5'h8 == _T_968 ? welem[8] : _GEN_9802; // @[Execute.scala 117:10]
  assign _GEN_9804 = 5'h9 == _T_968 ? welem[9] : _GEN_9803; // @[Execute.scala 117:10]
  assign _GEN_9805 = 5'ha == _T_968 ? welem[10] : _GEN_9804; // @[Execute.scala 117:10]
  assign _GEN_9806 = 5'hb == _T_968 ? welem[11] : _GEN_9805; // @[Execute.scala 117:10]
  assign _GEN_9807 = 5'hc == _T_968 ? welem[12] : _GEN_9806; // @[Execute.scala 117:10]
  assign _GEN_9808 = 5'hd == _T_968 ? welem[13] : _GEN_9807; // @[Execute.scala 117:10]
  assign _GEN_9809 = 5'he == _T_968 ? welem[14] : _GEN_9808; // @[Execute.scala 117:10]
  assign _GEN_9810 = 5'hf == _T_968 ? welem[15] : _GEN_9809; // @[Execute.scala 117:10]
  assign _GEN_9811 = 5'h10 == _T_968 ? welem[16] : _GEN_9810; // @[Execute.scala 117:10]
  assign _GEN_9812 = 5'h11 == _T_968 ? welem[17] : _GEN_9811; // @[Execute.scala 117:10]
  assign _GEN_9813 = 5'h12 == _T_968 ? welem[18] : _GEN_9812; // @[Execute.scala 117:10]
  assign _GEN_9814 = 5'h13 == _T_968 ? welem[19] : _GEN_9813; // @[Execute.scala 117:10]
  assign _GEN_9815 = 5'h14 == _T_968 ? welem[20] : _GEN_9814; // @[Execute.scala 117:10]
  assign _GEN_9816 = 5'h15 == _T_968 ? welem[21] : _GEN_9815; // @[Execute.scala 117:10]
  assign _GEN_9817 = 5'h16 == _T_968 ? welem[22] : _GEN_9816; // @[Execute.scala 117:10]
  assign _GEN_9818 = 5'h17 == _T_968 ? welem[23] : _GEN_9817; // @[Execute.scala 117:10]
  assign _GEN_9819 = 5'h18 == _T_968 ? welem[24] : _GEN_9818; // @[Execute.scala 117:10]
  assign _GEN_9820 = 5'h19 == _T_968 ? welem[25] : _GEN_9819; // @[Execute.scala 117:10]
  assign _GEN_9821 = 5'h1a == _T_968 ? welem[26] : _GEN_9820; // @[Execute.scala 117:10]
  assign _GEN_9822 = 5'h1b == _T_968 ? welem[27] : _GEN_9821; // @[Execute.scala 117:10]
  assign _GEN_9823 = 5'h1c == _T_968 ? welem[28] : _GEN_9822; // @[Execute.scala 117:10]
  assign _GEN_9824 = 5'h1d == _T_968 ? welem[29] : _GEN_9823; // @[Execute.scala 117:10]
  assign _GEN_9825 = 5'h1e == _T_968 ? welem[30] : _GEN_9824; // @[Execute.scala 117:10]
  assign _GEN_9826 = 5'h1f == _T_968 ? welem[31] : _GEN_9825; // @[Execute.scala 117:10]
  assign _GEN_9828 = 5'h1 == _T_970 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9829 = 5'h2 == _T_970 ? welem[2] : _GEN_9828; // @[Execute.scala 117:10]
  assign _GEN_9830 = 5'h3 == _T_970 ? welem[3] : _GEN_9829; // @[Execute.scala 117:10]
  assign _GEN_9831 = 5'h4 == _T_970 ? welem[4] : _GEN_9830; // @[Execute.scala 117:10]
  assign _GEN_9832 = 5'h5 == _T_970 ? welem[5] : _GEN_9831; // @[Execute.scala 117:10]
  assign _GEN_9833 = 5'h6 == _T_970 ? welem[6] : _GEN_9832; // @[Execute.scala 117:10]
  assign _GEN_9834 = 5'h7 == _T_970 ? welem[7] : _GEN_9833; // @[Execute.scala 117:10]
  assign _GEN_9835 = 5'h8 == _T_970 ? welem[8] : _GEN_9834; // @[Execute.scala 117:10]
  assign _GEN_9836 = 5'h9 == _T_970 ? welem[9] : _GEN_9835; // @[Execute.scala 117:10]
  assign _GEN_9837 = 5'ha == _T_970 ? welem[10] : _GEN_9836; // @[Execute.scala 117:10]
  assign _GEN_9838 = 5'hb == _T_970 ? welem[11] : _GEN_9837; // @[Execute.scala 117:10]
  assign _GEN_9839 = 5'hc == _T_970 ? welem[12] : _GEN_9838; // @[Execute.scala 117:10]
  assign _GEN_9840 = 5'hd == _T_970 ? welem[13] : _GEN_9839; // @[Execute.scala 117:10]
  assign _GEN_9841 = 5'he == _T_970 ? welem[14] : _GEN_9840; // @[Execute.scala 117:10]
  assign _GEN_9842 = 5'hf == _T_970 ? welem[15] : _GEN_9841; // @[Execute.scala 117:10]
  assign _GEN_9843 = 5'h10 == _T_970 ? welem[16] : _GEN_9842; // @[Execute.scala 117:10]
  assign _GEN_9844 = 5'h11 == _T_970 ? welem[17] : _GEN_9843; // @[Execute.scala 117:10]
  assign _GEN_9845 = 5'h12 == _T_970 ? welem[18] : _GEN_9844; // @[Execute.scala 117:10]
  assign _GEN_9846 = 5'h13 == _T_970 ? welem[19] : _GEN_9845; // @[Execute.scala 117:10]
  assign _GEN_9847 = 5'h14 == _T_970 ? welem[20] : _GEN_9846; // @[Execute.scala 117:10]
  assign _GEN_9848 = 5'h15 == _T_970 ? welem[21] : _GEN_9847; // @[Execute.scala 117:10]
  assign _GEN_9849 = 5'h16 == _T_970 ? welem[22] : _GEN_9848; // @[Execute.scala 117:10]
  assign _GEN_9850 = 5'h17 == _T_970 ? welem[23] : _GEN_9849; // @[Execute.scala 117:10]
  assign _GEN_9851 = 5'h18 == _T_970 ? welem[24] : _GEN_9850; // @[Execute.scala 117:10]
  assign _GEN_9852 = 5'h19 == _T_970 ? welem[25] : _GEN_9851; // @[Execute.scala 117:10]
  assign _GEN_9853 = 5'h1a == _T_970 ? welem[26] : _GEN_9852; // @[Execute.scala 117:10]
  assign _GEN_9854 = 5'h1b == _T_970 ? welem[27] : _GEN_9853; // @[Execute.scala 117:10]
  assign _GEN_9855 = 5'h1c == _T_970 ? welem[28] : _GEN_9854; // @[Execute.scala 117:10]
  assign _GEN_9856 = 5'h1d == _T_970 ? welem[29] : _GEN_9855; // @[Execute.scala 117:10]
  assign _GEN_9857 = 5'h1e == _T_970 ? welem[30] : _GEN_9856; // @[Execute.scala 117:10]
  assign _GEN_9858 = 5'h1f == _T_970 ? welem[31] : _GEN_9857; // @[Execute.scala 117:10]
  assign _T_971 = _T_966 ? _GEN_9826 : _GEN_9858; // @[Execute.scala 117:10]
  assign _T_972 = r[4:0] < 5'h9; // @[Execute.scala 117:15]
  assign _T_974 = r[4:0] - 5'h9; // @[Execute.scala 117:37]
  assign _T_976 = 5'h17 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9860 = 5'h1 == _T_974 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9861 = 5'h2 == _T_974 ? welem[2] : _GEN_9860; // @[Execute.scala 117:10]
  assign _GEN_9862 = 5'h3 == _T_974 ? welem[3] : _GEN_9861; // @[Execute.scala 117:10]
  assign _GEN_9863 = 5'h4 == _T_974 ? welem[4] : _GEN_9862; // @[Execute.scala 117:10]
  assign _GEN_9864 = 5'h5 == _T_974 ? welem[5] : _GEN_9863; // @[Execute.scala 117:10]
  assign _GEN_9865 = 5'h6 == _T_974 ? welem[6] : _GEN_9864; // @[Execute.scala 117:10]
  assign _GEN_9866 = 5'h7 == _T_974 ? welem[7] : _GEN_9865; // @[Execute.scala 117:10]
  assign _GEN_9867 = 5'h8 == _T_974 ? welem[8] : _GEN_9866; // @[Execute.scala 117:10]
  assign _GEN_9868 = 5'h9 == _T_974 ? welem[9] : _GEN_9867; // @[Execute.scala 117:10]
  assign _GEN_9869 = 5'ha == _T_974 ? welem[10] : _GEN_9868; // @[Execute.scala 117:10]
  assign _GEN_9870 = 5'hb == _T_974 ? welem[11] : _GEN_9869; // @[Execute.scala 117:10]
  assign _GEN_9871 = 5'hc == _T_974 ? welem[12] : _GEN_9870; // @[Execute.scala 117:10]
  assign _GEN_9872 = 5'hd == _T_974 ? welem[13] : _GEN_9871; // @[Execute.scala 117:10]
  assign _GEN_9873 = 5'he == _T_974 ? welem[14] : _GEN_9872; // @[Execute.scala 117:10]
  assign _GEN_9874 = 5'hf == _T_974 ? welem[15] : _GEN_9873; // @[Execute.scala 117:10]
  assign _GEN_9875 = 5'h10 == _T_974 ? welem[16] : _GEN_9874; // @[Execute.scala 117:10]
  assign _GEN_9876 = 5'h11 == _T_974 ? welem[17] : _GEN_9875; // @[Execute.scala 117:10]
  assign _GEN_9877 = 5'h12 == _T_974 ? welem[18] : _GEN_9876; // @[Execute.scala 117:10]
  assign _GEN_9878 = 5'h13 == _T_974 ? welem[19] : _GEN_9877; // @[Execute.scala 117:10]
  assign _GEN_9879 = 5'h14 == _T_974 ? welem[20] : _GEN_9878; // @[Execute.scala 117:10]
  assign _GEN_9880 = 5'h15 == _T_974 ? welem[21] : _GEN_9879; // @[Execute.scala 117:10]
  assign _GEN_9881 = 5'h16 == _T_974 ? welem[22] : _GEN_9880; // @[Execute.scala 117:10]
  assign _GEN_9882 = 5'h17 == _T_974 ? welem[23] : _GEN_9881; // @[Execute.scala 117:10]
  assign _GEN_9883 = 5'h18 == _T_974 ? welem[24] : _GEN_9882; // @[Execute.scala 117:10]
  assign _GEN_9884 = 5'h19 == _T_974 ? welem[25] : _GEN_9883; // @[Execute.scala 117:10]
  assign _GEN_9885 = 5'h1a == _T_974 ? welem[26] : _GEN_9884; // @[Execute.scala 117:10]
  assign _GEN_9886 = 5'h1b == _T_974 ? welem[27] : _GEN_9885; // @[Execute.scala 117:10]
  assign _GEN_9887 = 5'h1c == _T_974 ? welem[28] : _GEN_9886; // @[Execute.scala 117:10]
  assign _GEN_9888 = 5'h1d == _T_974 ? welem[29] : _GEN_9887; // @[Execute.scala 117:10]
  assign _GEN_9889 = 5'h1e == _T_974 ? welem[30] : _GEN_9888; // @[Execute.scala 117:10]
  assign _GEN_9890 = 5'h1f == _T_974 ? welem[31] : _GEN_9889; // @[Execute.scala 117:10]
  assign _GEN_9892 = 5'h1 == _T_976 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9893 = 5'h2 == _T_976 ? welem[2] : _GEN_9892; // @[Execute.scala 117:10]
  assign _GEN_9894 = 5'h3 == _T_976 ? welem[3] : _GEN_9893; // @[Execute.scala 117:10]
  assign _GEN_9895 = 5'h4 == _T_976 ? welem[4] : _GEN_9894; // @[Execute.scala 117:10]
  assign _GEN_9896 = 5'h5 == _T_976 ? welem[5] : _GEN_9895; // @[Execute.scala 117:10]
  assign _GEN_9897 = 5'h6 == _T_976 ? welem[6] : _GEN_9896; // @[Execute.scala 117:10]
  assign _GEN_9898 = 5'h7 == _T_976 ? welem[7] : _GEN_9897; // @[Execute.scala 117:10]
  assign _GEN_9899 = 5'h8 == _T_976 ? welem[8] : _GEN_9898; // @[Execute.scala 117:10]
  assign _GEN_9900 = 5'h9 == _T_976 ? welem[9] : _GEN_9899; // @[Execute.scala 117:10]
  assign _GEN_9901 = 5'ha == _T_976 ? welem[10] : _GEN_9900; // @[Execute.scala 117:10]
  assign _GEN_9902 = 5'hb == _T_976 ? welem[11] : _GEN_9901; // @[Execute.scala 117:10]
  assign _GEN_9903 = 5'hc == _T_976 ? welem[12] : _GEN_9902; // @[Execute.scala 117:10]
  assign _GEN_9904 = 5'hd == _T_976 ? welem[13] : _GEN_9903; // @[Execute.scala 117:10]
  assign _GEN_9905 = 5'he == _T_976 ? welem[14] : _GEN_9904; // @[Execute.scala 117:10]
  assign _GEN_9906 = 5'hf == _T_976 ? welem[15] : _GEN_9905; // @[Execute.scala 117:10]
  assign _GEN_9907 = 5'h10 == _T_976 ? welem[16] : _GEN_9906; // @[Execute.scala 117:10]
  assign _GEN_9908 = 5'h11 == _T_976 ? welem[17] : _GEN_9907; // @[Execute.scala 117:10]
  assign _GEN_9909 = 5'h12 == _T_976 ? welem[18] : _GEN_9908; // @[Execute.scala 117:10]
  assign _GEN_9910 = 5'h13 == _T_976 ? welem[19] : _GEN_9909; // @[Execute.scala 117:10]
  assign _GEN_9911 = 5'h14 == _T_976 ? welem[20] : _GEN_9910; // @[Execute.scala 117:10]
  assign _GEN_9912 = 5'h15 == _T_976 ? welem[21] : _GEN_9911; // @[Execute.scala 117:10]
  assign _GEN_9913 = 5'h16 == _T_976 ? welem[22] : _GEN_9912; // @[Execute.scala 117:10]
  assign _GEN_9914 = 5'h17 == _T_976 ? welem[23] : _GEN_9913; // @[Execute.scala 117:10]
  assign _GEN_9915 = 5'h18 == _T_976 ? welem[24] : _GEN_9914; // @[Execute.scala 117:10]
  assign _GEN_9916 = 5'h19 == _T_976 ? welem[25] : _GEN_9915; // @[Execute.scala 117:10]
  assign _GEN_9917 = 5'h1a == _T_976 ? welem[26] : _GEN_9916; // @[Execute.scala 117:10]
  assign _GEN_9918 = 5'h1b == _T_976 ? welem[27] : _GEN_9917; // @[Execute.scala 117:10]
  assign _GEN_9919 = 5'h1c == _T_976 ? welem[28] : _GEN_9918; // @[Execute.scala 117:10]
  assign _GEN_9920 = 5'h1d == _T_976 ? welem[29] : _GEN_9919; // @[Execute.scala 117:10]
  assign _GEN_9921 = 5'h1e == _T_976 ? welem[30] : _GEN_9920; // @[Execute.scala 117:10]
  assign _GEN_9922 = 5'h1f == _T_976 ? welem[31] : _GEN_9921; // @[Execute.scala 117:10]
  assign _T_977 = _T_972 ? _GEN_9890 : _GEN_9922; // @[Execute.scala 117:10]
  assign _T_978 = r[4:0] < 5'h8; // @[Execute.scala 117:15]
  assign _T_980 = r[4:0] - 5'h8; // @[Execute.scala 117:37]
  assign _T_982 = 5'h18 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9924 = 5'h1 == _T_980 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9925 = 5'h2 == _T_980 ? welem[2] : _GEN_9924; // @[Execute.scala 117:10]
  assign _GEN_9926 = 5'h3 == _T_980 ? welem[3] : _GEN_9925; // @[Execute.scala 117:10]
  assign _GEN_9927 = 5'h4 == _T_980 ? welem[4] : _GEN_9926; // @[Execute.scala 117:10]
  assign _GEN_9928 = 5'h5 == _T_980 ? welem[5] : _GEN_9927; // @[Execute.scala 117:10]
  assign _GEN_9929 = 5'h6 == _T_980 ? welem[6] : _GEN_9928; // @[Execute.scala 117:10]
  assign _GEN_9930 = 5'h7 == _T_980 ? welem[7] : _GEN_9929; // @[Execute.scala 117:10]
  assign _GEN_9931 = 5'h8 == _T_980 ? welem[8] : _GEN_9930; // @[Execute.scala 117:10]
  assign _GEN_9932 = 5'h9 == _T_980 ? welem[9] : _GEN_9931; // @[Execute.scala 117:10]
  assign _GEN_9933 = 5'ha == _T_980 ? welem[10] : _GEN_9932; // @[Execute.scala 117:10]
  assign _GEN_9934 = 5'hb == _T_980 ? welem[11] : _GEN_9933; // @[Execute.scala 117:10]
  assign _GEN_9935 = 5'hc == _T_980 ? welem[12] : _GEN_9934; // @[Execute.scala 117:10]
  assign _GEN_9936 = 5'hd == _T_980 ? welem[13] : _GEN_9935; // @[Execute.scala 117:10]
  assign _GEN_9937 = 5'he == _T_980 ? welem[14] : _GEN_9936; // @[Execute.scala 117:10]
  assign _GEN_9938 = 5'hf == _T_980 ? welem[15] : _GEN_9937; // @[Execute.scala 117:10]
  assign _GEN_9939 = 5'h10 == _T_980 ? welem[16] : _GEN_9938; // @[Execute.scala 117:10]
  assign _GEN_9940 = 5'h11 == _T_980 ? welem[17] : _GEN_9939; // @[Execute.scala 117:10]
  assign _GEN_9941 = 5'h12 == _T_980 ? welem[18] : _GEN_9940; // @[Execute.scala 117:10]
  assign _GEN_9942 = 5'h13 == _T_980 ? welem[19] : _GEN_9941; // @[Execute.scala 117:10]
  assign _GEN_9943 = 5'h14 == _T_980 ? welem[20] : _GEN_9942; // @[Execute.scala 117:10]
  assign _GEN_9944 = 5'h15 == _T_980 ? welem[21] : _GEN_9943; // @[Execute.scala 117:10]
  assign _GEN_9945 = 5'h16 == _T_980 ? welem[22] : _GEN_9944; // @[Execute.scala 117:10]
  assign _GEN_9946 = 5'h17 == _T_980 ? welem[23] : _GEN_9945; // @[Execute.scala 117:10]
  assign _GEN_9947 = 5'h18 == _T_980 ? welem[24] : _GEN_9946; // @[Execute.scala 117:10]
  assign _GEN_9948 = 5'h19 == _T_980 ? welem[25] : _GEN_9947; // @[Execute.scala 117:10]
  assign _GEN_9949 = 5'h1a == _T_980 ? welem[26] : _GEN_9948; // @[Execute.scala 117:10]
  assign _GEN_9950 = 5'h1b == _T_980 ? welem[27] : _GEN_9949; // @[Execute.scala 117:10]
  assign _GEN_9951 = 5'h1c == _T_980 ? welem[28] : _GEN_9950; // @[Execute.scala 117:10]
  assign _GEN_9952 = 5'h1d == _T_980 ? welem[29] : _GEN_9951; // @[Execute.scala 117:10]
  assign _GEN_9953 = 5'h1e == _T_980 ? welem[30] : _GEN_9952; // @[Execute.scala 117:10]
  assign _GEN_9954 = 5'h1f == _T_980 ? welem[31] : _GEN_9953; // @[Execute.scala 117:10]
  assign _GEN_9956 = 5'h1 == _T_982 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9957 = 5'h2 == _T_982 ? welem[2] : _GEN_9956; // @[Execute.scala 117:10]
  assign _GEN_9958 = 5'h3 == _T_982 ? welem[3] : _GEN_9957; // @[Execute.scala 117:10]
  assign _GEN_9959 = 5'h4 == _T_982 ? welem[4] : _GEN_9958; // @[Execute.scala 117:10]
  assign _GEN_9960 = 5'h5 == _T_982 ? welem[5] : _GEN_9959; // @[Execute.scala 117:10]
  assign _GEN_9961 = 5'h6 == _T_982 ? welem[6] : _GEN_9960; // @[Execute.scala 117:10]
  assign _GEN_9962 = 5'h7 == _T_982 ? welem[7] : _GEN_9961; // @[Execute.scala 117:10]
  assign _GEN_9963 = 5'h8 == _T_982 ? welem[8] : _GEN_9962; // @[Execute.scala 117:10]
  assign _GEN_9964 = 5'h9 == _T_982 ? welem[9] : _GEN_9963; // @[Execute.scala 117:10]
  assign _GEN_9965 = 5'ha == _T_982 ? welem[10] : _GEN_9964; // @[Execute.scala 117:10]
  assign _GEN_9966 = 5'hb == _T_982 ? welem[11] : _GEN_9965; // @[Execute.scala 117:10]
  assign _GEN_9967 = 5'hc == _T_982 ? welem[12] : _GEN_9966; // @[Execute.scala 117:10]
  assign _GEN_9968 = 5'hd == _T_982 ? welem[13] : _GEN_9967; // @[Execute.scala 117:10]
  assign _GEN_9969 = 5'he == _T_982 ? welem[14] : _GEN_9968; // @[Execute.scala 117:10]
  assign _GEN_9970 = 5'hf == _T_982 ? welem[15] : _GEN_9969; // @[Execute.scala 117:10]
  assign _GEN_9971 = 5'h10 == _T_982 ? welem[16] : _GEN_9970; // @[Execute.scala 117:10]
  assign _GEN_9972 = 5'h11 == _T_982 ? welem[17] : _GEN_9971; // @[Execute.scala 117:10]
  assign _GEN_9973 = 5'h12 == _T_982 ? welem[18] : _GEN_9972; // @[Execute.scala 117:10]
  assign _GEN_9974 = 5'h13 == _T_982 ? welem[19] : _GEN_9973; // @[Execute.scala 117:10]
  assign _GEN_9975 = 5'h14 == _T_982 ? welem[20] : _GEN_9974; // @[Execute.scala 117:10]
  assign _GEN_9976 = 5'h15 == _T_982 ? welem[21] : _GEN_9975; // @[Execute.scala 117:10]
  assign _GEN_9977 = 5'h16 == _T_982 ? welem[22] : _GEN_9976; // @[Execute.scala 117:10]
  assign _GEN_9978 = 5'h17 == _T_982 ? welem[23] : _GEN_9977; // @[Execute.scala 117:10]
  assign _GEN_9979 = 5'h18 == _T_982 ? welem[24] : _GEN_9978; // @[Execute.scala 117:10]
  assign _GEN_9980 = 5'h19 == _T_982 ? welem[25] : _GEN_9979; // @[Execute.scala 117:10]
  assign _GEN_9981 = 5'h1a == _T_982 ? welem[26] : _GEN_9980; // @[Execute.scala 117:10]
  assign _GEN_9982 = 5'h1b == _T_982 ? welem[27] : _GEN_9981; // @[Execute.scala 117:10]
  assign _GEN_9983 = 5'h1c == _T_982 ? welem[28] : _GEN_9982; // @[Execute.scala 117:10]
  assign _GEN_9984 = 5'h1d == _T_982 ? welem[29] : _GEN_9983; // @[Execute.scala 117:10]
  assign _GEN_9985 = 5'h1e == _T_982 ? welem[30] : _GEN_9984; // @[Execute.scala 117:10]
  assign _GEN_9986 = 5'h1f == _T_982 ? welem[31] : _GEN_9985; // @[Execute.scala 117:10]
  assign _T_983 = _T_978 ? _GEN_9954 : _GEN_9986; // @[Execute.scala 117:10]
  assign _T_984 = r[4:0] < 5'h7; // @[Execute.scala 117:15]
  assign _T_986 = r[4:0] - 5'h7; // @[Execute.scala 117:37]
  assign _T_988 = 5'h19 + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_9988 = 5'h1 == _T_986 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_9989 = 5'h2 == _T_986 ? welem[2] : _GEN_9988; // @[Execute.scala 117:10]
  assign _GEN_9990 = 5'h3 == _T_986 ? welem[3] : _GEN_9989; // @[Execute.scala 117:10]
  assign _GEN_9991 = 5'h4 == _T_986 ? welem[4] : _GEN_9990; // @[Execute.scala 117:10]
  assign _GEN_9992 = 5'h5 == _T_986 ? welem[5] : _GEN_9991; // @[Execute.scala 117:10]
  assign _GEN_9993 = 5'h6 == _T_986 ? welem[6] : _GEN_9992; // @[Execute.scala 117:10]
  assign _GEN_9994 = 5'h7 == _T_986 ? welem[7] : _GEN_9993; // @[Execute.scala 117:10]
  assign _GEN_9995 = 5'h8 == _T_986 ? welem[8] : _GEN_9994; // @[Execute.scala 117:10]
  assign _GEN_9996 = 5'h9 == _T_986 ? welem[9] : _GEN_9995; // @[Execute.scala 117:10]
  assign _GEN_9997 = 5'ha == _T_986 ? welem[10] : _GEN_9996; // @[Execute.scala 117:10]
  assign _GEN_9998 = 5'hb == _T_986 ? welem[11] : _GEN_9997; // @[Execute.scala 117:10]
  assign _GEN_9999 = 5'hc == _T_986 ? welem[12] : _GEN_9998; // @[Execute.scala 117:10]
  assign _GEN_10000 = 5'hd == _T_986 ? welem[13] : _GEN_9999; // @[Execute.scala 117:10]
  assign _GEN_10001 = 5'he == _T_986 ? welem[14] : _GEN_10000; // @[Execute.scala 117:10]
  assign _GEN_10002 = 5'hf == _T_986 ? welem[15] : _GEN_10001; // @[Execute.scala 117:10]
  assign _GEN_10003 = 5'h10 == _T_986 ? welem[16] : _GEN_10002; // @[Execute.scala 117:10]
  assign _GEN_10004 = 5'h11 == _T_986 ? welem[17] : _GEN_10003; // @[Execute.scala 117:10]
  assign _GEN_10005 = 5'h12 == _T_986 ? welem[18] : _GEN_10004; // @[Execute.scala 117:10]
  assign _GEN_10006 = 5'h13 == _T_986 ? welem[19] : _GEN_10005; // @[Execute.scala 117:10]
  assign _GEN_10007 = 5'h14 == _T_986 ? welem[20] : _GEN_10006; // @[Execute.scala 117:10]
  assign _GEN_10008 = 5'h15 == _T_986 ? welem[21] : _GEN_10007; // @[Execute.scala 117:10]
  assign _GEN_10009 = 5'h16 == _T_986 ? welem[22] : _GEN_10008; // @[Execute.scala 117:10]
  assign _GEN_10010 = 5'h17 == _T_986 ? welem[23] : _GEN_10009; // @[Execute.scala 117:10]
  assign _GEN_10011 = 5'h18 == _T_986 ? welem[24] : _GEN_10010; // @[Execute.scala 117:10]
  assign _GEN_10012 = 5'h19 == _T_986 ? welem[25] : _GEN_10011; // @[Execute.scala 117:10]
  assign _GEN_10013 = 5'h1a == _T_986 ? welem[26] : _GEN_10012; // @[Execute.scala 117:10]
  assign _GEN_10014 = 5'h1b == _T_986 ? welem[27] : _GEN_10013; // @[Execute.scala 117:10]
  assign _GEN_10015 = 5'h1c == _T_986 ? welem[28] : _GEN_10014; // @[Execute.scala 117:10]
  assign _GEN_10016 = 5'h1d == _T_986 ? welem[29] : _GEN_10015; // @[Execute.scala 117:10]
  assign _GEN_10017 = 5'h1e == _T_986 ? welem[30] : _GEN_10016; // @[Execute.scala 117:10]
  assign _GEN_10018 = 5'h1f == _T_986 ? welem[31] : _GEN_10017; // @[Execute.scala 117:10]
  assign _GEN_10020 = 5'h1 == _T_988 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10021 = 5'h2 == _T_988 ? welem[2] : _GEN_10020; // @[Execute.scala 117:10]
  assign _GEN_10022 = 5'h3 == _T_988 ? welem[3] : _GEN_10021; // @[Execute.scala 117:10]
  assign _GEN_10023 = 5'h4 == _T_988 ? welem[4] : _GEN_10022; // @[Execute.scala 117:10]
  assign _GEN_10024 = 5'h5 == _T_988 ? welem[5] : _GEN_10023; // @[Execute.scala 117:10]
  assign _GEN_10025 = 5'h6 == _T_988 ? welem[6] : _GEN_10024; // @[Execute.scala 117:10]
  assign _GEN_10026 = 5'h7 == _T_988 ? welem[7] : _GEN_10025; // @[Execute.scala 117:10]
  assign _GEN_10027 = 5'h8 == _T_988 ? welem[8] : _GEN_10026; // @[Execute.scala 117:10]
  assign _GEN_10028 = 5'h9 == _T_988 ? welem[9] : _GEN_10027; // @[Execute.scala 117:10]
  assign _GEN_10029 = 5'ha == _T_988 ? welem[10] : _GEN_10028; // @[Execute.scala 117:10]
  assign _GEN_10030 = 5'hb == _T_988 ? welem[11] : _GEN_10029; // @[Execute.scala 117:10]
  assign _GEN_10031 = 5'hc == _T_988 ? welem[12] : _GEN_10030; // @[Execute.scala 117:10]
  assign _GEN_10032 = 5'hd == _T_988 ? welem[13] : _GEN_10031; // @[Execute.scala 117:10]
  assign _GEN_10033 = 5'he == _T_988 ? welem[14] : _GEN_10032; // @[Execute.scala 117:10]
  assign _GEN_10034 = 5'hf == _T_988 ? welem[15] : _GEN_10033; // @[Execute.scala 117:10]
  assign _GEN_10035 = 5'h10 == _T_988 ? welem[16] : _GEN_10034; // @[Execute.scala 117:10]
  assign _GEN_10036 = 5'h11 == _T_988 ? welem[17] : _GEN_10035; // @[Execute.scala 117:10]
  assign _GEN_10037 = 5'h12 == _T_988 ? welem[18] : _GEN_10036; // @[Execute.scala 117:10]
  assign _GEN_10038 = 5'h13 == _T_988 ? welem[19] : _GEN_10037; // @[Execute.scala 117:10]
  assign _GEN_10039 = 5'h14 == _T_988 ? welem[20] : _GEN_10038; // @[Execute.scala 117:10]
  assign _GEN_10040 = 5'h15 == _T_988 ? welem[21] : _GEN_10039; // @[Execute.scala 117:10]
  assign _GEN_10041 = 5'h16 == _T_988 ? welem[22] : _GEN_10040; // @[Execute.scala 117:10]
  assign _GEN_10042 = 5'h17 == _T_988 ? welem[23] : _GEN_10041; // @[Execute.scala 117:10]
  assign _GEN_10043 = 5'h18 == _T_988 ? welem[24] : _GEN_10042; // @[Execute.scala 117:10]
  assign _GEN_10044 = 5'h19 == _T_988 ? welem[25] : _GEN_10043; // @[Execute.scala 117:10]
  assign _GEN_10045 = 5'h1a == _T_988 ? welem[26] : _GEN_10044; // @[Execute.scala 117:10]
  assign _GEN_10046 = 5'h1b == _T_988 ? welem[27] : _GEN_10045; // @[Execute.scala 117:10]
  assign _GEN_10047 = 5'h1c == _T_988 ? welem[28] : _GEN_10046; // @[Execute.scala 117:10]
  assign _GEN_10048 = 5'h1d == _T_988 ? welem[29] : _GEN_10047; // @[Execute.scala 117:10]
  assign _GEN_10049 = 5'h1e == _T_988 ? welem[30] : _GEN_10048; // @[Execute.scala 117:10]
  assign _GEN_10050 = 5'h1f == _T_988 ? welem[31] : _GEN_10049; // @[Execute.scala 117:10]
  assign _T_989 = _T_984 ? _GEN_10018 : _GEN_10050; // @[Execute.scala 117:10]
  assign _T_990 = r[4:0] < 5'h6; // @[Execute.scala 117:15]
  assign _T_992 = r[4:0] - 5'h6; // @[Execute.scala 117:37]
  assign _T_994 = 5'h1a + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_10052 = 5'h1 == _T_992 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10053 = 5'h2 == _T_992 ? welem[2] : _GEN_10052; // @[Execute.scala 117:10]
  assign _GEN_10054 = 5'h3 == _T_992 ? welem[3] : _GEN_10053; // @[Execute.scala 117:10]
  assign _GEN_10055 = 5'h4 == _T_992 ? welem[4] : _GEN_10054; // @[Execute.scala 117:10]
  assign _GEN_10056 = 5'h5 == _T_992 ? welem[5] : _GEN_10055; // @[Execute.scala 117:10]
  assign _GEN_10057 = 5'h6 == _T_992 ? welem[6] : _GEN_10056; // @[Execute.scala 117:10]
  assign _GEN_10058 = 5'h7 == _T_992 ? welem[7] : _GEN_10057; // @[Execute.scala 117:10]
  assign _GEN_10059 = 5'h8 == _T_992 ? welem[8] : _GEN_10058; // @[Execute.scala 117:10]
  assign _GEN_10060 = 5'h9 == _T_992 ? welem[9] : _GEN_10059; // @[Execute.scala 117:10]
  assign _GEN_10061 = 5'ha == _T_992 ? welem[10] : _GEN_10060; // @[Execute.scala 117:10]
  assign _GEN_10062 = 5'hb == _T_992 ? welem[11] : _GEN_10061; // @[Execute.scala 117:10]
  assign _GEN_10063 = 5'hc == _T_992 ? welem[12] : _GEN_10062; // @[Execute.scala 117:10]
  assign _GEN_10064 = 5'hd == _T_992 ? welem[13] : _GEN_10063; // @[Execute.scala 117:10]
  assign _GEN_10065 = 5'he == _T_992 ? welem[14] : _GEN_10064; // @[Execute.scala 117:10]
  assign _GEN_10066 = 5'hf == _T_992 ? welem[15] : _GEN_10065; // @[Execute.scala 117:10]
  assign _GEN_10067 = 5'h10 == _T_992 ? welem[16] : _GEN_10066; // @[Execute.scala 117:10]
  assign _GEN_10068 = 5'h11 == _T_992 ? welem[17] : _GEN_10067; // @[Execute.scala 117:10]
  assign _GEN_10069 = 5'h12 == _T_992 ? welem[18] : _GEN_10068; // @[Execute.scala 117:10]
  assign _GEN_10070 = 5'h13 == _T_992 ? welem[19] : _GEN_10069; // @[Execute.scala 117:10]
  assign _GEN_10071 = 5'h14 == _T_992 ? welem[20] : _GEN_10070; // @[Execute.scala 117:10]
  assign _GEN_10072 = 5'h15 == _T_992 ? welem[21] : _GEN_10071; // @[Execute.scala 117:10]
  assign _GEN_10073 = 5'h16 == _T_992 ? welem[22] : _GEN_10072; // @[Execute.scala 117:10]
  assign _GEN_10074 = 5'h17 == _T_992 ? welem[23] : _GEN_10073; // @[Execute.scala 117:10]
  assign _GEN_10075 = 5'h18 == _T_992 ? welem[24] : _GEN_10074; // @[Execute.scala 117:10]
  assign _GEN_10076 = 5'h19 == _T_992 ? welem[25] : _GEN_10075; // @[Execute.scala 117:10]
  assign _GEN_10077 = 5'h1a == _T_992 ? welem[26] : _GEN_10076; // @[Execute.scala 117:10]
  assign _GEN_10078 = 5'h1b == _T_992 ? welem[27] : _GEN_10077; // @[Execute.scala 117:10]
  assign _GEN_10079 = 5'h1c == _T_992 ? welem[28] : _GEN_10078; // @[Execute.scala 117:10]
  assign _GEN_10080 = 5'h1d == _T_992 ? welem[29] : _GEN_10079; // @[Execute.scala 117:10]
  assign _GEN_10081 = 5'h1e == _T_992 ? welem[30] : _GEN_10080; // @[Execute.scala 117:10]
  assign _GEN_10082 = 5'h1f == _T_992 ? welem[31] : _GEN_10081; // @[Execute.scala 117:10]
  assign _GEN_10084 = 5'h1 == _T_994 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10085 = 5'h2 == _T_994 ? welem[2] : _GEN_10084; // @[Execute.scala 117:10]
  assign _GEN_10086 = 5'h3 == _T_994 ? welem[3] : _GEN_10085; // @[Execute.scala 117:10]
  assign _GEN_10087 = 5'h4 == _T_994 ? welem[4] : _GEN_10086; // @[Execute.scala 117:10]
  assign _GEN_10088 = 5'h5 == _T_994 ? welem[5] : _GEN_10087; // @[Execute.scala 117:10]
  assign _GEN_10089 = 5'h6 == _T_994 ? welem[6] : _GEN_10088; // @[Execute.scala 117:10]
  assign _GEN_10090 = 5'h7 == _T_994 ? welem[7] : _GEN_10089; // @[Execute.scala 117:10]
  assign _GEN_10091 = 5'h8 == _T_994 ? welem[8] : _GEN_10090; // @[Execute.scala 117:10]
  assign _GEN_10092 = 5'h9 == _T_994 ? welem[9] : _GEN_10091; // @[Execute.scala 117:10]
  assign _GEN_10093 = 5'ha == _T_994 ? welem[10] : _GEN_10092; // @[Execute.scala 117:10]
  assign _GEN_10094 = 5'hb == _T_994 ? welem[11] : _GEN_10093; // @[Execute.scala 117:10]
  assign _GEN_10095 = 5'hc == _T_994 ? welem[12] : _GEN_10094; // @[Execute.scala 117:10]
  assign _GEN_10096 = 5'hd == _T_994 ? welem[13] : _GEN_10095; // @[Execute.scala 117:10]
  assign _GEN_10097 = 5'he == _T_994 ? welem[14] : _GEN_10096; // @[Execute.scala 117:10]
  assign _GEN_10098 = 5'hf == _T_994 ? welem[15] : _GEN_10097; // @[Execute.scala 117:10]
  assign _GEN_10099 = 5'h10 == _T_994 ? welem[16] : _GEN_10098; // @[Execute.scala 117:10]
  assign _GEN_10100 = 5'h11 == _T_994 ? welem[17] : _GEN_10099; // @[Execute.scala 117:10]
  assign _GEN_10101 = 5'h12 == _T_994 ? welem[18] : _GEN_10100; // @[Execute.scala 117:10]
  assign _GEN_10102 = 5'h13 == _T_994 ? welem[19] : _GEN_10101; // @[Execute.scala 117:10]
  assign _GEN_10103 = 5'h14 == _T_994 ? welem[20] : _GEN_10102; // @[Execute.scala 117:10]
  assign _GEN_10104 = 5'h15 == _T_994 ? welem[21] : _GEN_10103; // @[Execute.scala 117:10]
  assign _GEN_10105 = 5'h16 == _T_994 ? welem[22] : _GEN_10104; // @[Execute.scala 117:10]
  assign _GEN_10106 = 5'h17 == _T_994 ? welem[23] : _GEN_10105; // @[Execute.scala 117:10]
  assign _GEN_10107 = 5'h18 == _T_994 ? welem[24] : _GEN_10106; // @[Execute.scala 117:10]
  assign _GEN_10108 = 5'h19 == _T_994 ? welem[25] : _GEN_10107; // @[Execute.scala 117:10]
  assign _GEN_10109 = 5'h1a == _T_994 ? welem[26] : _GEN_10108; // @[Execute.scala 117:10]
  assign _GEN_10110 = 5'h1b == _T_994 ? welem[27] : _GEN_10109; // @[Execute.scala 117:10]
  assign _GEN_10111 = 5'h1c == _T_994 ? welem[28] : _GEN_10110; // @[Execute.scala 117:10]
  assign _GEN_10112 = 5'h1d == _T_994 ? welem[29] : _GEN_10111; // @[Execute.scala 117:10]
  assign _GEN_10113 = 5'h1e == _T_994 ? welem[30] : _GEN_10112; // @[Execute.scala 117:10]
  assign _GEN_10114 = 5'h1f == _T_994 ? welem[31] : _GEN_10113; // @[Execute.scala 117:10]
  assign _T_995 = _T_990 ? _GEN_10082 : _GEN_10114; // @[Execute.scala 117:10]
  assign _T_996 = r[4:0] < 5'h5; // @[Execute.scala 117:15]
  assign _T_998 = r[4:0] - 5'h5; // @[Execute.scala 117:37]
  assign _T_1000 = 5'h1b + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_10116 = 5'h1 == _T_998 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10117 = 5'h2 == _T_998 ? welem[2] : _GEN_10116; // @[Execute.scala 117:10]
  assign _GEN_10118 = 5'h3 == _T_998 ? welem[3] : _GEN_10117; // @[Execute.scala 117:10]
  assign _GEN_10119 = 5'h4 == _T_998 ? welem[4] : _GEN_10118; // @[Execute.scala 117:10]
  assign _GEN_10120 = 5'h5 == _T_998 ? welem[5] : _GEN_10119; // @[Execute.scala 117:10]
  assign _GEN_10121 = 5'h6 == _T_998 ? welem[6] : _GEN_10120; // @[Execute.scala 117:10]
  assign _GEN_10122 = 5'h7 == _T_998 ? welem[7] : _GEN_10121; // @[Execute.scala 117:10]
  assign _GEN_10123 = 5'h8 == _T_998 ? welem[8] : _GEN_10122; // @[Execute.scala 117:10]
  assign _GEN_10124 = 5'h9 == _T_998 ? welem[9] : _GEN_10123; // @[Execute.scala 117:10]
  assign _GEN_10125 = 5'ha == _T_998 ? welem[10] : _GEN_10124; // @[Execute.scala 117:10]
  assign _GEN_10126 = 5'hb == _T_998 ? welem[11] : _GEN_10125; // @[Execute.scala 117:10]
  assign _GEN_10127 = 5'hc == _T_998 ? welem[12] : _GEN_10126; // @[Execute.scala 117:10]
  assign _GEN_10128 = 5'hd == _T_998 ? welem[13] : _GEN_10127; // @[Execute.scala 117:10]
  assign _GEN_10129 = 5'he == _T_998 ? welem[14] : _GEN_10128; // @[Execute.scala 117:10]
  assign _GEN_10130 = 5'hf == _T_998 ? welem[15] : _GEN_10129; // @[Execute.scala 117:10]
  assign _GEN_10131 = 5'h10 == _T_998 ? welem[16] : _GEN_10130; // @[Execute.scala 117:10]
  assign _GEN_10132 = 5'h11 == _T_998 ? welem[17] : _GEN_10131; // @[Execute.scala 117:10]
  assign _GEN_10133 = 5'h12 == _T_998 ? welem[18] : _GEN_10132; // @[Execute.scala 117:10]
  assign _GEN_10134 = 5'h13 == _T_998 ? welem[19] : _GEN_10133; // @[Execute.scala 117:10]
  assign _GEN_10135 = 5'h14 == _T_998 ? welem[20] : _GEN_10134; // @[Execute.scala 117:10]
  assign _GEN_10136 = 5'h15 == _T_998 ? welem[21] : _GEN_10135; // @[Execute.scala 117:10]
  assign _GEN_10137 = 5'h16 == _T_998 ? welem[22] : _GEN_10136; // @[Execute.scala 117:10]
  assign _GEN_10138 = 5'h17 == _T_998 ? welem[23] : _GEN_10137; // @[Execute.scala 117:10]
  assign _GEN_10139 = 5'h18 == _T_998 ? welem[24] : _GEN_10138; // @[Execute.scala 117:10]
  assign _GEN_10140 = 5'h19 == _T_998 ? welem[25] : _GEN_10139; // @[Execute.scala 117:10]
  assign _GEN_10141 = 5'h1a == _T_998 ? welem[26] : _GEN_10140; // @[Execute.scala 117:10]
  assign _GEN_10142 = 5'h1b == _T_998 ? welem[27] : _GEN_10141; // @[Execute.scala 117:10]
  assign _GEN_10143 = 5'h1c == _T_998 ? welem[28] : _GEN_10142; // @[Execute.scala 117:10]
  assign _GEN_10144 = 5'h1d == _T_998 ? welem[29] : _GEN_10143; // @[Execute.scala 117:10]
  assign _GEN_10145 = 5'h1e == _T_998 ? welem[30] : _GEN_10144; // @[Execute.scala 117:10]
  assign _GEN_10146 = 5'h1f == _T_998 ? welem[31] : _GEN_10145; // @[Execute.scala 117:10]
  assign _GEN_10148 = 5'h1 == _T_1000 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10149 = 5'h2 == _T_1000 ? welem[2] : _GEN_10148; // @[Execute.scala 117:10]
  assign _GEN_10150 = 5'h3 == _T_1000 ? welem[3] : _GEN_10149; // @[Execute.scala 117:10]
  assign _GEN_10151 = 5'h4 == _T_1000 ? welem[4] : _GEN_10150; // @[Execute.scala 117:10]
  assign _GEN_10152 = 5'h5 == _T_1000 ? welem[5] : _GEN_10151; // @[Execute.scala 117:10]
  assign _GEN_10153 = 5'h6 == _T_1000 ? welem[6] : _GEN_10152; // @[Execute.scala 117:10]
  assign _GEN_10154 = 5'h7 == _T_1000 ? welem[7] : _GEN_10153; // @[Execute.scala 117:10]
  assign _GEN_10155 = 5'h8 == _T_1000 ? welem[8] : _GEN_10154; // @[Execute.scala 117:10]
  assign _GEN_10156 = 5'h9 == _T_1000 ? welem[9] : _GEN_10155; // @[Execute.scala 117:10]
  assign _GEN_10157 = 5'ha == _T_1000 ? welem[10] : _GEN_10156; // @[Execute.scala 117:10]
  assign _GEN_10158 = 5'hb == _T_1000 ? welem[11] : _GEN_10157; // @[Execute.scala 117:10]
  assign _GEN_10159 = 5'hc == _T_1000 ? welem[12] : _GEN_10158; // @[Execute.scala 117:10]
  assign _GEN_10160 = 5'hd == _T_1000 ? welem[13] : _GEN_10159; // @[Execute.scala 117:10]
  assign _GEN_10161 = 5'he == _T_1000 ? welem[14] : _GEN_10160; // @[Execute.scala 117:10]
  assign _GEN_10162 = 5'hf == _T_1000 ? welem[15] : _GEN_10161; // @[Execute.scala 117:10]
  assign _GEN_10163 = 5'h10 == _T_1000 ? welem[16] : _GEN_10162; // @[Execute.scala 117:10]
  assign _GEN_10164 = 5'h11 == _T_1000 ? welem[17] : _GEN_10163; // @[Execute.scala 117:10]
  assign _GEN_10165 = 5'h12 == _T_1000 ? welem[18] : _GEN_10164; // @[Execute.scala 117:10]
  assign _GEN_10166 = 5'h13 == _T_1000 ? welem[19] : _GEN_10165; // @[Execute.scala 117:10]
  assign _GEN_10167 = 5'h14 == _T_1000 ? welem[20] : _GEN_10166; // @[Execute.scala 117:10]
  assign _GEN_10168 = 5'h15 == _T_1000 ? welem[21] : _GEN_10167; // @[Execute.scala 117:10]
  assign _GEN_10169 = 5'h16 == _T_1000 ? welem[22] : _GEN_10168; // @[Execute.scala 117:10]
  assign _GEN_10170 = 5'h17 == _T_1000 ? welem[23] : _GEN_10169; // @[Execute.scala 117:10]
  assign _GEN_10171 = 5'h18 == _T_1000 ? welem[24] : _GEN_10170; // @[Execute.scala 117:10]
  assign _GEN_10172 = 5'h19 == _T_1000 ? welem[25] : _GEN_10171; // @[Execute.scala 117:10]
  assign _GEN_10173 = 5'h1a == _T_1000 ? welem[26] : _GEN_10172; // @[Execute.scala 117:10]
  assign _GEN_10174 = 5'h1b == _T_1000 ? welem[27] : _GEN_10173; // @[Execute.scala 117:10]
  assign _GEN_10175 = 5'h1c == _T_1000 ? welem[28] : _GEN_10174; // @[Execute.scala 117:10]
  assign _GEN_10176 = 5'h1d == _T_1000 ? welem[29] : _GEN_10175; // @[Execute.scala 117:10]
  assign _GEN_10177 = 5'h1e == _T_1000 ? welem[30] : _GEN_10176; // @[Execute.scala 117:10]
  assign _GEN_10178 = 5'h1f == _T_1000 ? welem[31] : _GEN_10177; // @[Execute.scala 117:10]
  assign _T_1001 = _T_996 ? _GEN_10146 : _GEN_10178; // @[Execute.scala 117:10]
  assign _T_1002 = r[4:0] < 5'h4; // @[Execute.scala 117:15]
  assign _T_1004 = r[4:0] - 5'h4; // @[Execute.scala 117:37]
  assign _T_1006 = 5'h1c + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_10180 = 5'h1 == _T_1004 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10181 = 5'h2 == _T_1004 ? welem[2] : _GEN_10180; // @[Execute.scala 117:10]
  assign _GEN_10182 = 5'h3 == _T_1004 ? welem[3] : _GEN_10181; // @[Execute.scala 117:10]
  assign _GEN_10183 = 5'h4 == _T_1004 ? welem[4] : _GEN_10182; // @[Execute.scala 117:10]
  assign _GEN_10184 = 5'h5 == _T_1004 ? welem[5] : _GEN_10183; // @[Execute.scala 117:10]
  assign _GEN_10185 = 5'h6 == _T_1004 ? welem[6] : _GEN_10184; // @[Execute.scala 117:10]
  assign _GEN_10186 = 5'h7 == _T_1004 ? welem[7] : _GEN_10185; // @[Execute.scala 117:10]
  assign _GEN_10187 = 5'h8 == _T_1004 ? welem[8] : _GEN_10186; // @[Execute.scala 117:10]
  assign _GEN_10188 = 5'h9 == _T_1004 ? welem[9] : _GEN_10187; // @[Execute.scala 117:10]
  assign _GEN_10189 = 5'ha == _T_1004 ? welem[10] : _GEN_10188; // @[Execute.scala 117:10]
  assign _GEN_10190 = 5'hb == _T_1004 ? welem[11] : _GEN_10189; // @[Execute.scala 117:10]
  assign _GEN_10191 = 5'hc == _T_1004 ? welem[12] : _GEN_10190; // @[Execute.scala 117:10]
  assign _GEN_10192 = 5'hd == _T_1004 ? welem[13] : _GEN_10191; // @[Execute.scala 117:10]
  assign _GEN_10193 = 5'he == _T_1004 ? welem[14] : _GEN_10192; // @[Execute.scala 117:10]
  assign _GEN_10194 = 5'hf == _T_1004 ? welem[15] : _GEN_10193; // @[Execute.scala 117:10]
  assign _GEN_10195 = 5'h10 == _T_1004 ? welem[16] : _GEN_10194; // @[Execute.scala 117:10]
  assign _GEN_10196 = 5'h11 == _T_1004 ? welem[17] : _GEN_10195; // @[Execute.scala 117:10]
  assign _GEN_10197 = 5'h12 == _T_1004 ? welem[18] : _GEN_10196; // @[Execute.scala 117:10]
  assign _GEN_10198 = 5'h13 == _T_1004 ? welem[19] : _GEN_10197; // @[Execute.scala 117:10]
  assign _GEN_10199 = 5'h14 == _T_1004 ? welem[20] : _GEN_10198; // @[Execute.scala 117:10]
  assign _GEN_10200 = 5'h15 == _T_1004 ? welem[21] : _GEN_10199; // @[Execute.scala 117:10]
  assign _GEN_10201 = 5'h16 == _T_1004 ? welem[22] : _GEN_10200; // @[Execute.scala 117:10]
  assign _GEN_10202 = 5'h17 == _T_1004 ? welem[23] : _GEN_10201; // @[Execute.scala 117:10]
  assign _GEN_10203 = 5'h18 == _T_1004 ? welem[24] : _GEN_10202; // @[Execute.scala 117:10]
  assign _GEN_10204 = 5'h19 == _T_1004 ? welem[25] : _GEN_10203; // @[Execute.scala 117:10]
  assign _GEN_10205 = 5'h1a == _T_1004 ? welem[26] : _GEN_10204; // @[Execute.scala 117:10]
  assign _GEN_10206 = 5'h1b == _T_1004 ? welem[27] : _GEN_10205; // @[Execute.scala 117:10]
  assign _GEN_10207 = 5'h1c == _T_1004 ? welem[28] : _GEN_10206; // @[Execute.scala 117:10]
  assign _GEN_10208 = 5'h1d == _T_1004 ? welem[29] : _GEN_10207; // @[Execute.scala 117:10]
  assign _GEN_10209 = 5'h1e == _T_1004 ? welem[30] : _GEN_10208; // @[Execute.scala 117:10]
  assign _GEN_10210 = 5'h1f == _T_1004 ? welem[31] : _GEN_10209; // @[Execute.scala 117:10]
  assign _GEN_10212 = 5'h1 == _T_1006 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10213 = 5'h2 == _T_1006 ? welem[2] : _GEN_10212; // @[Execute.scala 117:10]
  assign _GEN_10214 = 5'h3 == _T_1006 ? welem[3] : _GEN_10213; // @[Execute.scala 117:10]
  assign _GEN_10215 = 5'h4 == _T_1006 ? welem[4] : _GEN_10214; // @[Execute.scala 117:10]
  assign _GEN_10216 = 5'h5 == _T_1006 ? welem[5] : _GEN_10215; // @[Execute.scala 117:10]
  assign _GEN_10217 = 5'h6 == _T_1006 ? welem[6] : _GEN_10216; // @[Execute.scala 117:10]
  assign _GEN_10218 = 5'h7 == _T_1006 ? welem[7] : _GEN_10217; // @[Execute.scala 117:10]
  assign _GEN_10219 = 5'h8 == _T_1006 ? welem[8] : _GEN_10218; // @[Execute.scala 117:10]
  assign _GEN_10220 = 5'h9 == _T_1006 ? welem[9] : _GEN_10219; // @[Execute.scala 117:10]
  assign _GEN_10221 = 5'ha == _T_1006 ? welem[10] : _GEN_10220; // @[Execute.scala 117:10]
  assign _GEN_10222 = 5'hb == _T_1006 ? welem[11] : _GEN_10221; // @[Execute.scala 117:10]
  assign _GEN_10223 = 5'hc == _T_1006 ? welem[12] : _GEN_10222; // @[Execute.scala 117:10]
  assign _GEN_10224 = 5'hd == _T_1006 ? welem[13] : _GEN_10223; // @[Execute.scala 117:10]
  assign _GEN_10225 = 5'he == _T_1006 ? welem[14] : _GEN_10224; // @[Execute.scala 117:10]
  assign _GEN_10226 = 5'hf == _T_1006 ? welem[15] : _GEN_10225; // @[Execute.scala 117:10]
  assign _GEN_10227 = 5'h10 == _T_1006 ? welem[16] : _GEN_10226; // @[Execute.scala 117:10]
  assign _GEN_10228 = 5'h11 == _T_1006 ? welem[17] : _GEN_10227; // @[Execute.scala 117:10]
  assign _GEN_10229 = 5'h12 == _T_1006 ? welem[18] : _GEN_10228; // @[Execute.scala 117:10]
  assign _GEN_10230 = 5'h13 == _T_1006 ? welem[19] : _GEN_10229; // @[Execute.scala 117:10]
  assign _GEN_10231 = 5'h14 == _T_1006 ? welem[20] : _GEN_10230; // @[Execute.scala 117:10]
  assign _GEN_10232 = 5'h15 == _T_1006 ? welem[21] : _GEN_10231; // @[Execute.scala 117:10]
  assign _GEN_10233 = 5'h16 == _T_1006 ? welem[22] : _GEN_10232; // @[Execute.scala 117:10]
  assign _GEN_10234 = 5'h17 == _T_1006 ? welem[23] : _GEN_10233; // @[Execute.scala 117:10]
  assign _GEN_10235 = 5'h18 == _T_1006 ? welem[24] : _GEN_10234; // @[Execute.scala 117:10]
  assign _GEN_10236 = 5'h19 == _T_1006 ? welem[25] : _GEN_10235; // @[Execute.scala 117:10]
  assign _GEN_10237 = 5'h1a == _T_1006 ? welem[26] : _GEN_10236; // @[Execute.scala 117:10]
  assign _GEN_10238 = 5'h1b == _T_1006 ? welem[27] : _GEN_10237; // @[Execute.scala 117:10]
  assign _GEN_10239 = 5'h1c == _T_1006 ? welem[28] : _GEN_10238; // @[Execute.scala 117:10]
  assign _GEN_10240 = 5'h1d == _T_1006 ? welem[29] : _GEN_10239; // @[Execute.scala 117:10]
  assign _GEN_10241 = 5'h1e == _T_1006 ? welem[30] : _GEN_10240; // @[Execute.scala 117:10]
  assign _GEN_10242 = 5'h1f == _T_1006 ? welem[31] : _GEN_10241; // @[Execute.scala 117:10]
  assign _T_1007 = _T_1002 ? _GEN_10210 : _GEN_10242; // @[Execute.scala 117:10]
  assign _T_1008 = r[4:0] < 5'h3; // @[Execute.scala 117:15]
  assign _T_1010 = r[4:0] - 5'h3; // @[Execute.scala 117:37]
  assign _T_1012 = 5'h1d + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_10244 = 5'h1 == _T_1010 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10245 = 5'h2 == _T_1010 ? welem[2] : _GEN_10244; // @[Execute.scala 117:10]
  assign _GEN_10246 = 5'h3 == _T_1010 ? welem[3] : _GEN_10245; // @[Execute.scala 117:10]
  assign _GEN_10247 = 5'h4 == _T_1010 ? welem[4] : _GEN_10246; // @[Execute.scala 117:10]
  assign _GEN_10248 = 5'h5 == _T_1010 ? welem[5] : _GEN_10247; // @[Execute.scala 117:10]
  assign _GEN_10249 = 5'h6 == _T_1010 ? welem[6] : _GEN_10248; // @[Execute.scala 117:10]
  assign _GEN_10250 = 5'h7 == _T_1010 ? welem[7] : _GEN_10249; // @[Execute.scala 117:10]
  assign _GEN_10251 = 5'h8 == _T_1010 ? welem[8] : _GEN_10250; // @[Execute.scala 117:10]
  assign _GEN_10252 = 5'h9 == _T_1010 ? welem[9] : _GEN_10251; // @[Execute.scala 117:10]
  assign _GEN_10253 = 5'ha == _T_1010 ? welem[10] : _GEN_10252; // @[Execute.scala 117:10]
  assign _GEN_10254 = 5'hb == _T_1010 ? welem[11] : _GEN_10253; // @[Execute.scala 117:10]
  assign _GEN_10255 = 5'hc == _T_1010 ? welem[12] : _GEN_10254; // @[Execute.scala 117:10]
  assign _GEN_10256 = 5'hd == _T_1010 ? welem[13] : _GEN_10255; // @[Execute.scala 117:10]
  assign _GEN_10257 = 5'he == _T_1010 ? welem[14] : _GEN_10256; // @[Execute.scala 117:10]
  assign _GEN_10258 = 5'hf == _T_1010 ? welem[15] : _GEN_10257; // @[Execute.scala 117:10]
  assign _GEN_10259 = 5'h10 == _T_1010 ? welem[16] : _GEN_10258; // @[Execute.scala 117:10]
  assign _GEN_10260 = 5'h11 == _T_1010 ? welem[17] : _GEN_10259; // @[Execute.scala 117:10]
  assign _GEN_10261 = 5'h12 == _T_1010 ? welem[18] : _GEN_10260; // @[Execute.scala 117:10]
  assign _GEN_10262 = 5'h13 == _T_1010 ? welem[19] : _GEN_10261; // @[Execute.scala 117:10]
  assign _GEN_10263 = 5'h14 == _T_1010 ? welem[20] : _GEN_10262; // @[Execute.scala 117:10]
  assign _GEN_10264 = 5'h15 == _T_1010 ? welem[21] : _GEN_10263; // @[Execute.scala 117:10]
  assign _GEN_10265 = 5'h16 == _T_1010 ? welem[22] : _GEN_10264; // @[Execute.scala 117:10]
  assign _GEN_10266 = 5'h17 == _T_1010 ? welem[23] : _GEN_10265; // @[Execute.scala 117:10]
  assign _GEN_10267 = 5'h18 == _T_1010 ? welem[24] : _GEN_10266; // @[Execute.scala 117:10]
  assign _GEN_10268 = 5'h19 == _T_1010 ? welem[25] : _GEN_10267; // @[Execute.scala 117:10]
  assign _GEN_10269 = 5'h1a == _T_1010 ? welem[26] : _GEN_10268; // @[Execute.scala 117:10]
  assign _GEN_10270 = 5'h1b == _T_1010 ? welem[27] : _GEN_10269; // @[Execute.scala 117:10]
  assign _GEN_10271 = 5'h1c == _T_1010 ? welem[28] : _GEN_10270; // @[Execute.scala 117:10]
  assign _GEN_10272 = 5'h1d == _T_1010 ? welem[29] : _GEN_10271; // @[Execute.scala 117:10]
  assign _GEN_10273 = 5'h1e == _T_1010 ? welem[30] : _GEN_10272; // @[Execute.scala 117:10]
  assign _GEN_10274 = 5'h1f == _T_1010 ? welem[31] : _GEN_10273; // @[Execute.scala 117:10]
  assign _GEN_10276 = 5'h1 == _T_1012 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10277 = 5'h2 == _T_1012 ? welem[2] : _GEN_10276; // @[Execute.scala 117:10]
  assign _GEN_10278 = 5'h3 == _T_1012 ? welem[3] : _GEN_10277; // @[Execute.scala 117:10]
  assign _GEN_10279 = 5'h4 == _T_1012 ? welem[4] : _GEN_10278; // @[Execute.scala 117:10]
  assign _GEN_10280 = 5'h5 == _T_1012 ? welem[5] : _GEN_10279; // @[Execute.scala 117:10]
  assign _GEN_10281 = 5'h6 == _T_1012 ? welem[6] : _GEN_10280; // @[Execute.scala 117:10]
  assign _GEN_10282 = 5'h7 == _T_1012 ? welem[7] : _GEN_10281; // @[Execute.scala 117:10]
  assign _GEN_10283 = 5'h8 == _T_1012 ? welem[8] : _GEN_10282; // @[Execute.scala 117:10]
  assign _GEN_10284 = 5'h9 == _T_1012 ? welem[9] : _GEN_10283; // @[Execute.scala 117:10]
  assign _GEN_10285 = 5'ha == _T_1012 ? welem[10] : _GEN_10284; // @[Execute.scala 117:10]
  assign _GEN_10286 = 5'hb == _T_1012 ? welem[11] : _GEN_10285; // @[Execute.scala 117:10]
  assign _GEN_10287 = 5'hc == _T_1012 ? welem[12] : _GEN_10286; // @[Execute.scala 117:10]
  assign _GEN_10288 = 5'hd == _T_1012 ? welem[13] : _GEN_10287; // @[Execute.scala 117:10]
  assign _GEN_10289 = 5'he == _T_1012 ? welem[14] : _GEN_10288; // @[Execute.scala 117:10]
  assign _GEN_10290 = 5'hf == _T_1012 ? welem[15] : _GEN_10289; // @[Execute.scala 117:10]
  assign _GEN_10291 = 5'h10 == _T_1012 ? welem[16] : _GEN_10290; // @[Execute.scala 117:10]
  assign _GEN_10292 = 5'h11 == _T_1012 ? welem[17] : _GEN_10291; // @[Execute.scala 117:10]
  assign _GEN_10293 = 5'h12 == _T_1012 ? welem[18] : _GEN_10292; // @[Execute.scala 117:10]
  assign _GEN_10294 = 5'h13 == _T_1012 ? welem[19] : _GEN_10293; // @[Execute.scala 117:10]
  assign _GEN_10295 = 5'h14 == _T_1012 ? welem[20] : _GEN_10294; // @[Execute.scala 117:10]
  assign _GEN_10296 = 5'h15 == _T_1012 ? welem[21] : _GEN_10295; // @[Execute.scala 117:10]
  assign _GEN_10297 = 5'h16 == _T_1012 ? welem[22] : _GEN_10296; // @[Execute.scala 117:10]
  assign _GEN_10298 = 5'h17 == _T_1012 ? welem[23] : _GEN_10297; // @[Execute.scala 117:10]
  assign _GEN_10299 = 5'h18 == _T_1012 ? welem[24] : _GEN_10298; // @[Execute.scala 117:10]
  assign _GEN_10300 = 5'h19 == _T_1012 ? welem[25] : _GEN_10299; // @[Execute.scala 117:10]
  assign _GEN_10301 = 5'h1a == _T_1012 ? welem[26] : _GEN_10300; // @[Execute.scala 117:10]
  assign _GEN_10302 = 5'h1b == _T_1012 ? welem[27] : _GEN_10301; // @[Execute.scala 117:10]
  assign _GEN_10303 = 5'h1c == _T_1012 ? welem[28] : _GEN_10302; // @[Execute.scala 117:10]
  assign _GEN_10304 = 5'h1d == _T_1012 ? welem[29] : _GEN_10303; // @[Execute.scala 117:10]
  assign _GEN_10305 = 5'h1e == _T_1012 ? welem[30] : _GEN_10304; // @[Execute.scala 117:10]
  assign _GEN_10306 = 5'h1f == _T_1012 ? welem[31] : _GEN_10305; // @[Execute.scala 117:10]
  assign _T_1013 = _T_1008 ? _GEN_10274 : _GEN_10306; // @[Execute.scala 117:10]
  assign _T_1014 = r[4:0] < 5'h2; // @[Execute.scala 117:15]
  assign _T_1016 = r[4:0] - 5'h2; // @[Execute.scala 117:37]
  assign _T_1018 = 5'h1e + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_10308 = 5'h1 == _T_1016 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10309 = 5'h2 == _T_1016 ? welem[2] : _GEN_10308; // @[Execute.scala 117:10]
  assign _GEN_10310 = 5'h3 == _T_1016 ? welem[3] : _GEN_10309; // @[Execute.scala 117:10]
  assign _GEN_10311 = 5'h4 == _T_1016 ? welem[4] : _GEN_10310; // @[Execute.scala 117:10]
  assign _GEN_10312 = 5'h5 == _T_1016 ? welem[5] : _GEN_10311; // @[Execute.scala 117:10]
  assign _GEN_10313 = 5'h6 == _T_1016 ? welem[6] : _GEN_10312; // @[Execute.scala 117:10]
  assign _GEN_10314 = 5'h7 == _T_1016 ? welem[7] : _GEN_10313; // @[Execute.scala 117:10]
  assign _GEN_10315 = 5'h8 == _T_1016 ? welem[8] : _GEN_10314; // @[Execute.scala 117:10]
  assign _GEN_10316 = 5'h9 == _T_1016 ? welem[9] : _GEN_10315; // @[Execute.scala 117:10]
  assign _GEN_10317 = 5'ha == _T_1016 ? welem[10] : _GEN_10316; // @[Execute.scala 117:10]
  assign _GEN_10318 = 5'hb == _T_1016 ? welem[11] : _GEN_10317; // @[Execute.scala 117:10]
  assign _GEN_10319 = 5'hc == _T_1016 ? welem[12] : _GEN_10318; // @[Execute.scala 117:10]
  assign _GEN_10320 = 5'hd == _T_1016 ? welem[13] : _GEN_10319; // @[Execute.scala 117:10]
  assign _GEN_10321 = 5'he == _T_1016 ? welem[14] : _GEN_10320; // @[Execute.scala 117:10]
  assign _GEN_10322 = 5'hf == _T_1016 ? welem[15] : _GEN_10321; // @[Execute.scala 117:10]
  assign _GEN_10323 = 5'h10 == _T_1016 ? welem[16] : _GEN_10322; // @[Execute.scala 117:10]
  assign _GEN_10324 = 5'h11 == _T_1016 ? welem[17] : _GEN_10323; // @[Execute.scala 117:10]
  assign _GEN_10325 = 5'h12 == _T_1016 ? welem[18] : _GEN_10324; // @[Execute.scala 117:10]
  assign _GEN_10326 = 5'h13 == _T_1016 ? welem[19] : _GEN_10325; // @[Execute.scala 117:10]
  assign _GEN_10327 = 5'h14 == _T_1016 ? welem[20] : _GEN_10326; // @[Execute.scala 117:10]
  assign _GEN_10328 = 5'h15 == _T_1016 ? welem[21] : _GEN_10327; // @[Execute.scala 117:10]
  assign _GEN_10329 = 5'h16 == _T_1016 ? welem[22] : _GEN_10328; // @[Execute.scala 117:10]
  assign _GEN_10330 = 5'h17 == _T_1016 ? welem[23] : _GEN_10329; // @[Execute.scala 117:10]
  assign _GEN_10331 = 5'h18 == _T_1016 ? welem[24] : _GEN_10330; // @[Execute.scala 117:10]
  assign _GEN_10332 = 5'h19 == _T_1016 ? welem[25] : _GEN_10331; // @[Execute.scala 117:10]
  assign _GEN_10333 = 5'h1a == _T_1016 ? welem[26] : _GEN_10332; // @[Execute.scala 117:10]
  assign _GEN_10334 = 5'h1b == _T_1016 ? welem[27] : _GEN_10333; // @[Execute.scala 117:10]
  assign _GEN_10335 = 5'h1c == _T_1016 ? welem[28] : _GEN_10334; // @[Execute.scala 117:10]
  assign _GEN_10336 = 5'h1d == _T_1016 ? welem[29] : _GEN_10335; // @[Execute.scala 117:10]
  assign _GEN_10337 = 5'h1e == _T_1016 ? welem[30] : _GEN_10336; // @[Execute.scala 117:10]
  assign _GEN_10338 = 5'h1f == _T_1016 ? welem[31] : _GEN_10337; // @[Execute.scala 117:10]
  assign _GEN_10340 = 5'h1 == _T_1018 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10341 = 5'h2 == _T_1018 ? welem[2] : _GEN_10340; // @[Execute.scala 117:10]
  assign _GEN_10342 = 5'h3 == _T_1018 ? welem[3] : _GEN_10341; // @[Execute.scala 117:10]
  assign _GEN_10343 = 5'h4 == _T_1018 ? welem[4] : _GEN_10342; // @[Execute.scala 117:10]
  assign _GEN_10344 = 5'h5 == _T_1018 ? welem[5] : _GEN_10343; // @[Execute.scala 117:10]
  assign _GEN_10345 = 5'h6 == _T_1018 ? welem[6] : _GEN_10344; // @[Execute.scala 117:10]
  assign _GEN_10346 = 5'h7 == _T_1018 ? welem[7] : _GEN_10345; // @[Execute.scala 117:10]
  assign _GEN_10347 = 5'h8 == _T_1018 ? welem[8] : _GEN_10346; // @[Execute.scala 117:10]
  assign _GEN_10348 = 5'h9 == _T_1018 ? welem[9] : _GEN_10347; // @[Execute.scala 117:10]
  assign _GEN_10349 = 5'ha == _T_1018 ? welem[10] : _GEN_10348; // @[Execute.scala 117:10]
  assign _GEN_10350 = 5'hb == _T_1018 ? welem[11] : _GEN_10349; // @[Execute.scala 117:10]
  assign _GEN_10351 = 5'hc == _T_1018 ? welem[12] : _GEN_10350; // @[Execute.scala 117:10]
  assign _GEN_10352 = 5'hd == _T_1018 ? welem[13] : _GEN_10351; // @[Execute.scala 117:10]
  assign _GEN_10353 = 5'he == _T_1018 ? welem[14] : _GEN_10352; // @[Execute.scala 117:10]
  assign _GEN_10354 = 5'hf == _T_1018 ? welem[15] : _GEN_10353; // @[Execute.scala 117:10]
  assign _GEN_10355 = 5'h10 == _T_1018 ? welem[16] : _GEN_10354; // @[Execute.scala 117:10]
  assign _GEN_10356 = 5'h11 == _T_1018 ? welem[17] : _GEN_10355; // @[Execute.scala 117:10]
  assign _GEN_10357 = 5'h12 == _T_1018 ? welem[18] : _GEN_10356; // @[Execute.scala 117:10]
  assign _GEN_10358 = 5'h13 == _T_1018 ? welem[19] : _GEN_10357; // @[Execute.scala 117:10]
  assign _GEN_10359 = 5'h14 == _T_1018 ? welem[20] : _GEN_10358; // @[Execute.scala 117:10]
  assign _GEN_10360 = 5'h15 == _T_1018 ? welem[21] : _GEN_10359; // @[Execute.scala 117:10]
  assign _GEN_10361 = 5'h16 == _T_1018 ? welem[22] : _GEN_10360; // @[Execute.scala 117:10]
  assign _GEN_10362 = 5'h17 == _T_1018 ? welem[23] : _GEN_10361; // @[Execute.scala 117:10]
  assign _GEN_10363 = 5'h18 == _T_1018 ? welem[24] : _GEN_10362; // @[Execute.scala 117:10]
  assign _GEN_10364 = 5'h19 == _T_1018 ? welem[25] : _GEN_10363; // @[Execute.scala 117:10]
  assign _GEN_10365 = 5'h1a == _T_1018 ? welem[26] : _GEN_10364; // @[Execute.scala 117:10]
  assign _GEN_10366 = 5'h1b == _T_1018 ? welem[27] : _GEN_10365; // @[Execute.scala 117:10]
  assign _GEN_10367 = 5'h1c == _T_1018 ? welem[28] : _GEN_10366; // @[Execute.scala 117:10]
  assign _GEN_10368 = 5'h1d == _T_1018 ? welem[29] : _GEN_10367; // @[Execute.scala 117:10]
  assign _GEN_10369 = 5'h1e == _T_1018 ? welem[30] : _GEN_10368; // @[Execute.scala 117:10]
  assign _GEN_10370 = 5'h1f == _T_1018 ? welem[31] : _GEN_10369; // @[Execute.scala 117:10]
  assign _T_1019 = _T_1014 ? _GEN_10338 : _GEN_10370; // @[Execute.scala 117:10]
  assign _T_1020 = r[4:0] < 5'h1; // @[Execute.scala 117:15]
  assign _T_1022 = r[4:0] - 5'h1; // @[Execute.scala 117:37]
  assign _T_1024 = 5'h1f + r[4:0]; // @[Execute.scala 117:60]
  assign _GEN_10372 = 5'h1 == _T_1022 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10373 = 5'h2 == _T_1022 ? welem[2] : _GEN_10372; // @[Execute.scala 117:10]
  assign _GEN_10374 = 5'h3 == _T_1022 ? welem[3] : _GEN_10373; // @[Execute.scala 117:10]
  assign _GEN_10375 = 5'h4 == _T_1022 ? welem[4] : _GEN_10374; // @[Execute.scala 117:10]
  assign _GEN_10376 = 5'h5 == _T_1022 ? welem[5] : _GEN_10375; // @[Execute.scala 117:10]
  assign _GEN_10377 = 5'h6 == _T_1022 ? welem[6] : _GEN_10376; // @[Execute.scala 117:10]
  assign _GEN_10378 = 5'h7 == _T_1022 ? welem[7] : _GEN_10377; // @[Execute.scala 117:10]
  assign _GEN_10379 = 5'h8 == _T_1022 ? welem[8] : _GEN_10378; // @[Execute.scala 117:10]
  assign _GEN_10380 = 5'h9 == _T_1022 ? welem[9] : _GEN_10379; // @[Execute.scala 117:10]
  assign _GEN_10381 = 5'ha == _T_1022 ? welem[10] : _GEN_10380; // @[Execute.scala 117:10]
  assign _GEN_10382 = 5'hb == _T_1022 ? welem[11] : _GEN_10381; // @[Execute.scala 117:10]
  assign _GEN_10383 = 5'hc == _T_1022 ? welem[12] : _GEN_10382; // @[Execute.scala 117:10]
  assign _GEN_10384 = 5'hd == _T_1022 ? welem[13] : _GEN_10383; // @[Execute.scala 117:10]
  assign _GEN_10385 = 5'he == _T_1022 ? welem[14] : _GEN_10384; // @[Execute.scala 117:10]
  assign _GEN_10386 = 5'hf == _T_1022 ? welem[15] : _GEN_10385; // @[Execute.scala 117:10]
  assign _GEN_10387 = 5'h10 == _T_1022 ? welem[16] : _GEN_10386; // @[Execute.scala 117:10]
  assign _GEN_10388 = 5'h11 == _T_1022 ? welem[17] : _GEN_10387; // @[Execute.scala 117:10]
  assign _GEN_10389 = 5'h12 == _T_1022 ? welem[18] : _GEN_10388; // @[Execute.scala 117:10]
  assign _GEN_10390 = 5'h13 == _T_1022 ? welem[19] : _GEN_10389; // @[Execute.scala 117:10]
  assign _GEN_10391 = 5'h14 == _T_1022 ? welem[20] : _GEN_10390; // @[Execute.scala 117:10]
  assign _GEN_10392 = 5'h15 == _T_1022 ? welem[21] : _GEN_10391; // @[Execute.scala 117:10]
  assign _GEN_10393 = 5'h16 == _T_1022 ? welem[22] : _GEN_10392; // @[Execute.scala 117:10]
  assign _GEN_10394 = 5'h17 == _T_1022 ? welem[23] : _GEN_10393; // @[Execute.scala 117:10]
  assign _GEN_10395 = 5'h18 == _T_1022 ? welem[24] : _GEN_10394; // @[Execute.scala 117:10]
  assign _GEN_10396 = 5'h19 == _T_1022 ? welem[25] : _GEN_10395; // @[Execute.scala 117:10]
  assign _GEN_10397 = 5'h1a == _T_1022 ? welem[26] : _GEN_10396; // @[Execute.scala 117:10]
  assign _GEN_10398 = 5'h1b == _T_1022 ? welem[27] : _GEN_10397; // @[Execute.scala 117:10]
  assign _GEN_10399 = 5'h1c == _T_1022 ? welem[28] : _GEN_10398; // @[Execute.scala 117:10]
  assign _GEN_10400 = 5'h1d == _T_1022 ? welem[29] : _GEN_10399; // @[Execute.scala 117:10]
  assign _GEN_10401 = 5'h1e == _T_1022 ? welem[30] : _GEN_10400; // @[Execute.scala 117:10]
  assign _GEN_10402 = 5'h1f == _T_1022 ? welem[31] : _GEN_10401; // @[Execute.scala 117:10]
  assign _GEN_10404 = 5'h1 == _T_1024 ? welem[1] : welem[0]; // @[Execute.scala 117:10]
  assign _GEN_10405 = 5'h2 == _T_1024 ? welem[2] : _GEN_10404; // @[Execute.scala 117:10]
  assign _GEN_10406 = 5'h3 == _T_1024 ? welem[3] : _GEN_10405; // @[Execute.scala 117:10]
  assign _GEN_10407 = 5'h4 == _T_1024 ? welem[4] : _GEN_10406; // @[Execute.scala 117:10]
  assign _GEN_10408 = 5'h5 == _T_1024 ? welem[5] : _GEN_10407; // @[Execute.scala 117:10]
  assign _GEN_10409 = 5'h6 == _T_1024 ? welem[6] : _GEN_10408; // @[Execute.scala 117:10]
  assign _GEN_10410 = 5'h7 == _T_1024 ? welem[7] : _GEN_10409; // @[Execute.scala 117:10]
  assign _GEN_10411 = 5'h8 == _T_1024 ? welem[8] : _GEN_10410; // @[Execute.scala 117:10]
  assign _GEN_10412 = 5'h9 == _T_1024 ? welem[9] : _GEN_10411; // @[Execute.scala 117:10]
  assign _GEN_10413 = 5'ha == _T_1024 ? welem[10] : _GEN_10412; // @[Execute.scala 117:10]
  assign _GEN_10414 = 5'hb == _T_1024 ? welem[11] : _GEN_10413; // @[Execute.scala 117:10]
  assign _GEN_10415 = 5'hc == _T_1024 ? welem[12] : _GEN_10414; // @[Execute.scala 117:10]
  assign _GEN_10416 = 5'hd == _T_1024 ? welem[13] : _GEN_10415; // @[Execute.scala 117:10]
  assign _GEN_10417 = 5'he == _T_1024 ? welem[14] : _GEN_10416; // @[Execute.scala 117:10]
  assign _GEN_10418 = 5'hf == _T_1024 ? welem[15] : _GEN_10417; // @[Execute.scala 117:10]
  assign _GEN_10419 = 5'h10 == _T_1024 ? welem[16] : _GEN_10418; // @[Execute.scala 117:10]
  assign _GEN_10420 = 5'h11 == _T_1024 ? welem[17] : _GEN_10419; // @[Execute.scala 117:10]
  assign _GEN_10421 = 5'h12 == _T_1024 ? welem[18] : _GEN_10420; // @[Execute.scala 117:10]
  assign _GEN_10422 = 5'h13 == _T_1024 ? welem[19] : _GEN_10421; // @[Execute.scala 117:10]
  assign _GEN_10423 = 5'h14 == _T_1024 ? welem[20] : _GEN_10422; // @[Execute.scala 117:10]
  assign _GEN_10424 = 5'h15 == _T_1024 ? welem[21] : _GEN_10423; // @[Execute.scala 117:10]
  assign _GEN_10425 = 5'h16 == _T_1024 ? welem[22] : _GEN_10424; // @[Execute.scala 117:10]
  assign _GEN_10426 = 5'h17 == _T_1024 ? welem[23] : _GEN_10425; // @[Execute.scala 117:10]
  assign _GEN_10427 = 5'h18 == _T_1024 ? welem[24] : _GEN_10426; // @[Execute.scala 117:10]
  assign _GEN_10428 = 5'h19 == _T_1024 ? welem[25] : _GEN_10427; // @[Execute.scala 117:10]
  assign _GEN_10429 = 5'h1a == _T_1024 ? welem[26] : _GEN_10428; // @[Execute.scala 117:10]
  assign _GEN_10430 = 5'h1b == _T_1024 ? welem[27] : _GEN_10429; // @[Execute.scala 117:10]
  assign _GEN_10431 = 5'h1c == _T_1024 ? welem[28] : _GEN_10430; // @[Execute.scala 117:10]
  assign _GEN_10432 = 5'h1d == _T_1024 ? welem[29] : _GEN_10431; // @[Execute.scala 117:10]
  assign _GEN_10433 = 5'h1e == _T_1024 ? welem[30] : _GEN_10432; // @[Execute.scala 117:10]
  assign _GEN_10434 = 5'h1f == _T_1024 ? welem[31] : _GEN_10433; // @[Execute.scala 117:10]
  assign _T_1025 = _T_1020 ? _GEN_10402 : _GEN_10434; // @[Execute.scala 117:10]
  assign _T_1033 = {_T_881,_T_875,_T_869,_T_863,_T_857,_T_851,_T_845,_GEN_8418}; // @[Execute.scala 311:68]
  assign _T_1041 = {_T_929,_T_923,_T_917,_T_911,_T_905,_T_899,_T_893,_T_887,_T_1033}; // @[Execute.scala 311:68]
  assign _T_1048 = {_T_977,_T_971,_T_965,_T_959,_T_953,_T_947,_T_941,_T_935}; // @[Execute.scala 311:68]
  assign _T_1057 = {_T_1025,_T_1019,_T_1013,_T_1007,_T_1001,_T_995,_T_989,_T_983,_T_1048,_T_1041}; // @[Execute.scala 311:68]
  assign _T_1058 = {{32'd0}, _T_1057}; // @[Execute.scala 311:78]
  assign io_wmask = io_is32bit ? _T_1058 : _T_795; // @[Execute.scala 307:12]
  assign io_tmask = 7'h40 == onesD[6:0] ? 64'hffffffffffffffff : _GEN_8385; // @[Execute.scala 308:12]
endmodule
