// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

module cl_dma_pcis_slv #(parameter SCRB_MAX_ADDR = 64'h3FFFFFFFF, parameter SCRB_BURST_LEN_MINUS1 = 15, parameter NO_SCRB_INST = 1)

(
    input aclk,
    input aresetn,

    cfg_bus_t.master ddra_tst_cfg_bus,
    cfg_bus_t.master ddrb_tst_cfg_bus,
    cfg_bus_t.master ddrc_tst_cfg_bus,
    cfg_bus_t.master ddrd_tst_cfg_bus,

    scrb_bus_t.master ddra_scrb_bus,
    scrb_bus_t.master ddrb_scrb_bus,
    scrb_bus_t.master ddrc_scrb_bus,
    scrb_bus_t.master ddrd_scrb_bus,

    axi_bus_t.master cl_pcis_dram,
    axi_bus_t.master cl_rtl_m_axi,

    axi_bus_t.slave lcl_cl_sh_ddra,
    axi_bus_t.slave lcl_cl_sh_ddrb,
    axi_bus_t.slave lcl_cl_sh_ddrc,
    axi_bus_t.slave lcl_cl_sh_ddrd,

    axi_bus_t cl_pcis_dram_q
);
localparam NUM_CFG_STGS_CL_DDR_ATG = 4;
localparam NUM_CFG_STGS_SH_DDR_ATG = 4;

//----------------------------
// Internal signals
//----------------------------
axi_bus_t axi_m_00G_16G_();
axi_bus_t axi_m_32G_48G_();
axi_bus_t axi_m_16G_32G_();
axi_bus_t axi_m_48G_64G_();
// Register Slice
axi_bus_t axi_m_00G_16G_2();
axi_bus_t axi_m_16G_32G_2();
axi_bus_t axi_m_32G_48G_2();
axi_bus_t axi_m_48G_64G_2();
// Register Slice:
axi_bus_t axi_m_00G_16G_out();
axi_bus_t axi_m_16G_32G_out();
axi_bus_t axi_m_32G_48G_out();
axi_bus_t axi_m_48G_64G_out();

axi_bus_t sh_cl_pcis();

cfg_bus_t ddra_tst_cfg_bus_q();
cfg_bus_t ddrb_tst_cfg_bus_q();
cfg_bus_t ddrc_tst_cfg_bus_q();
cfg_bus_t ddrd_tst_cfg_bus_q();

scrb_bus_t ddra_scrb_bus_q();
scrb_bus_t ddrb_scrb_bus_q();
scrb_bus_t ddrc_scrb_bus_q();
scrb_bus_t ddrd_scrb_bus_q();

//----------------------------
// End Internal signals
//----------------------------


//reset synchronizers
(* dont_touch = "true" *) logic slr0_sync_aresetn;
(* dont_touch = "true" *) logic slr1_sync_aresetn;
(* dont_touch = "true" *) logic slr2_sync_aresetn;
lib_pipe #(.WIDTH(1), .STAGES(4)) SLR0_PIPE_RST_N (.clk(aclk), .rst_n(1'b1), .in_bus(aresetn), .out_bus(slr0_sync_aresetn));
lib_pipe #(.WIDTH(1), .STAGES(4)) SLR1_PIPE_RST_N (.clk(aclk), .rst_n(1'b1), .in_bus(aresetn), .out_bus(slr1_sync_aresetn));
lib_pipe #(.WIDTH(1), .STAGES(4)) SLR2_PIPE_RST_N (.clk(aclk), .rst_n(1'b1), .in_bus(aresetn), .out_bus(slr2_sync_aresetn));

//----------------------------
// flop the dma_pcis interface input of CL
//----------------------------

   // AXI4 Register Slice for dma_pcis interface
   axi_register_slice PCI_AXL_REG_SLC (
       .aclk          (aclk),
       .aresetn       (slr0_sync_aresetn),
       .s_axi_awid    (cl_pcis_dram.awid),
       .s_axi_awaddr  (cl_pcis_dram.awaddr),
       .s_axi_awlen   (cl_pcis_dram.awlen),
       .s_axi_awvalid (cl_pcis_dram.awvalid),
       .s_axi_awsize  (cl_pcis_dram.awsize),
       .s_axi_awready (cl_pcis_dram.awready),
       .s_axi_wdata   (cl_pcis_dram.wdata),
       .s_axi_wstrb   (cl_pcis_dram.wstrb),
       .s_axi_wlast   (cl_pcis_dram.wlast),
       .s_axi_wvalid  (cl_pcis_dram.wvalid),
       .s_axi_wready  (cl_pcis_dram.wready),
       .s_axi_bid     (cl_pcis_dram.bid),
       .s_axi_bresp   (cl_pcis_dram.bresp),
       .s_axi_bvalid  (cl_pcis_dram.bvalid),
       .s_axi_bready  (cl_pcis_dram.bready),
       .s_axi_arid    (cl_pcis_dram.arid),
       .s_axi_araddr  (cl_pcis_dram.araddr),
       .s_axi_arlen   (cl_pcis_dram.arlen),
       .s_axi_arvalid (cl_pcis_dram.arvalid),
       .s_axi_arsize  (cl_pcis_dram.arsize),
       .s_axi_arready (cl_pcis_dram.arready),
       .s_axi_rid     (cl_pcis_dram.rid),
       .s_axi_rdata   (cl_pcis_dram.rdata),
       .s_axi_rresp   (cl_pcis_dram.rresp),
       .s_axi_rlast   (cl_pcis_dram.rlast),
       .s_axi_rvalid  (cl_pcis_dram.rvalid),
       .s_axi_rready  (cl_pcis_dram.rready),

       .m_axi_awid    (cl_pcis_dram_q.awid),
       .m_axi_awaddr  (cl_pcis_dram_q.awaddr),
       .m_axi_awlen   (cl_pcis_dram_q.awlen),
       .m_axi_awvalid (cl_pcis_dram_q.awvalid),
       .m_axi_awsize  (cl_pcis_dram_q.awsize),
       .m_axi_awready (cl_pcis_dram_q.awready),
       .m_axi_wdata   (cl_pcis_dram_q.wdata),
       .m_axi_wstrb   (cl_pcis_dram_q.wstrb),
       .m_axi_wvalid  (cl_pcis_dram_q.wvalid),
       .m_axi_wlast   (cl_pcis_dram_q.wlast),
       .m_axi_wready  (cl_pcis_dram_q.wready),
       .m_axi_bresp   (cl_pcis_dram_q.bresp),
       .m_axi_bvalid  (cl_pcis_dram_q.bvalid),
       .m_axi_bid     (cl_pcis_dram_q.bid),
       .m_axi_bready  (cl_pcis_dram_q.bready),
       .m_axi_arid    (cl_pcis_dram_q.arid),
       .m_axi_araddr  (cl_pcis_dram_q.araddr),
       .m_axi_arlen   (cl_pcis_dram_q.arlen),
       .m_axi_arsize  (cl_pcis_dram_q.arsize),
       .m_axi_arvalid (cl_pcis_dram_q.arvalid),
       .m_axi_arready (cl_pcis_dram_q.arready),
       .m_axi_rid     (cl_pcis_dram_q.rid),
       .m_axi_rdata   (cl_pcis_dram_q.rdata),
       .m_axi_rresp   (cl_pcis_dram_q.rresp),
       .m_axi_rlast   (cl_pcis_dram_q.rlast),
       .m_axi_rvalid  (cl_pcis_dram_q.rvalid),
       .m_axi_rready  (cl_pcis_dram_q.rready)
   );

//-----------------------------------------------------
//TIE-OFF unused signals to prevent critical warnings
//-----------------------------------------------------
   assign cl_pcis_dram_q.rid[15:6] = 10'b0 ;
   assign cl_pcis_dram_q.bid[15:6] = 10'b0 ;

//----------------------------
// axi interconnect for DDR address decodes
//----------------------------
(* dont_touch = "true" *) cl_axi_interconnect AXI_CROSSBAR
       (.ACLK(aclk),
        .ARESETN(slr1_sync_aresetn),

        .M00_AXI_araddr    (axi_m_00G_16G_0.araddr),
        .M00_AXI_arburst   (),
        .M00_AXI_arcache   (),
        .M00_AXI_arid      (axi_m_00G_16G_0.arid[6:0]),
        .M00_AXI_arlen     (axi_m_00G_16G_0.arlen),
        .M00_AXI_arlock    (),
        .M00_AXI_arprot    (),
        .M00_AXI_arqos     (),
        .M00_AXI_arready   (axi_m_00G_16G_0.arready),
        .M00_AXI_arregion  (),
        .M00_AXI_arsize    (axi_m_00G_16G_0.arsize),
        .M00_AXI_arvalid   (axi_m_00G_16G_0.arvalid),
        .M00_AXI_awaddr    (axi_m_00G_16G_0.awaddr),
        .M00_AXI_awburst   (),
        .M00_AXI_awcache   (),
        .M00_AXI_awid      (axi_m_00G_16G_0.awid[6:0]),
        .M00_AXI_awlen     (axi_m_00G_16G_0.awlen),
        .M00_AXI_awlock    (),
        .M00_AXI_awprot    (),
        .M00_AXI_awqos     (),
        .M00_AXI_awready   (axi_m_00G_16G_0.awready),
        .M00_AXI_awregion  (),
        .M00_AXI_awsize    (axi_m_00G_16G_0.awsize),
        .M00_AXI_awvalid   (axi_m_00G_16G_0.awvalid),
        .M00_AXI_bid       (axi_m_00G_16G_0.bid[6:0]),
        .M00_AXI_bready    (axi_m_00G_16G_0.bready),
        .M00_AXI_bresp     (axi_m_00G_16G_0.bresp),
        .M00_AXI_bvalid    (axi_m_00G_16G_0.bvalid),
        .M00_AXI_rdata     (axi_m_00G_16G_0.rdata),
        .M00_AXI_rid       (axi_m_00G_16G_0.rid[6:0]),
        .M00_AXI_rlast     (axi_m_00G_16G_0.rlast),
        .M00_AXI_rready    (axi_m_00G_16G_0.rready),
        .M00_AXI_rresp     (axi_m_00G_16G_0.rresp),
        .M00_AXI_rvalid    (axi_m_00G_16G_0.rvalid),
        .M00_AXI_wdata     (axi_m_00G_16G_0.wdata),
        .M00_AXI_wlast     (axi_m_00G_16G_0.wlast),
        .M00_AXI_wready    (axi_m_00G_16G_0.wready),
        .M00_AXI_wstrb     (axi_m_00G_16G_0.wstrb),
        .M00_AXI_wvalid    (axi_m_00G_16G_0.wvalid),

        .M01_AXI_araddr    (axi_m_16G_32G_0.araddr),
        .M01_AXI_arburst   (),
        .M01_AXI_arcache   (),
        .M01_AXI_arid      (axi_m_16G_32G_0.arid[6:0]),
        .M01_AXI_arlen     (axi_m_16G_32G_0.arlen),
        .M01_AXI_arlock    (),
        .M01_AXI_arprot    (),
        .M01_AXI_arqos     (),
        .M01_AXI_arready   (axi_m_16G_32G_0.arready),
        .M01_AXI_arregion  (),
        .M01_AXI_arsize    (axi_m_16G_32G_0.arsize),
        .M01_AXI_arvalid   (axi_m_16G_32G_0.arvalid),
        .M01_AXI_awaddr    (axi_m_16G_32G_0.awaddr),
        .M01_AXI_awburst   (),
        .M01_AXI_awcache   (),
        .M01_AXI_awid      (axi_m_16G_32G_0.awid[6:0]),
        .M01_AXI_awlen     (axi_m_16G_32G_0.awlen),
        .M01_AXI_awlock    (),
        .M01_AXI_awprot    (),
        .M01_AXI_awqos     (),
        .M01_AXI_awready   (axi_m_16G_32G_0.awready),
        .M01_AXI_awregion  (),
        .M01_AXI_awsize    (axi_m_16G_32G_0.awsize),
        .M01_AXI_awvalid   (axi_m_16G_32G_0.awvalid),
        .M01_AXI_bid       (axi_m_16G_32G_0.bid[6:0]),
        .M01_AXI_bready    (axi_m_16G_32G_0.bready),
        .M01_AXI_bresp     (axi_m_16G_32G_0.bresp),
        .M01_AXI_bvalid    (axi_m_16G_32G_0.bvalid),
        .M01_AXI_rdata     (axi_m_16G_32G_0.rdata),
        .M01_AXI_rid       (axi_m_16G_32G_0.rid[6:0]),
        .M01_AXI_rlast     (axi_m_16G_32G_0.rlast),
        .M01_AXI_rready    (axi_m_16G_32G_0.rready),
        .M01_AXI_rresp     (axi_m_16G_32G_0.rresp),
        .M01_AXI_rvalid    (axi_m_16G_32G_0.rvalid),
        .M01_AXI_wdata     (axi_m_16G_32G_0.wdata),
        .M01_AXI_wlast     (axi_m_16G_32G_0.wlast),
        .M01_AXI_wready    (axi_m_16G_32G_0.wready),
        .M01_AXI_wstrb     (axi_m_16G_32G_0.wstrb),
        .M01_AXI_wvalid    (axi_m_16G_32G_0.wvalid),


        .M02_AXI_araddr    (axi_m_32G_48G_0.araddr),
        .M02_AXI_arburst   (),
        .M02_AXI_arcache   (),
        .M02_AXI_arid      (axi_m_32G_48G_0.arid[6:0]),
        .M02_AXI_arlen     (axi_m_32G_48G_0.arlen),
        .M02_AXI_arlock    (),
        .M02_AXI_arprot    (),
        .M02_AXI_arqos     (),
        .M02_AXI_arready   (axi_m_32G_48G_0.arready),
        .M02_AXI_arregion  (),
        .M02_AXI_arsize    (axi_m_32G_48G_0.arsize),
        .M02_AXI_arvalid   (axi_m_32G_48G_0.arvalid),
        .M02_AXI_awaddr    (axi_m_32G_48G_0.awaddr),
        .M02_AXI_awburst   (),
        .M02_AXI_awcache   (),
        .M02_AXI_awid      (axi_m_32G_48G_0.awid[6:0]),
        .M02_AXI_awlen     (axi_m_32G_48G_0.awlen),
        .M02_AXI_awlock    (),
        .M02_AXI_awprot    (),
        .M02_AXI_awqos     (),
        .M02_AXI_awready   (axi_m_32G_48G_0.awready),
        .M02_AXI_awregion  (),
        .M02_AXI_awsize    (axi_m_32G_48G_0.awsize),
        .M02_AXI_awvalid   (axi_m_32G_48G_0.awvalid),
        .M02_AXI_bid       (axi_m_32G_48G_0.bid[6:0]),
        .M02_AXI_bready    (axi_m_32G_48G_0.bready),
        .M02_AXI_bresp     (axi_m_32G_48G_0.bresp),
        .M02_AXI_bvalid    (axi_m_32G_48G_0.bvalid),
        .M02_AXI_rdata     (axi_m_32G_48G_0.rdata),
        .M02_AXI_rid       (axi_m_32G_48G_0.rid[6:0]),
        .M02_AXI_rlast     (axi_m_32G_48G_0.rlast),
        .M02_AXI_rready    (axi_m_32G_48G_0.rready),
        .M02_AXI_rresp     (axi_m_32G_48G_0.rresp),
        .M02_AXI_rvalid    (axi_m_32G_48G_0.rvalid),
        .M02_AXI_wdata     (axi_m_32G_48G_0.wdata),
        .M02_AXI_wlast     (axi_m_32G_48G_0.wlast),
        .M02_AXI_wready    (axi_m_32G_48G_0.wready),
        .M02_AXI_wstrb     (axi_m_32G_48G_0.wstrb),
        .M02_AXI_wvalid    (axi_m_32G_48G_0.wvalid),

        .M03_AXI_araddr    (axi_m_48G_64G_0.araddr),
        .M03_AXI_arburst   (),
        .M03_AXI_arcache   (),
        .M03_AXI_arid      (axi_m_48G_64G_0.arid[6:0]),
        .M03_AXI_arlen     (axi_m_48G_64G_0.arlen),
        .M03_AXI_arlock    (),
        .M03_AXI_arprot    (),
        .M03_AXI_arqos     (),
        .M03_AXI_arready   (axi_m_48G_64G_0.arready),
        .M03_AXI_arregion  (),
        .M03_AXI_arsize    (axi_m_48G_64G_0.arsize),
        .M03_AXI_arvalid   (axi_m_48G_64G_0.arvalid),
        .M03_AXI_awaddr    (axi_m_48G_64G_0.awaddr),
        .M03_AXI_awburst   (),
        .M03_AXI_awcache   (),
        .M03_AXI_awid      (axi_m_48G_64G_0.awid[6:0]),
        .M03_AXI_awlen     (axi_m_48G_64G_0.awlen),
        .M03_AXI_awlock    (),
        .M03_AXI_awprot    (),
        .M03_AXI_awqos     (),
        .M03_AXI_awready   (axi_m_48G_64G_0.awready),
        .M03_AXI_awregion  (),
        .M03_AXI_awsize    (axi_m_48G_64G_0.awsize),
        .M03_AXI_awvalid   (axi_m_48G_64G_0.awvalid),
        .M03_AXI_bid       (axi_m_48G_64G_0.bid[6:0]),
        .M03_AXI_bready    (axi_m_48G_64G_0.bready),
        .M03_AXI_bresp     (axi_m_48G_64G_0.bresp),
        .M03_AXI_bvalid    (axi_m_48G_64G_0.bvalid),
        .M03_AXI_rdata     (axi_m_48G_64G_0.rdata),
        .M03_AXI_rid       (axi_m_48G_64G_0.rid[6:0]),
        .M03_AXI_rlast     (axi_m_48G_64G_0.rlast),
        .M03_AXI_rready    (axi_m_48G_64G_0.rready),
        .M03_AXI_rresp     (axi_m_48G_64G_0.rresp),
        .M03_AXI_rvalid    (axi_m_48G_64G_0.rvalid),
        .M03_AXI_wdata     (axi_m_48G_64G_0.wdata),
        .M03_AXI_wlast     (axi_m_48G_64G_0.wlast),
        .M03_AXI_wready    (axi_m_48G_64G_0.wready),
        .M03_AXI_wstrb     (axi_m_48G_64G_0.wstrb),
        .M03_AXI_wvalid    (axi_m_48G_64G_0.wvalid),



        .S00_AXI_araddr    ({cl_pcis_dram_q.araddr[63:37], 1'b0, cl_pcis_dram_q.araddr[35:0]}),
        .S00_AXI_arburst   (2'b1),
        .S00_AXI_arcache   (4'b11),
        .S00_AXI_arid      (cl_pcis_dram_q.arid[5:0]),
        .S00_AXI_arlen     (cl_pcis_dram_q.arlen),
        .S00_AXI_arlock    (1'b0),
        .S00_AXI_arprot    (3'b10),
        .S00_AXI_arqos     (4'b0),
        .S00_AXI_arready   (cl_pcis_dram_q.arready),
        .S00_AXI_arregion  (4'b0),
        .S00_AXI_arsize    (cl_pcis_dram_q.arsize),
        .S00_AXI_arvalid   (cl_pcis_dram_q.arvalid),
        .S00_AXI_awaddr    ({cl_pcis_dram_q.awaddr[63:37], 1'b0, cl_pcis_dram_q.awaddr[35:0]}),
        .S00_AXI_awburst   (2'b1),
        .S00_AXI_awcache   (4'b11),
        .S00_AXI_awid      (cl_pcis_dram_q.awid[5:0]),
        .S00_AXI_awlen     (cl_pcis_dram_q.awlen),
        .S00_AXI_awlock    (1'b0),
        .S00_AXI_awprot    (3'b10),
        .S00_AXI_awqos     (4'b0),
        .S00_AXI_awready   (cl_pcis_dram_q.awready),
        .S00_AXI_awregion  (4'b0),
        .S00_AXI_awsize    (cl_pcis_dram_q.awsize),
        .S00_AXI_awvalid   (cl_pcis_dram_q.awvalid),
        .S00_AXI_bid       (cl_pcis_dram_q.bid[5:0]),
        .S00_AXI_bready    (cl_pcis_dram_q.bready),
        .S00_AXI_bresp     (cl_pcis_dram_q.bresp),
        .S00_AXI_bvalid    (cl_pcis_dram_q.bvalid),
        .S00_AXI_rdata     (cl_pcis_dram_q.rdata),
        .S00_AXI_rid       (cl_pcis_dram_q.rid[5:0]),
        .S00_AXI_rlast     (cl_pcis_dram_q.rlast),
        .S00_AXI_rready    (cl_pcis_dram_q.rready),
        .S00_AXI_rresp     (cl_pcis_dram_q.rresp),
        .S00_AXI_rvalid    (cl_pcis_dram_q.rvalid),
        .S00_AXI_wdata     (cl_pcis_dram_q.wdata),
        .S00_AXI_wlast     (cl_pcis_dram_q.wlast),
        .S00_AXI_wready    (cl_pcis_dram_q.wready),
        .S00_AXI_wstrb     (cl_pcis_dram_q.wstrb),
        .S00_AXI_wvalid    (cl_pcis_dram_q.wvalid),

        .S01_AXI_araddr    ({cl_rtl_m_axi.araddr[63:37], 1'b0, cl_rtl_m_axi.araddr[35:0]}),
        .S01_AXI_arburst   (2'b1),
        .S01_AXI_arcache   (4'b11),
        .S01_AXI_arid      (cl_rtl_m_axi.arid[5:0]),
        .S01_AXI_arlen     (cl_rtl_m_axi.arlen),
        .S01_AXI_arlock    (1'b0),
        .S01_AXI_arprot    (3'b10),
        .S01_AXI_arqos     (4'b0),
        .S01_AXI_arready   (cl_rtl_m_axi.arready),
        .S01_AXI_arregion  (4'b0),
        .S01_AXI_arsize    (cl_rtl_m_axi.arsize),
        .S01_AXI_arvalid   (cl_rtl_m_axi.arvalid),
        .S01_AXI_awaddr    ({cl_rtl_m_axi.awaddr[63:37], 1'b0, cl_rtl_m_axi.awaddr[35:0]}),
        .S01_AXI_awburst   (2'b1),
        .S01_AXI_awcache   (4'b11),
        .S01_AXI_awid      (cl_rtl_m_axi.awid[5:0]),
        .S01_AXI_awlen     (cl_rtl_m_axi.awlen),
        .S01_AXI_awlock    (1'b0),
        .S01_AXI_awprot    (3'b10),
        .S01_AXI_awqos     (4'b0),
        .S01_AXI_awready   (cl_rtl_m_axi.awready),
        .S01_AXI_awregion  (4'b0),
        .S01_AXI_awsize    (cl_rtl_m_axi.awsize),
        .S01_AXI_awvalid   (cl_rtl_m_axi.awvalid),
        .S01_AXI_bid       (cl_rtl_m_axi.bid[5:0]),
        .S01_AXI_bready    (cl_rtl_m_axi.bready),
        .S01_AXI_bresp     (cl_rtl_m_axi.bresp),
        .S01_AXI_bvalid    (cl_rtl_m_axi.bvalid),
        .S01_AXI_rdata     (cl_rtl_m_axi.rdata),
        .S01_AXI_rid       (cl_rtl_m_axi.rid[5:0]),
        .S01_AXI_rlast     (cl_rtl_m_axi.rlast),
        .S01_AXI_rready    (cl_rtl_m_axi.rready),
        .S01_AXI_rresp     (cl_rtl_m_axi.rresp),
        .S01_AXI_rvalid    (cl_rtl_m_axi.rvalid),
        .S01_AXI_wdata     (cl_rtl_m_axi.wdata),
        .S01_AXI_wlast     (cl_rtl_m_axi.wlast),
        .S01_AXI_wready    (cl_rtl_m_axi.wready),
        .S01_AXI_wstrb     (cl_rtl_m_axi.wstrb),
        .S01_AXI_wvalid    (cl_rtl_m_axi.wvalid));

//----------------------------
//                    flop the output of interconnect for 00G-16G
// back to back for SLR crossing
//----------------------------
   //back to back register slices for SLR crossing
   src_register_slice AXI4_REG_SLC_00G_16G_1 (
       .aclk           (aclk),
       .aresetn        (slr1_sync_aresetn),
       .s_axi_awid     (axi_m_00G_16G_0.awid),
       .s_axi_awaddr   ({axi_m_00G_16G_0.awaddr[63:36], 2'b0, axi_m_00G_16G_0.awaddr[33:0]}),
       .s_axi_awlen    (axi_m_00G_16G_0.awlen),
       .s_axi_awsize   (axi_m_00G_16G_0.awsize),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (axi_m_00G_16G_0.awvalid),
       .s_axi_awready  (axi_m_00G_16G_0.awready),
       .s_axi_wdata    (axi_m_00G_16G_0.wdata),
       .s_axi_wstrb    (axi_m_00G_16G_0.wstrb),
       .s_axi_wlast    (axi_m_00G_16G_0.wlast),
       .s_axi_wvalid   (axi_m_00G_16G_0.wvalid),
       .s_axi_wready   (axi_m_00G_16G_0.wready),
       .s_axi_bid      (axi_m_00G_16G_0.bid),
       .s_axi_bresp    (axi_m_00G_16G_0.bresp),
       .s_axi_bvalid   (axi_m_00G_16G_0.bvalid),
       .s_axi_bready   (axi_m_00G_16G_0.bready),
       .s_axi_arid     (axi_m_00G_16G_0.arid),
       .s_axi_araddr   ({axi_m_00G_16G_0.araddr[63:36], 2'b0, axi_m_00G_16G_0.araddr[33:0]}),
       .s_axi_arlen    (axi_m_00G_16G_0.arlen),
       .s_axi_arsize   (axi_m_00G_16G_0.arsize),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (axi_m_00G_16G_0.arvalid),
       .s_axi_arready  (axi_m_00G_16G_0.arready),
       .s_axi_rid      (axi_m_00G_16G_0.rid),
       .s_axi_rdata    (axi_m_00G_16G_0.rdata),
       .s_axi_rresp    (axi_m_00G_16G_0.rresp),
       .s_axi_rlast    (axi_m_00G_16G_0.rlast),
       .s_axi_rvalid   (axi_m_00G_16G_0.rvalid),
       .s_axi_rready   (axi_m_00G_16G_0.rready),
       .m_axi_awid     (axi_m_00G_16G_0.awid),
       .m_axi_awaddr   (axi_m_00G_16G_2.awaddr),
       .m_axi_awlen    (axi_m_00G_16G_2.awlen),
       .m_axi_awsize   (axi_m_00G_16G_2.awsize),
       .m_axi_awburst  (),
       .m_axi_awlock   (),
       .m_axi_awcache  (),
       .m_axi_awprot   (),
       .m_axi_awregion (),
       .m_axi_awqos    (),
       .m_axi_awvalid  (axi_m_00G_16G_2.awvalid),
       .m_axi_awready  (axi_m_00G_16G_2.awready),
       .m_axi_wdata    (axi_m_00G_16G_2.wdata),
       .m_axi_wstrb    (axi_m_00G_16G_2.wstrb),
       .m_axi_wlast    (axi_m_00G_16G_2.wlast),
       .m_axi_wvalid   (axi_m_00G_16G_2.wvalid),
       .m_axi_wready   (axi_m_00G_16G_2.wready),
       .m_axi_bid      (axi_m_00G_16G_2.bid),
       .m_axi_bresp    (axi_m_00G_16G_2.bresp),
       .m_axi_bvalid   (axi_m_00G_16G_2.bvalid),
       .m_axi_bready   (axi_m_00G_16G_2.bready),
       .m_axi_arid     (axi_m_00G_16G_2.arid),
       .m_axi_araddr   (axi_m_00G_16G_2.araddr),
       .m_axi_arlen    (axi_m_00G_16G_2.arlen),
       .m_axi_arsize   (axi_m_00G_16G_2.arsize),
       .m_axi_arburst  (),
       .m_axi_arlock   (),
       .m_axi_arcache  (),
       .m_axi_arprot   (),
       .m_axi_arregion (),
       .m_axi_arqos    (),
       .m_axi_arvalid  (axi_m_00G_16G_2.arvalid),
       .m_axi_arready  (axi_m_00G_16G_2.arready),
       .m_axi_rid      (axi_m_00G_16G_2.rid),
       .m_axi_rdata    (axi_m_00G_16G_2.rdata),
       .m_axi_rresp    (axi_m_00G_16G_2.rresp),
       .m_axi_rlast    (axi_m_00G_16G_2.rlast),
       .m_axi_rvalid   (axi_m_00G_16G_2.rvalid),
       .m_axi_rready   (axi_m_00G_16G_2.rready)
       );
   dest_register_slice AXI4_REG_SLC_00G_16G_2 (
       .aclk           (aclk),
       .aresetn        (slr2_sync_aresetn),
       .s_axi_awid     (axi_m_00G_16G_2.awid),
       .s_axi_awaddr   (axi_m_00G_16G_2.awaddr),
       .s_axi_awlen    (axi_m_00G_16G_2.awlen),
       .s_axi_awsize   (axi_m_00G_16G_2.awsize),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (axi_m_00G_16G_2.awvalid),
       .s_axi_awready  (axi_m_00G_16G_2.awready),
       .s_axi_wdata    (axi_m_00G_16G_2.wdata),
       .s_axi_wstrb    (axi_m_00G_16G_2.wstrb),
       .s_axi_wlast    (axi_m_00G_16G_2.wlast),
       .s_axi_wvalid   (axi_m_00G_16G_2.wvalid),
       .s_axi_wready   (axi_m_00G_16G_2.wready),
       .s_axi_bid      (axi_m_00G_16G_2.bid),
       .s_axi_bresp    (axi_m_00G_16G_2.bresp),
       .s_axi_bvalid   (axi_m_00G_16G_2.bvalid),
       .s_axi_bready   (axi_m_00G_16G_2.bready),
       .s_axi_arid     (axi_m_00G_16G_2.arid),
       .s_axi_araddr   (axi_m_00G_16G_2.araddr),
       .s_axi_arlen    (axi_m_00G_16G_2.arlen),
       .s_axi_arsize   (axi_m_00G_16G_2.arsize),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (axi_m_00G_16G_2.arvalid),
       .s_axi_arready  (axi_m_00G_16G_2.arready),
       .s_axi_rid      (axi_m_00G_16G_2.rid),
       .s_axi_rdata    (axi_m_00G_16G_2.rdata),
       .s_axi_rresp    (axi_m_00G_16G_2.rresp),
       .s_axi_rlast    (axi_m_00G_16G_2.rlast),
       .s_axi_rvalid   (axi_m_00G_16G_2.rvalid),
       .s_axi_rready   (axi_m_00G_16G_2.rready),
       .m_axi_awid     (axi_m_00G_16G_out.awid),
       .m_axi_awaddr   (axi_m_00G_16G_out.awaddr),
       .m_axi_awlen    (axi_m_00G_16G_out.awlen),
       .m_axi_awsize   (axi_m_00G_16G_out.awsize),
       .m_axi_awburst  (),
       .m_axi_awlock   (),
       .m_axi_awcache  (),
       .m_axi_awprot   (),
       .m_axi_awregion (),
       .m_axi_awqos    (),
       .m_axi_awvalid  (axi_m_00G_16G_out.awvalid),
       .m_axi_awready  (axi_m_00G_16G_out.awready),
       .m_axi_wdata    (axi_m_00G_16G_out.wdata),
       .m_axi_wstrb    (axi_m_00G_16G_out.wstrb),
       .m_axi_wlast    (axi_m_00G_16G_out.wlast),
       .m_axi_wvalid   (axi_m_00G_16G_out.wvalid),
       .m_axi_wready   (axi_m_00G_16G_out.wready),
       .m_axi_bid      (axi_m_00G_16G_out.bid),
       .m_axi_bresp    (axi_m_00G_16G_out.bresp),
       .m_axi_bvalid   (axi_m_00G_16G_out.bvalid),
       .m_axi_bready   (axi_m_00G_16G_out.bready),
       .m_axi_arid     (axi_m_00G_16G_out.arid),
       .m_axi_araddr   (axi_m_00G_16G_out.araddr),
       .m_axi_arlen    (axi_m_00G_16G_out.arlen),
       .m_axi_arsize   (axi_m_00G_16G_out.arsize),
       .m_axi_arburst  (),
       .m_axi_arlock   (),
       .m_axi_arcache  (),
       .m_axi_arprot   (),
       .m_axi_arregion (),
       .m_axi_arqos    (),
       .m_axi_arvalid  (axi_m_00G_16G_out.arvalid),
       .m_axi_arready  (axi_m_00G_16G_out.arready),
       .m_axi_rid      (axi_m_00G_16G_out.rid),
       .m_axi_rdata    (axi_m_00G_16G_out.rdata),
       .m_axi_rresp    (axi_m_00G_16G_out.rresp),
       .m_axi_rlast    (axi_m_00G_16G_out.rlast),
       .m_axi_rvalid   (axi_m_00G_16G_out.rvalid),
       .m_axi_rready   (axi_m_00G_16G_out.rready)
       );

//----------------------------
// flop the output of interconnect 32G-48G
//----------------------------
   axi_register_slice AXI4_REG_SLC_32G_48G_1 (
       .aclk           (aclk),
       .aresetn        (slr1_sync_aresetn),

       .s_axi_awid     (axi_m_32G_48G_0.awid),
       .s_axi_awaddr   ({axi_m_32G_48G_0.awaddr[63:36], 2'b0, axi_m_32G_48G_0.awaddr[33:0]}),
       .s_axi_awlen    (axi_m_32G_48G_0.awlen),
       .s_axi_awsize   (axi_m_32G_48G_0.awsize),
       .s_axi_awvalid  (axi_m_32G_48G_0.awvalid),
       .s_axi_awready  (axi_m_32G_48G_0.awready),
       .s_axi_wdata    (axi_m_32G_48G_0.wdata),
       .s_axi_wstrb    (axi_m_32G_48G_0.wstrb),
       .s_axi_wlast    (axi_m_32G_48G_0.wlast),
       .s_axi_wvalid   (axi_m_32G_48G_0.wvalid),
       .s_axi_wready   (axi_m_32G_48G_0.wready),
       .s_axi_bid      (axi_m_32G_48G_0.bid),
       .s_axi_bresp    (axi_m_32G_48G_0.bresp),
       .s_axi_bvalid   (axi_m_32G_48G_0.bvalid),
       .s_axi_bready   (axi_m_32G_48G_0.bready),
       .s_axi_arid     (axi_m_32G_48G_0.arid),
       .s_axi_araddr   ({axi_m_32G_48G_0.araddr[63:36], 2'b0, axi_m_32G_48G_0.araddr[33:0]}),
       .s_axi_arlen    (axi_m_32G_48G_0.arlen),
       .s_axi_arsize   (axi_m_32G_48G_0.arsize),
       .s_axi_arvalid  (axi_m_32G_48G_0.arvalid),
       .s_axi_arready  (axi_m_32G_48G_0.arready),
       .s_axi_rid      (axi_m_32G_48G_0.rid),
       .s_axi_rdata    (axi_m_32G_48G_0.rdata),
       .s_axi_rresp    (axi_m_32G_48G_0.rresp),
       .s_axi_rlast    (axi_m_32G_48G_0.rlast),
       .s_axi_rvalid   (axi_m_32G_48G_0.rvalid),
       .s_axi_rready   (axi_m_32G_48G_0.rready),
       .m_axi_awid     (axi_m_32G_48G_2.awid),
       .m_axi_awaddr   (axi_m_32G_48G_2.awaddr),
       .m_axi_awlen    (axi_m_32G_48G_2.awlen),
       .m_axi_awsize   (axi_m_32G_48G_2.awsize),
       .m_axi_awvalid  (axi_m_32G_48G_2.awvalid),
       .m_axi_awready  (axi_m_32G_48G_2.awready),
       .m_axi_wdata    (axi_m_32G_48G_2.wdata),
       .m_axi_wstrb    (axi_m_32G_48G_2.wstrb),
       .m_axi_wlast    (axi_m_32G_48G_2.wlast),
       .m_axi_wvalid   (axi_m_32G_48G_2.wvalid),
       .m_axi_wready   (axi_m_32G_48G_2.wready),
       .m_axi_bid      (axi_m_32G_48G_2.bid),
       .m_axi_bresp    (axi_m_32G_48G_2.bresp),
       .m_axi_bvalid   (axi_m_32G_48G_2.bvalid),
       .m_axi_bready   (axi_m_32G_48G_2.bready),
       .m_axi_arid     (axi_m_32G_48G_2.arid),
       .m_axi_araddr   (axi_m_32G_48G_2.araddr),
       .m_axi_arlen    (axi_m_32G_48G_2.arlen),
       .m_axi_arsize   (axi_m_32G_48G_2.arsize),
       .m_axi_arvalid  (axi_m_32G_48G_2.arvalid),
       .m_axi_arready  (axi_m_32G_48G_2.arready),
       .m_axi_rid      (axi_m_32G_48G_2.rid),
       .m_axi_rdata    (axi_m_32G_48G_2.rdata),
       .m_axi_rresp    (axi_m_32G_48G_2.rresp),
       .m_axi_rlast    (axi_m_32G_48G_2.rlast),
       .m_axi_rvalid   (axi_m_32G_48G_2.rvalid),
       .m_axi_rready   (axi_m_32G_48G_2.rready)
   );
   axi_register_slice AXI4_REG_SLC_32G_48G_2 (
       .aclk           (aclk),
       .aresetn        (slr1_sync_aresetn),

       .s_axi_awid     (axi_m_32G_48G_2.awid),
       .s_axi_awaddr   ({axi_m_32G_48G_2.awaddr[63:36], 2'b0, axi_m_32G_48G_2.awaddr[33:0]}),
       .s_axi_awlen    (axi_m_32G_48G_2.awlen),
       .s_axi_awsize   (axi_m_32G_48G_2.awsize),
       .s_axi_awvalid  (axi_m_32G_48G_2.awvalid),
       .s_axi_awready  (axi_m_32G_48G_2.awready),
       .s_axi_wdata    (axi_m_32G_48G_2.wdata),
       .s_axi_wstrb    (axi_m_32G_48G_2.wstrb),
       .s_axi_wlast    (axi_m_32G_48G_2.wlast),
       .s_axi_wvalid   (axi_m_32G_48G_2.wvalid),
       .s_axi_wready   (axi_m_32G_48G_2.wready),
       .s_axi_bid      (axi_m_32G_48G_2.bid),
       .s_axi_bresp    (axi_m_32G_48G_2.bresp),
       .s_axi_bvalid   (axi_m_32G_48G_2.bvalid),
       .s_axi_bready   (axi_m_32G_48G_2.bready),
       .s_axi_arid     (axi_m_32G_48G_2.arid),
       .s_axi_araddr   ({axi_m_32G_48G_2.araddr[63:36], 2'b0, axi_m_32G_48G_2.araddr[33:0]}),
       .s_axi_arlen    (axi_m_32G_48G_2.arlen),
       .s_axi_arsize   (axi_m_32G_48G_2.arsize),
       .s_axi_arvalid  (axi_m_32G_48G_2.arvalid),
       .s_axi_arready  (axi_m_32G_48G_2.arready),
       .s_axi_rid      (axi_m_32G_48G_2.rid),
       .s_axi_rdata    (axi_m_32G_48G_2.rdata),
       .s_axi_rresp    (axi_m_32G_48G_2.rresp),
       .s_axi_rlast    (axi_m_32G_48G_2.rlast),
       .s_axi_rvalid   (axi_m_32G_48G_2.rvalid),
       .s_axi_rready   (axi_m_32G_48G_2.rready),
       .m_axi_awid     (axi_m_32G_48G_out.awid),
       .m_axi_awaddr   (axi_m_32G_48G_out.awaddr),
       .m_axi_awlen    (axi_m_32G_48G_out.awlen),
       .m_axi_awsize   (axi_m_32G_48G_out.awsize),
       .m_axi_awvalid  (axi_m_32G_48G_out.awvalid),
       .m_axi_awready  (axi_m_32G_48G_out.awready),
       .m_axi_wdata    (axi_m_32G_48G_out.wdata),
       .m_axi_wstrb    (axi_m_32G_48G_out.wstrb),
       .m_axi_wlast    (axi_m_32G_48G_out.wlast),
       .m_axi_wvalid   (axi_m_32G_48G_out.wvalid),
       .m_axi_wready   (axi_m_32G_48G_out.wready),
       .m_axi_bid      (axi_m_32G_48G_out.bid),
       .m_axi_bresp    (axi_m_32G_48G_out.bresp),
       .m_axi_bvalid   (axi_m_32G_48G_out.bvalid),
       .m_axi_bready   (axi_m_32G_48G_out.bready),
       .m_axi_arid     (axi_m_32G_48G_out.arid),
       .m_axi_araddr   (axi_m_32G_48G_out.araddr),
       .m_axi_arlen    (axi_m_32G_48G_out.arlen),
       .m_axi_arsize   (axi_m_32G_48G_out.arsize),
       .m_axi_arvalid  (axi_m_32G_48G_out.arvalid),
       .m_axi_arready  (axi_m_32G_48G_out.arready),
       .m_axi_rid      (axi_m_32G_48G_out.rid),
       .m_axi_rdata    (axi_m_32G_48G_out.rdata),
       .m_axi_rresp    (axi_m_32G_48G_out.rresp),
       .m_axi_rlast    (axi_m_32G_48G_out.rlast),
       .m_axi_rvalid   (axi_m_32G_48G_out.rvalid),
       .m_axi_rready   (axi_m_32G_48G_out.rready)
   );

//----------------------------
// flop the output of interconnect for DDRB
// back to back for SLR crossing
//----------------------------

  //back to back register slices for SLR crossing
   src_register_slice DDR_B_TST_AXI4_REG_SLC_1 (
       .aclk           (aclk),
       .aresetn        (slr1_sync_aresetn),
       .s_axi_awid     (axi_m_16G_32G_0.awid),
       .s_axi_awaddr   ({axi_m_16G_32G_0.awaddr[63:36], 2'b0, axi_m_16G_32G_0.awaddr[33:0]}),
       .s_axi_awlen    (axi_m_16G_32G_0.awlen),
       .s_axi_awsize   (axi_m_16G_32G_0.awsize),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (axi_m_16G_32G_0.awvalid),
       .s_axi_awready  (axi_m_16G_32G_0.awready),
       .s_axi_wdata    (axi_m_16G_32G_0.wdata),
       .s_axi_wstrb    (axi_m_16G_32G_0.wstrb),
       .s_axi_wlast    (axi_m_16G_32G_0.wlast),
       .s_axi_wvalid   (axi_m_16G_32G_0.wvalid),
       .s_axi_wready   (axi_m_16G_32G_0.wready),
       .s_axi_bid      (axi_m_16G_32G_0.bid),
       .s_axi_bresp    (axi_m_16G_32G_0.bresp),
       .s_axi_bvalid   (axi_m_16G_32G_0.bvalid),
       .s_axi_bready   (axi_m_16G_32G_0.bready),
       .s_axi_arid     (axi_m_16G_32G_0.arid),
       .s_axi_araddr   ({axi_m_16G_32G_0.araddr[63:36], 2'b0, axi_m_16G_32G_0.araddr[33:0]}),
       .s_axi_arlen    (axi_m_16G_32G_0.arlen),
       .s_axi_arsize   (axi_m_16G_32G_0.arsize),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (axi_m_16G_32G_0.arvalid),
       .s_axi_arready  (axi_m_16G_32G_0.arready),
       .s_axi_rid      (axi_m_16G_32G_0.rid),
       .s_axi_rdata    (axi_m_16G_32G_0.rdata),
       .s_axi_rresp    (axi_m_16G_32G_0.rresp),
       .s_axi_rlast    (axi_m_16G_32G_0.rlast),
       .s_axi_rvalid   (axi_m_16G_32G_0.rvalid),
       .s_axi_rready   (axi_m_16G_32G_0.rready),
       .m_axi_awid     (axi_m_16G_32G_2.awid),
       .m_axi_awaddr   (axi_m_16G_32G_2.awaddr),
       .m_axi_awlen    (axi_m_16G_32G_2.awlen),
       .m_axi_awsize   (axi_m_16G_32G_2.awsize),
       .m_axi_awburst  (),
       .m_axi_awlock   (),
       .m_axi_awcache  (),
       .m_axi_awprot   (),
       .m_axi_awregion (),
       .m_axi_awqos    (),
       .m_axi_awvalid  (axi_m_16G_32G_2.awvalid),
       .m_axi_awready  (axi_m_16G_32G_2.awready),
       .m_axi_wdata    (axi_m_16G_32G_2.wdata),
       .m_axi_wstrb    (axi_m_16G_32G_2.wstrb),
       .m_axi_wlast    (axi_m_16G_32G_2.wlast),
       .m_axi_wvalid   (axi_m_16G_32G_2.wvalid),
       .m_axi_wready   (axi_m_16G_32G_2.wready),
       .m_axi_bid      (axi_m_16G_32G_2.bid),
       .m_axi_bresp    (axi_m_16G_32G_2.bresp),
       .m_axi_bvalid   (axi_m_16G_32G_2.bvalid),
       .m_axi_bready   (axi_m_16G_32G_2.bready),
       .m_axi_arid     (axi_m_16G_32G_2.arid),
       .m_axi_araddr   (axi_m_16G_32G_2.araddr),
       .m_axi_arlen    (axi_m_16G_32G_2.arlen),
       .m_axi_arsize   (axi_m_16G_32G_2.arsize),
       .m_axi_arburst  (),
       .m_axi_arlock   (),
       .m_axi_arcache  (),
       .m_axi_arprot   (),
       .m_axi_arregion (),
       .m_axi_arqos    (),
       .m_axi_arvalid  (axi_m_16G_32G_2.arvalid),
       .m_axi_arready  (axi_m_16G_32G_2.arready),
       .m_axi_rid      (axi_m_16G_32G_2.rid),
       .m_axi_rdata    (axi_m_16G_32G_2.rdata),
       .m_axi_rresp    (axi_m_16G_32G_2.rresp),
       .m_axi_rlast    (axi_m_16G_32G_2.rlast),
       .m_axi_rvalid   (axi_m_16G_32G_2.rvalid),
       .m_axi_rready   (axi_m_16G_32G_2.rready)
       );
   dest_register_slice DDR_B_TST_AXI4_REG_SLC_2 (
       .aclk           (aclk),
       .aresetn        (slr1_sync_aresetn),
       .s_axi_awid     (axi_m_16G_32G_2.awid),
       .s_axi_awaddr   (axi_m_16G_32G_2.awaddr),
       .s_axi_awlen    (axi_m_16G_32G_2.awlen),
       .s_axi_awsize   (axi_m_16G_32G_2.awsize),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (axi_m_16G_32G_2.awvalid),
       .s_axi_awready  (axi_m_16G_32G_2.awready),
       .s_axi_wdata    (axi_m_16G_32G_2.wdata),
       .s_axi_wstrb    (axi_m_16G_32G_2.wstrb),
       .s_axi_wlast    (axi_m_16G_32G_2.wlast),
       .s_axi_wvalid   (axi_m_16G_32G_2.wvalid),
       .s_axi_wready   (axi_m_16G_32G_2.wready),
       .s_axi_bid      (axi_m_16G_32G_2.bid),
       .s_axi_bresp    (axi_m_16G_32G_2.bresp),
       .s_axi_bvalid   (axi_m_16G_32G_2.bvalid),
       .s_axi_bready   (axi_m_16G_32G_2.bready),
       .s_axi_arid     (axi_m_16G_32G_2.arid),
       .s_axi_araddr   (axi_m_16G_32G_2.araddr),
       .s_axi_arlen    (axi_m_16G_32G_2.arlen),
       .s_axi_arsize   (axi_m_16G_32G_2.arsize),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (axi_m_16G_32G_2.arvalid),
       .s_axi_arready  (axi_m_16G_32G_2.arready),
       .s_axi_rid      (axi_m_16G_32G_2.rid),
       .s_axi_rdata    (axi_m_16G_32G_2.rdata),
       .s_axi_rresp    (axi_m_16G_32G_2.rresp),
       .s_axi_rlast    (axi_m_16G_32G_2.rlast),
       .s_axi_rvalid   (axi_m_16G_32G_2.rvalid),
       .s_axi_rready   (axi_m_16G_32G_2.rready),
       .m_axi_awid     (axi_m_16G_32G_out.awid),
       .m_axi_awaddr   (axi_m_16G_32G_out.awaddr),
       .m_axi_awlen    (axi_m_16G_32G_out.awlen),
       .m_axi_awsize   (axi_m_16G_32G_out.awsize),
       .m_axi_awburst  (),
       .m_axi_awlock   (),
       .m_axi_awcache  (),
       .m_axi_awprot   (),
       .m_axi_awregion (),
       .m_axi_awqos    (),
       .m_axi_awvalid  (axi_m_16G_32G_out.awvalid),
       .m_axi_awready  (axi_m_16G_32G_out.awready),
       .m_axi_wdata    (axi_m_16G_32G_out.wdata),
       .m_axi_wstrb    (axi_m_16G_32G_out.wstrb),
       .m_axi_wlast    (axi_m_16G_32G_out.wlast),
       .m_axi_wvalid   (axi_m_16G_32G_out.wvalid),
       .m_axi_wready   (axi_m_16G_32G_out.wready),
       .m_axi_bid      (axi_m_16G_32G_out.bid),
       .m_axi_bresp    (axi_m_16G_32G_out.bresp),
       .m_axi_bvalid   (axi_m_16G_32G_out.bvalid),
       .m_axi_bready   (axi_m_16G_32G_out.bready),
       .m_axi_arid     (axi_m_16G_32G_out.arid),
       .m_axi_araddr   (axi_m_16G_32G_out.araddr),
       .m_axi_arlen    (axi_m_16G_32G_out.arlen),
       .m_axi_arsize   (axi_m_16G_32G_out.arsize),
       .m_axi_arburst  (),
       .m_axi_arlock   (),
       .m_axi_arcache  (),
       .m_axi_arprot   (),
       .m_axi_arregion (),
       .m_axi_arqos    (),
       .m_axi_arvalid  (axi_m_16G_32G_out.arvalid),
       .m_axi_arready  (axi_m_16G_32G_out.arready),
       .m_axi_rid      (axi_m_16G_32G_out.rid),
       .m_axi_rdata    (axi_m_16G_32G_out.rdata),
       .m_axi_rresp    (axi_m_16G_32G_out.rresp),
       .m_axi_rlast    (axi_m_16G_32G_out.rlast),
       .m_axi_rvalid   (axi_m_16G_32G_out.rvalid),
       .m_axi_rready   (axi_m_16G_32G_out.rready)
       );

//----------------------------
// ATG/scrubber for DDRA
//----------------------------
   lib_pipe #(.WIDTH(32+32+1+1), .STAGES(NUM_CFG_STGS_CL_DDR_ATG)) PIPE_CFG_REQ_DDR_A (.clk (aclk),
                                                              .rst_n (aresetn),
                                                              .in_bus({ddra_tst_cfg_bus.addr, ddra_tst_cfg_bus.wdata, ddra_tst_cfg_bus.wr, ddra_tst_cfg_bus.rd}),
                                                              .out_bus({ddra_tst_cfg_bus_q.addr, ddra_tst_cfg_bus_q.wdata, ddra_tst_cfg_bus_q.wr, ddra_tst_cfg_bus_q.rd})
                                                              );

   lib_pipe #(.WIDTH(32+1), .STAGES(NUM_CFG_STGS_CL_DDR_ATG)) PIPE_CFG_ACK_DDR_A (.clk (aclk),
                                                              .rst_n (aresetn),
                                                              .in_bus({ddra_tst_cfg_bus_q.ack, ddra_tst_cfg_bus_q.rdata}),
                                                              .out_bus({ddra_tst_cfg_bus.ack, ddra_tst_cfg_bus.rdata})
                                                              );


   lib_pipe #(.WIDTH(2+3+64), .STAGES(NUM_CFG_STGS_CL_DDR_ATG)) PIPE_SCRB_DDR_A (.clk(aclk),
                                                              .rst_n(aresetn),
                                                              .in_bus({ddra_scrb_bus.enable, ddra_scrb_bus_q.done, ddra_scrb_bus_q.state, ddra_scrb_bus_q.addr}),
                                                              .out_bus({ddra_scrb_bus_q.enable, ddra_scrb_bus.done, ddra_scrb_bus.state, ddra_scrb_bus.addr})
                                                              );

   cl_tst_scrb #(.DATA_WIDTH(512),
                    .SCRB_BURST_LEN_MINUS1(SCRB_BURST_LEN_MINUS1),
                    .SCRB_MAX_ADDR(SCRB_MAX_ADDR),
                    .NO_SCRB_INST(NO_SCRB_INST)) CL_TST_DDR_A (

         .clk(aclk),
         .rst_n(slr2_sync_aresetn),

         .cfg_addr(ddra_tst_cfg_bus_q.addr),
         .cfg_wdata(ddra_tst_cfg_bus_q.wdata),
         .cfg_wr(ddra_tst_cfg_bus_q.wr),
         .cfg_rd(ddra_tst_cfg_bus_q.rd),
         .tst_cfg_ack(ddra_tst_cfg_bus_q.ack),
         .tst_cfg_rdata(ddra_tst_cfg_bus_q.rdata),

         .slv_awid(ddra_axi_slv.awid[6:0]),
         .slv_awaddr(ddra_axi_slv.awaddr),
         .slv_awlen(ddra_axi_slv.awlen),
         .slv_awsize(ddra_axi_slv.awsize),
         .slv_awvalid(ddra_axi_slv.awvalid),
         .slv_awuser(11'b0),
         .slv_awready(ddra_axi_slv.awready),

         .slv_wid(7'b0),
         .slv_wdata(ddra_axi_slv.wdata),
         .slv_wstrb(ddra_axi_slv.wstrb),
         .slv_wlast(ddra_axi_slv.wlast),
         .slv_wvalid(ddra_axi_slv.wvalid),
         .slv_wready(ddra_axi_slv.wready),

         .slv_bid(ddra_axi_slv.bid[6:0]),
         .slv_bresp(ddra_axi_slv.bresp),
         .slv_buser(),
         .slv_bvalid(ddra_axi_slv.bvalid),
         .slv_bready(ddra_axi_slv.bready),

         .slv_arid(ddra_axi_slv.arid[6:0]),
         .slv_araddr(ddra_axi_slv.araddr),
         .slv_arlen(ddra_axi_slv.arlen),
         .slv_arsize(ddra_axi_slv.arsize),
         .slv_arvalid(ddra_axi_slv.arvalid),
         .slv_aruser(11'b0),
         .slv_arready(ddra_axi_slv.arready),

         .slv_rid(ddra_axi_slv.rid[6:0]),
         .slv_rdata(ddra_axi_slv.rdata),
         .slv_rresp(ddra_axi_slv.rresp),
         .slv_rlast(ddra_axi_slv.rlast),
         .slv_ruser(),
         .slv_rvalid(ddra_axi_slv.rvalid),
         .slv_rready(ddra_axi_slv.rready),


         .awid(lcl_cl_sh_ddra.awid[8:0]),
         .awaddr(lcl_cl_sh_ddra.awaddr),
         .awlen(lcl_cl_sh_ddra.awlen),
         .awsize(lcl_cl_sh_ddra.awsize),
         .awvalid(lcl_cl_sh_ddra.awvalid),
         .awuser(),
         .awready(lcl_cl_sh_ddra.awready),

         .wid(lcl_cl_sh_ddra.wid[8:0]),
         .wdata(lcl_cl_sh_ddra.wdata),
         .wstrb(lcl_cl_sh_ddra.wstrb),
         .wlast(lcl_cl_sh_ddra.wlast),
         .wvalid(lcl_cl_sh_ddra.wvalid),
         .wready(lcl_cl_sh_ddra.wready),

         .bid(lcl_cl_sh_ddra.bid[8:0]),
         .bresp(lcl_cl_sh_ddra.bresp),
         .buser(18'h0),
         .bvalid(lcl_cl_sh_ddra.bvalid),
         .bready(lcl_cl_sh_ddra.bready),

         .arid(lcl_cl_sh_ddra.arid[8:0]),
         .araddr(lcl_cl_sh_ddra.araddr),
         .arlen(lcl_cl_sh_ddra.arlen),
         .arsize(lcl_cl_sh_ddra.arsize),
         .arvalid(lcl_cl_sh_ddra.arvalid),
         .aruser(),
         .arready(lcl_cl_sh_ddra.arready),

         .rid(lcl_cl_sh_ddra.rid[8:0]),
         .rdata(lcl_cl_sh_ddra.rdata),
         .rresp(lcl_cl_sh_ddra.rresp),
         .rlast(lcl_cl_sh_ddra.rlast),
         .ruser(18'h0),
         .rvalid(lcl_cl_sh_ddra.rvalid),
         .rready(lcl_cl_sh_ddra.rready),

         .scrb_enable(ddra_scrb_bus_q.enable),
         .scrb_done  (ddra_scrb_bus_q.done),

         .scrb_dbg_state(ddra_scrb_bus_q.state),
         .scrb_dbg_addr (ddra_scrb_bus_q.addr)
      );
      assign lcl_cl_sh_ddra.awid[15:9] = 7'b0;
      assign lcl_cl_sh_ddra.wid[15:9] = 7'b0;
      assign lcl_cl_sh_ddra.arid[15:9] = 7'b0;

//----------------------------
// ATG/scrubber for DDRB
//----------------------------
   lib_pipe #(.WIDTH(32+32+1+1), .STAGES(NUM_CFG_STGS_CL_DDR_ATG)) PIPE_CFG_REQ_DDR_B (.clk (aclk),
                                                              .rst_n (aresetn),
                                                              .in_bus({ddrb_tst_cfg_bus.addr, ddrb_tst_cfg_bus.wdata, ddrb_tst_cfg_bus.wr, ddrb_tst_cfg_bus.rd}),
                                                              .out_bus({ddrb_tst_cfg_bus_q.addr, ddrb_tst_cfg_bus_q.wdata, ddrb_tst_cfg_bus_q.wr, ddrb_tst_cfg_bus_q.rd})
                                                              );

   lib_pipe #(.WIDTH(32+1), .STAGES(NUM_CFG_STGS_CL_DDR_ATG)) PIPE_CFG_ACK_DDR_B (.clk (aclk),
                                                              .rst_n (aresetn),
                                                              .in_bus({ddrb_tst_cfg_bus_q.ack, ddrb_tst_cfg_bus_q.rdata}),
                                                              .out_bus({ddrb_tst_cfg_bus.ack, ddrb_tst_cfg_bus.rdata})
                                                              );


   lib_pipe #(.WIDTH(2+3+64), .STAGES(NUM_CFG_STGS_CL_DDR_ATG)) PIPE_SCRB_DDR_B (.clk(aclk),
                                                              .rst_n(aresetn),
                                                              .in_bus({ddrb_scrb_bus.enable, ddrb_scrb_bus_q.done, ddrb_scrb_bus_q.state, ddrb_scrb_bus_q.addr}),
                                                              .out_bus({ddrb_scrb_bus_q.enable, ddrb_scrb_bus.done, ddrb_scrb_bus.state, ddrb_scrb_bus.addr})
                                                              );

   cl_tst_scrb #(.DATA_WIDTH(512),
                    .SCRB_BURST_LEN_MINUS1(SCRB_BURST_LEN_MINUS1),
                    .SCRB_MAX_ADDR(SCRB_MAX_ADDR),
                    .NO_SCRB_INST(NO_SCRB_INST)) CL_TST_DDR_B (

         .clk(aclk),
         .rst_n(slr1_sync_aresetn),

         .cfg_addr(ddrb_tst_cfg_bus_q.addr),
         .cfg_wdata(ddrb_tst_cfg_bus_q.wdata),
         .cfg_wr(ddrb_tst_cfg_bus_q.wr),
         .cfg_rd(ddrb_tst_cfg_bus_q.rd),
         .tst_cfg_ack(ddrb_tst_cfg_bus_q.ack),
         .tst_cfg_rdata(ddrb_tst_cfg_bus_q.rdata),

         .slv_awid(ddrb_axi_slv.awid[6:0]),
         .slv_awaddr(ddrb_axi_slv.awaddr),
         .slv_awlen(ddrb_axi_slv.awlen),
         .slv_awsize(ddrb_axi_slv.awsize),
         .slv_awvalid(ddrb_axi_slv.awvalid),
         .slv_awuser(11'b0),
         .slv_awready(ddrb_axi_slv.awready),

         .slv_wid(7'b0),
         .slv_wdata(ddrb_axi_slv.wdata),
         .slv_wstrb(ddrb_axi_slv.wstrb),
         .slv_wlast(ddrb_axi_slv.wlast),
         .slv_wvalid(ddrb_axi_slv.wvalid),
         .slv_wready(ddrb_axi_slv.wready),

         .slv_bid(ddrb_axi_slv.bid[6:0]),
         .slv_bresp(ddrb_axi_slv.bresp),
         .slv_buser(),
         .slv_bvalid(ddrb_axi_slv.bvalid),
         .slv_bready(ddrb_axi_slv.bready),

         .slv_arid(ddrb_axi_slv.arid[6:0]),
         .slv_araddr(ddrb_axi_slv.araddr),
         .slv_arlen(ddrb_axi_slv.arlen),
         .slv_arsize(ddrb_axi_slv.arsize),
         .slv_arvalid(ddrb_axi_slv.arvalid),
         .slv_aruser(11'b0),
         .slv_arready(ddrb_axi_slv.arready),

         .slv_rid(ddrb_axi_slv.rid[6:0]),
         .slv_rdata(ddrb_axi_slv.rdata),
         .slv_rresp(ddrb_axi_slv.rresp),
         .slv_rlast(ddrb_axi_slv.rlast),
         .slv_ruser(),
         .slv_rvalid(ddrb_axi_slv.rvalid),
         .slv_rready(ddrb_axi_slv.rready),


         .awid(lcl_cl_sh_ddrb.awid[8:0]),
         .awaddr(lcl_cl_sh_ddrb.awaddr),
         .awlen(lcl_cl_sh_ddrb.awlen),
         .awsize(lcl_cl_sh_ddrb.awsize),
         .awvalid(lcl_cl_sh_ddrb.awvalid),
         .awuser(),
         .awready(lcl_cl_sh_ddrb.awready),

         .wid(lcl_cl_sh_ddrb.wid[8:0]),
         .wdata(lcl_cl_sh_ddrb.wdata),
         .wstrb(lcl_cl_sh_ddrb.wstrb),
         .wlast(lcl_cl_sh_ddrb.wlast),
         .wvalid(lcl_cl_sh_ddrb.wvalid),
         .wready(lcl_cl_sh_ddrb.wready),

         .bid(lcl_cl_sh_ddrb.bid[8:0]),
         .bresp(lcl_cl_sh_ddrb.bresp),
         .buser(18'h0),
         .bvalid(lcl_cl_sh_ddrb.bvalid),
         .bready(lcl_cl_sh_ddrb.bready),

         .arid(lcl_cl_sh_ddrb.arid[8:0]),
         .araddr(lcl_cl_sh_ddrb.araddr),
         .arlen(lcl_cl_sh_ddrb.arlen),
         .arsize(lcl_cl_sh_ddrb.arsize),
         .arvalid(lcl_cl_sh_ddrb.arvalid),
         .aruser(),
         .arready(lcl_cl_sh_ddrb.arready),

         .rid(lcl_cl_sh_ddrb.rid[8:0]),
         .rdata(lcl_cl_sh_ddrb.rdata),
         .rresp(lcl_cl_sh_ddrb.rresp),
         .rlast(lcl_cl_sh_ddrb.rlast),
         .ruser(18'h0),
         .rvalid(lcl_cl_sh_ddrb.rvalid),
         .rready(lcl_cl_sh_ddrb.rready),

         .scrb_enable(ddrb_scrb_bus_q.enable),
         .scrb_done  (ddrb_scrb_bus_q.done),

         .scrb_dbg_state(ddrb_scrb_bus_q.state),
         .scrb_dbg_addr (ddrb_scrb_bus_q.addr)
      );
      assign lcl_cl_sh_ddrb.awid[15:9] = 7'b0;
      assign lcl_cl_sh_ddrb.wid[15:9] = 7'b0;
      assign lcl_cl_sh_ddrb.arid[15:9] = 7'b0;


//----------------------------
// ATG/scrubber for DDRC
//----------------------------

   lib_pipe #(.WIDTH(32+32+1+1), .STAGES(NUM_CFG_STGS_SH_DDR_ATG)) PIPE_CFG_REQ_DDR_C (.clk (aclk),
                                                              .rst_n (aresetn),
                                                              .in_bus({ddrc_tst_cfg_bus.addr, ddrc_tst_cfg_bus.wdata, ddrc_tst_cfg_bus.wr, ddrc_tst_cfg_bus.rd}),
                                                              .out_bus({ddrc_tst_cfg_bus_q.addr, ddrc_tst_cfg_bus_q.wdata, ddrc_tst_cfg_bus_q.wr, ddrc_tst_cfg_bus_q.rd})
                                                              );

   lib_pipe #(.WIDTH(32+1), .STAGES(NUM_CFG_STGS_SH_DDR_ATG)) PIPE_CFG_ACK_DDR_C (.clk (aclk),
                                                              .rst_n (aresetn),
                                                              .in_bus({ddrc_tst_cfg_bus_q.ack, ddrc_tst_cfg_bus_q.rdata}),
                                                              .out_bus({ddrc_tst_cfg_bus.ack, ddrc_tst_cfg_bus.rdata})
                                                              );


   lib_pipe #(.WIDTH(2+3+64), .STAGES(NUM_CFG_STGS_SH_DDR_ATG)) PIPE_SCRB_DDR_C (.clk(aclk),
                                                              .rst_n(aresetn),
                                                              .in_bus({ddrc_scrb_bus.enable, ddrc_scrb_bus_q.done, ddrc_scrb_bus_q.state, ddrc_scrb_bus_q.addr}),
                                                              .out_bus({ddrc_scrb_bus_q.enable, ddrc_scrb_bus.done, ddrc_scrb_bus.state, ddrc_scrb_bus.addr})
                                                              );
   cl_tst_scrb #(.DATA_WIDTH(512),
                    .SCRB_BURST_LEN_MINUS1(SCRB_BURST_LEN_MINUS1),
                    .SCRB_MAX_ADDR(SCRB_MAX_ADDR),
                    .NO_SCRB_INST(NO_SCRB_INST)) CL_TST_DDR_C (

         .clk(aclk),
         .rst_n(slr1_sync_aresetn),

         .cfg_addr(ddrc_tst_cfg_bus_q.addr),
         .cfg_wdata(ddrc_tst_cfg_bus_q.wdata),
         .cfg_wr(ddrc_tst_cfg_bus_q.wr),
         .cfg_rd(ddrc_tst_cfg_bus_q.rd),
         .tst_cfg_ack(ddrc_tst_cfg_bus_q.ack),
         .tst_cfg_rdata(ddrc_tst_cfg_bus_q.rdata),

         .slv_awid(ddrc_axi_slv.awid[6:0]),
         .slv_awaddr(ddrc_axi_slv.awaddr),
         .slv_awlen(ddrc_axi_slv.awlen),
         .slv_awvalid(ddrc_axi_slv.awvalid),
         .slv_awsize(ddrc_axi_slv.awsize),
         .slv_awuser(11'b0),
         .slv_awready(ddrc_axi_slv.awready),

         .slv_wid(7'b0),
         .slv_wdata(ddrc_axi_slv.wdata),
         .slv_wstrb(ddrc_axi_slv.wstrb),
         .slv_wlast(ddrc_axi_slv.wlast),
         .slv_wvalid(ddrc_axi_slv.wvalid),
         .slv_wready(ddrc_axi_slv.wready),

         .slv_bid(ddrc_axi_slv.bid[6:0]),
         .slv_bresp(ddrc_axi_slv.bresp),
         .slv_buser(),
         .slv_bvalid(ddrc_axi_slv.bvalid),
         .slv_bready(ddrc_axi_slv.bready),

         .slv_arid(ddrc_axi_slv.arid[6:0]),
         .slv_araddr(ddrc_axi_slv.araddr),
         .slv_arlen(ddrc_axi_slv.arlen),
         .slv_arvalid(ddrc_axi_slv.arvalid),
         .slv_arsize(ddrc_axi_slv.arsize),
         .slv_aruser(11'b0),
         .slv_arready(ddrc_axi_slv.arready),

         .slv_rid(ddrc_axi_slv.rid[6:0]),
         .slv_rdata(ddrc_axi_slv.rdata),
         .slv_rresp(ddrc_axi_slv.rresp),
         .slv_rlast(ddrc_axi_slv.rlast),
         .slv_ruser(),
         .slv_rvalid(ddrc_axi_slv.rvalid),
         .slv_rready(ddrc_axi_slv.rready),


         .awid(ddrc_axi_mstr.awid[8:0]),
         .awaddr(ddrc_axi_mstr.awaddr),
         .awlen(ddrc_axi_mstr.awlen),
         .awvalid(ddrc_axi_mstr.awvalid),
         .awsize(ddrc_axi_mstr.awsize),
         .awuser(),
         .awready(ddrc_axi_mstr.awready),

         //.wid(ddrc_axi_mstr.wid),
         .wid(),
         .wdata(ddrc_axi_mstr.wdata),
         .wstrb(ddrc_axi_mstr.wstrb),
         .wlast(ddrc_axi_mstr.wlast),
         .wvalid(ddrc_axi_mstr.wvalid),
         .wready(ddrc_axi_mstr.wready),

         .bid(ddrc_axi_mstr.bid[8:0]),
         .bresp(ddrc_axi_mstr.bresp),
         .buser(18'h0),
         .bvalid(ddrc_axi_mstr.bvalid),
         .bready(ddrc_axi_mstr.bready),

         .arid(ddrc_axi_mstr.arid[8:0]),
         .araddr(ddrc_axi_mstr.araddr),
         .arlen(ddrc_axi_mstr.arlen),
         .arvalid(ddrc_axi_mstr.arvalid),
         .arsize(ddrc_axi_mstr.arsize),
         .aruser(),
         .arready(ddrc_axi_mstr.arready),

         .rid(ddrc_axi_mstr.rid[8:0]),
         .rdata(ddrc_axi_mstr.rdata),
         .rresp(ddrc_axi_mstr.rresp),
         .rlast(ddrc_axi_mstr.rlast),
         .ruser(18'h0),
         .rvalid(ddrc_axi_mstr.rvalid),
         .rready(ddrc_axi_mstr.rready),

         .scrb_enable(ddrc_scrb_bus_q.enable),
         .scrb_done  (ddrc_scrb_bus_q.done),

         .scrb_dbg_state(ddrc_scrb_bus_q.state),
         .scrb_dbg_addr (ddrc_scrb_bus_q.addr)
   );

//----------------------------
// flop the output of ATG/Scrubber for DDRC
//----------------------------

   axi_register_slice DDR_C_TST_AXI4_REG_SLC_1 (
     .aclk           (aclk),
     .aresetn        (slr1_sync_aresetn),

     .s_axi_awid     (ddrc_axi_mstr.awid),
     .s_axi_awaddr   (ddrc_axi_mstr.awaddr),
     .s_axi_awlen    (ddrc_axi_mstr.awlen),
     .s_axi_awsize   (ddrc_axi_mstr.awsize),
     .s_axi_awvalid  (ddrc_axi_mstr.awvalid),
     .s_axi_awready  (ddrc_axi_mstr.awready),
     .s_axi_wdata    (ddrc_axi_mstr.wdata),
     .s_axi_wstrb    (ddrc_axi_mstr.wstrb),
     .s_axi_wlast    (ddrc_axi_mstr.wlast),
     .s_axi_wvalid   (ddrc_axi_mstr.wvalid),
     .s_axi_wready   (ddrc_axi_mstr.wready),
     .s_axi_bid      (ddrc_axi_mstr.bid),
     .s_axi_bresp    (ddrc_axi_mstr.bresp),
     .s_axi_bvalid   (ddrc_axi_mstr.bvalid),
     .s_axi_bready   (ddrc_axi_mstr.bready),
     .s_axi_arid     (ddrc_axi_mstr.arid),
     .s_axi_araddr   (ddrc_axi_mstr.araddr),
     .s_axi_arlen    (ddrc_axi_mstr.arlen),
     .s_axi_arsize   (ddrc_axi_mstr.arsize),
     .s_axi_arvalid  (ddrc_axi_mstr.arvalid),
     .s_axi_arready  (ddrc_axi_mstr.arready),
     .s_axi_rid      (ddrc_axi_mstr.rid),
     .s_axi_rdata    (ddrc_axi_mstr.rdata),
     .s_axi_rresp    (ddrc_axi_mstr.rresp),
     .s_axi_rlast    (ddrc_axi_mstr.rlast),
     .s_axi_rvalid   (ddrc_axi_mstr.rvalid),
     .s_axi_rready   (ddrc_axi_mstr.rready),

     .m_axi_awid     (lcl_cl_sh_ddrc.awid),
     .m_axi_awaddr   (lcl_cl_sh_ddrc.awaddr),
     .m_axi_awlen    (lcl_cl_sh_ddrc.awlen),
     .m_axi_awsize   (lcl_cl_sh_ddrc.awsize),
     .m_axi_awvalid  (lcl_cl_sh_ddrc.awvalid),
     .m_axi_awready  (lcl_cl_sh_ddrc.awready),
     .m_axi_wdata    (lcl_cl_sh_ddrc.wdata),
     .m_axi_wstrb    (lcl_cl_sh_ddrc.wstrb),
     .m_axi_wlast    (lcl_cl_sh_ddrc.wlast),
     .m_axi_wvalid   (lcl_cl_sh_ddrc.wvalid),
     .m_axi_wready   (lcl_cl_sh_ddrc.wready),
     .m_axi_bid      (lcl_cl_sh_ddrc.bid),
     .m_axi_bresp    (lcl_cl_sh_ddrc.bresp),
     .m_axi_bvalid   (lcl_cl_sh_ddrc.bvalid),
     .m_axi_bready   (lcl_cl_sh_ddrc.bready),
     .m_axi_arid     (lcl_cl_sh_ddrc.arid),
     .m_axi_araddr   (lcl_cl_sh_ddrc.araddr),
     .m_axi_arlen    (lcl_cl_sh_ddrc.arlen),
     .m_axi_arsize   (lcl_cl_sh_ddrc.arsize),
     .m_axi_arvalid  (lcl_cl_sh_ddrc.arvalid),
     .m_axi_arready  (lcl_cl_sh_ddrc.arready),
     .m_axi_rid      (lcl_cl_sh_ddrc.rid),
     .m_axi_rdata    (lcl_cl_sh_ddrc.rdata),
     .m_axi_rresp    (lcl_cl_sh_ddrc.rresp),
     .m_axi_rlast    (lcl_cl_sh_ddrc.rlast),
     .m_axi_rvalid   (lcl_cl_sh_ddrc.rvalid),
     .m_axi_rready   (lcl_cl_sh_ddrc.rready)
   );


//----------------------------
// flop the output of interconnect for DDRD
// back to back for SLR crossing
//----------------------------

  //back to back register slices for SLR crossing
   src_register_slice DDR_D_TST_AXI4_REG_SLC_1 (
       .aclk           (aclk),
       .aresetn        (slr1_sync_aresetn),
       .s_axi_awid     (axi_m_48G_64G_.awid),
       .s_axi_awaddr   ({axi_m_48G_64G_.awaddr[63:36], 2'b0, axi_m_48G_64G_.awaddr[33:0]}),
       .s_axi_awlen    (axi_m_48G_64G_.awlen),
       .s_axi_awsize   (axi_m_48G_64G_.awsize),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (axi_m_48G_64G_.awvalid),
       .s_axi_awready  (axi_m_48G_64G_.awready),
       .s_axi_wdata    (axi_m_48G_64G_.wdata),
       .s_axi_wstrb    (axi_m_48G_64G_.wstrb),
       .s_axi_wlast    (axi_m_48G_64G_.wlast),
       .s_axi_wvalid   (axi_m_48G_64G_.wvalid),
       .s_axi_wready   (axi_m_48G_64G_.wready),
       .s_axi_bid      (axi_m_48G_64G_.bid),
       .s_axi_bresp    (axi_m_48G_64G_.bresp),
       .s_axi_bvalid   (axi_m_48G_64G_.bvalid),
       .s_axi_bready   (axi_m_48G_64G_.bready),
       .s_axi_arid     (axi_m_48G_64G_.arid),
       .s_axi_araddr   ({axi_m_48G_64G_.araddr[63:36], 2'b0, axi_m_48G_64G_.araddr[33:0]}),
       .s_axi_arlen    (axi_m_48G_64G_.arlen),
       .s_axi_arsize   (axi_m_48G_64G_.arsize),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (axi_m_48G_64G_.arvalid),
       .s_axi_arready  (axi_m_48G_64G_.arready),
       .s_axi_rid      (axi_m_48G_64G_.rid),
       .s_axi_rdata    (axi_m_48G_64G_.rdata),
       .s_axi_rresp    (axi_m_48G_64G_.rresp),
       .s_axi_rlast    (axi_m_48G_64G_.rlast),
       .s_axi_rvalid   (axi_m_48G_64G_.rvalid),
       .s_axi_rready   (axi_m_48G_64G_.rready),
       .m_axi_awid     (axi_m_48G_64G_2.awid),
       .m_axi_awaddr   (axi_m_48G_64G_2.awaddr),
       .m_axi_awlen    (axi_m_48G_64G_2.awlen),
       .m_axi_awsize   (axi_m_48G_64G_2.awsize),
       .m_axi_awburst  (),
       .m_axi_awlock   (),
       .m_axi_awcache  (),
       .m_axi_awprot   (),
       .m_axi_awregion (),
       .m_axi_awqos    (),
       .m_axi_awvalid  (axi_m_48G_64G_2.awvalid),
       .m_axi_awready  (axi_m_48G_64G_2.awready),
       .m_axi_wdata    (axi_m_48G_64G_2.wdata),
       .m_axi_wstrb    (axi_m_48G_64G_2.wstrb),
       .m_axi_wlast    (axi_m_48G_64G_2.wlast),
       .m_axi_wvalid   (axi_m_48G_64G_2.wvalid),
       .m_axi_wready   (axi_m_48G_64G_2.wready),
       .m_axi_bid      (axi_m_48G_64G_2.bid),
       .m_axi_bresp    (axi_m_48G_64G_2.bresp),
       .m_axi_bvalid   (axi_m_48G_64G_2.bvalid),
       .m_axi_bready   (axi_m_48G_64G_2.bready),
       .m_axi_arid     (axi_m_48G_64G_2.arid),
       .m_axi_araddr   (axi_m_48G_64G_2.araddr),
       .m_axi_arlen    (axi_m_48G_64G_2.arlen),
       .m_axi_arsize   (axi_m_48G_64G_2.arsize),
       .m_axi_arburst  (),
       .m_axi_arlock   (),
       .m_axi_arcache  (),
       .m_axi_arprot   (),
       .m_axi_arregion (),
       .m_axi_arqos    (),
       .m_axi_arvalid  (axi_m_48G_64G_2.arvalid),
       .m_axi_arready  (axi_m_48G_64G_2.arready),
       .m_axi_rid      (axi_m_48G_64G_2.rid),
       .m_axi_rdata    (axi_m_48G_64G_2.rdata),
       .m_axi_rresp    (axi_m_48G_64G_2.rresp),
       .m_axi_rlast    (axi_m_48G_64G_2.rlast),
       .m_axi_rvalid   (axi_m_48G_64G_2.rvalid),
       .m_axi_rready   (axi_m_48G_64G_2.rready)
       );
   dest_register_slice DDR_D_TST_AXI4_REG_SLC_2 (
       .aclk           (aclk),
       .aresetn        (slr0_sync_aresetn),
       .s_axi_awid     (axi_m_48G_64G_2.awid),
       .s_axi_awaddr   (axi_m_48G_64G_2.awaddr),
       .s_axi_awlen    (axi_m_48G_64G_2.awlen),
       .s_axi_awsize   (axi_m_48G_64G_2.awsize),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (axi_m_48G_64G_2.awvalid),
       .s_axi_awready  (axi_m_48G_64G_2.awready),
       .s_axi_wdata    (axi_m_48G_64G_2.wdata),
       .s_axi_wstrb    (axi_m_48G_64G_2.wstrb),
       .s_axi_wlast    (axi_m_48G_64G_2.wlast),
       .s_axi_wvalid   (axi_m_48G_64G_2.wvalid),
       .s_axi_wready   (axi_m_48G_64G_2.wready),
       .s_axi_bid      (axi_m_48G_64G_2.bid),
       .s_axi_bresp    (axi_m_48G_64G_2.bresp),
       .s_axi_bvalid   (axi_m_48G_64G_2.bvalid),
       .s_axi_bready   (axi_m_48G_64G_2.bready),
       .s_axi_arid     (axi_m_48G_64G_2.arid),
       .s_axi_araddr   (axi_m_48G_64G_2.araddr),
       .s_axi_arlen    (axi_m_48G_64G_2.arlen),
       .s_axi_arsize   (axi_m_48G_64G_2.arsize),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (axi_m_48G_64G_2.arvalid),
       .s_axi_arready  (axi_m_48G_64G_2.arready),
       .s_axi_rid      (axi_m_48G_64G_2.rid),
       .s_axi_rdata    (axi_m_48G_64G_2.rdata),
       .s_axi_rresp    (axi_m_48G_64G_2.rresp),
       .s_axi_rlast    (axi_m_48G_64G_2.rlast),
       .s_axi_rvalid   (axi_m_48G_64G_2.rvalid),
       .s_axi_rready   (axi_m_48G_64G_2.rready),
       .m_axi_awid     (axi_m_48G_64G_out.awid),
       .m_axi_awaddr   (axi_m_48G_64G_out.awaddr),
       .m_axi_awlen    (axi_m_48G_64G_out.awlen),
       .m_axi_awsize   (axi_m_48G_64G_out.awsize),
       .m_axi_awburst  (),
       .m_axi_awlock   (),
       .m_axi_awcache  (),
       .m_axi_awprot   (),
       .m_axi_awregion (),
       .m_axi_awqos    (),
       .m_axi_awvalid  (axi_m_48G_64G_out.awvalid),
       .m_axi_awready  (axi_m_48G_64G_out.awready),
       .m_axi_wdata    (axi_m_48G_64G_out.wdata),
       .m_axi_wstrb    (axi_m_48G_64G_out.wstrb),
       .m_axi_wlast    (axi_m_48G_64G_out.wlast),
       .m_axi_wvalid   (axi_m_48G_64G_out.wvalid),
       .m_axi_wready   (axi_m_48G_64G_out.wready),
       .m_axi_bid      (axi_m_48G_64G_out.bid),
       .m_axi_bresp    (axi_m_48G_64G_out.bresp),
       .m_axi_bvalid   (axi_m_48G_64G_out.bvalid),
       .m_axi_bready   (axi_m_48G_64G_out.bready),
       .m_axi_arid     (axi_m_48G_64G_out.arid),
       .m_axi_araddr   (axi_m_48G_64G_out.araddr),
       .m_axi_arlen    (axi_m_48G_64G_out.arlen),
       .m_axi_arsize   (axi_m_48G_64G_out.arsize),
       .m_axi_arburst  (),
       .m_axi_arlock   (),
       .m_axi_arcache  (),
       .m_axi_arprot   (),
       .m_axi_arregion (),
       .m_axi_arqos    (),
       .m_axi_arvalid  (axi_m_48G_64G_out.arvalid),
       .m_axi_arready  (axi_m_48G_64G_out.arready),
       .m_axi_rid      (axi_m_48G_64G_out.rid),
       .m_axi_rdata    (axi_m_48G_64G_out.rdata),
       .m_axi_rresp    (axi_m_48G_64G_out.rresp),
       .m_axi_rlast    (axi_m_48G_64G_out.rlast),
       .m_axi_rvalid   (axi_m_48G_64G_out.rvalid),
       .m_axi_rready   (axi_m_48G_64G_out.rready)
       );

//----------------------------
// ATG/scrubber for DDRD
//----------------------------
   lib_pipe #(.WIDTH(32+32+1+1), .STAGES(NUM_CFG_STGS_CL_DDR_ATG)) PIPE_CFG_REQ_DDR_D (.clk (aclk),
                                                              .rst_n (aresetn),
                                                              .in_bus({ddrd_tst_cfg_bus.addr, ddrd_tst_cfg_bus.wdata, ddrd_tst_cfg_bus.wr, ddrd_tst_cfg_bus.rd}),
                                                              .out_bus({ddrd_tst_cfg_bus_q.addr, ddrd_tst_cfg_bus_q.wdata, ddrd_tst_cfg_bus_q.wr, ddrd_tst_cfg_bus_q.rd})
                                                              );

   lib_pipe #(.WIDTH(32+1), .STAGES(NUM_CFG_STGS_CL_DDR_ATG)) PIPE_CFG_ACK_DDR_D (.clk (aclk),
                                                              .rst_n (aresetn),
                                                              .in_bus({ddrd_tst_cfg_bus_q.ack, ddrd_tst_cfg_bus_q.rdata}),
                                                              .out_bus({ddrd_tst_cfg_bus.ack, ddrd_tst_cfg_bus.rdata})
                                                              );


   lib_pipe #(.WIDTH(2+3+64), .STAGES(NUM_CFG_STGS_CL_DDR_ATG)) PIPE_SCRB_DDR_D (.clk(aclk),
                                                              .rst_n(aresetn),
                                                              .in_bus({ddrd_scrb_bus.enable, ddrd_scrb_bus_q.done, ddrd_scrb_bus_q.state, ddrd_scrb_bus_q.addr}),
                                                              .out_bus({ddrd_scrb_bus_q.enable, ddrd_scrb_bus.done, ddrd_scrb_bus.state, ddrd_scrb_bus.addr})
                                                              );

   cl_tst_scrb #(.DATA_WIDTH(512),
                    .SCRB_BURST_LEN_MINUS1(SCRB_BURST_LEN_MINUS1),
                    .SCRB_MAX_ADDR(SCRB_MAX_ADDR),
                    .NO_SCRB_INST(NO_SCRB_INST)) CL_TST_DDR_D (

         .clk(aclk),
         .rst_n(slr0_sync_aresetn),

         .cfg_addr(ddrd_tst_cfg_bus_q.addr),
         .cfg_wdata(ddrd_tst_cfg_bus_q.wdata),
         .cfg_wr(ddrd_tst_cfg_bus_q.wr),
         .cfg_rd(ddrd_tst_cfg_bus_q.rd),
         .tst_cfg_ack(ddrd_tst_cfg_bus_q.ack),
         .tst_cfg_rdata(ddrd_tst_cfg_bus_q.rdata),

         .slv_awid(ddrd_axi_slv.awid[6:0]),
         .slv_awaddr(ddrd_axi_slv.awaddr),
         .slv_awlen(ddrd_axi_slv.awlen),
         .slv_awsize(ddrd_axi_slv.awsize),
         .slv_awvalid(ddrd_axi_slv.awvalid),
         .slv_awuser(11'b0),
         .slv_awready(ddrd_axi_slv.awready),

         .slv_wid(7'b0),
         .slv_wdata(ddrd_axi_slv.wdata),
         .slv_wstrb(ddrd_axi_slv.wstrb),
         .slv_wlast(ddrd_axi_slv.wlast),
         .slv_wvalid(ddrd_axi_slv.wvalid),
         .slv_wready(ddrd_axi_slv.wready),

         .slv_bid(ddrd_axi_slv.bid[6:0]),
         .slv_bresp(ddrd_axi_slv.bresp),
         .slv_buser(),
         .slv_bvalid(ddrd_axi_slv.bvalid),
         .slv_bready(ddrd_axi_slv.bready),

         .slv_arid(ddrd_axi_slv.arid[6:0]),
         .slv_araddr(ddrd_axi_slv.araddr),
         .slv_arlen(ddrd_axi_slv.arlen),
         .slv_arsize(ddrd_axi_slv.arsize),
         .slv_arvalid(ddrd_axi_slv.arvalid),
         .slv_aruser(11'b0),
         .slv_arready(ddrd_axi_slv.arready),

         .slv_rid(ddrd_axi_slv.rid[6:0]),
         .slv_rdata(ddrd_axi_slv.rdata),
         .slv_rresp(ddrd_axi_slv.rresp),
         .slv_rlast(ddrd_axi_slv.rlast),
         .slv_ruser(),
         .slv_rvalid(ddrd_axi_slv.rvalid),
         .slv_rready(ddrd_axi_slv.rready),

         .awid(lcl_cl_sh_ddrd.awid[8:0]),
         .awaddr(lcl_cl_sh_ddrd.awaddr),
         .awlen(lcl_cl_sh_ddrd.awlen),
         .awvalid(lcl_cl_sh_ddrd.awvalid),
         .awsize(lcl_cl_sh_ddrd.awsize),
         .awuser(),
         .awready(lcl_cl_sh_ddrd.awready),

         .wid(lcl_cl_sh_ddrd.wid[8:0]),
         .wdata(lcl_cl_sh_ddrd.wdata),
         .wstrb(lcl_cl_sh_ddrd.wstrb),
         .wlast(lcl_cl_sh_ddrd.wlast),
         .wvalid(lcl_cl_sh_ddrd.wvalid),
         .wready(lcl_cl_sh_ddrd.wready),

         .bid(lcl_cl_sh_ddrd.bid[8:0]),
         .bresp(lcl_cl_sh_ddrd.bresp),
         .buser(18'h0),
         .bvalid(lcl_cl_sh_ddrd.bvalid),
         .bready(lcl_cl_sh_ddrd.bready),

         .arid(lcl_cl_sh_ddrd.arid[8:0]),
         .araddr(lcl_cl_sh_ddrd.araddr),
         .arlen(lcl_cl_sh_ddrd.arlen),
         .arsize(lcl_cl_sh_ddrd.arsize),
         .arvalid(lcl_cl_sh_ddrd.arvalid),
         .aruser(),
         .arready(lcl_cl_sh_ddrd.arready),

         .rid(lcl_cl_sh_ddrd.rid[8:0]),
         .rdata(lcl_cl_sh_ddrd.rdata),
         .rresp(lcl_cl_sh_ddrd.rresp),
         .rlast(lcl_cl_sh_ddrd.rlast),
         .ruser(18'h0),
         .rvalid(lcl_cl_sh_ddrd.rvalid),
         .rready(lcl_cl_sh_ddrd.rready),

         .scrb_enable(ddrd_scrb_bus_q.enable),
         .scrb_done  (ddrd_scrb_bus_q.done),

         .scrb_dbg_state(ddrd_scrb_bus_q.state),
         .scrb_dbg_addr (ddrd_scrb_bus_q.addr)
      );
      assign lcl_cl_sh_ddrd.awid[15:9] = 7'b0;
      assign lcl_cl_sh_ddrd.wid[15:9] = 7'b0;
      assign lcl_cl_sh_ddrd.arid[15:9] = 7'b0;


endmodule

