module BranchUnit(
  input  [4:0]  io_dinst_rd_bits,
  input  [25:0] io_dinst_imm,
  input         io_dinst_is32bit,
  input  [4:0]  io_dinst_itype,
  input  [3:0]  io_dinst_op,
  input  [63:0] io_rVal1,
  input  [63:0] io_rVal2,
  input         io_cond,
  input  [63:0] io_pc,
  output        io_binst_valid,
  output [63:0] io_binst_bits_pc,
  output        io_binst_bits_unalignedExcp,
  output        io_pcrel_valid,
  output [4:0]  io_pcrel_bits_rd,
  output [63:0] io_pcrel_bits_res
);
  wire [27:0] immS2; // @[Cat.scala 29:58]
  wire [15:0] _T_2; // @[Branch.scala 39:40]
  wire [63:0] imm14S2; // @[Branch.scala 39:50]
  wire [27:0] _T_5; // @[Branch.scala 40:40]
  wire [63:0] imm26S2; // @[Branch.scala 40:50]
  wire [20:0] _T_8; // @[Branch.scala 41:40]
  wire [63:0] imm19S2; // @[Branch.scala 41:50]
  wire [20:0] _T_11; // @[Branch.scala 42:45]
  wire [63:0] imm21S0; // @[Branch.scala 42:55]
  wire [32:0] _T_15; // @[Branch.scala 43:62]
  wire [63:0] imm21S12; // @[Branch.scala 43:72]
  wire  _T_17; // @[Branch.scala 49:52]
  wire [63:0] _T_18; // @[Branch.scala 49:39]
  wire  _T_19; // @[Mux.scala 80:60]
  wire [63:0] _T_20; // @[Mux.scala 80:57]
  wire  _T_21; // @[Mux.scala 80:60]
  wire [63:0] _T_22; // @[Mux.scala 80:57]
  wire  _T_23; // @[Mux.scala 80:60]
  wire [63:0] _T_24; // @[Mux.scala 80:57]
  wire  _T_25; // @[Mux.scala 80:60]
  wire [63:0] _T_26; // @[Mux.scala 80:57]
  wire  _T_27; // @[Mux.scala 80:60]
  wire [63:0] immSExt; // @[Mux.scala 80:57]
  wire  _T_28; // @[Branch.scala 53:23]
  wire  _T_30; // @[Branch.scala 53:35]
  wire [63:0] _T_32; // @[Cat.scala 29:58]
  wire [63:0] pc; // @[Branch.scala 53:63]
  wire [64:0] _T_33; // @[Branch.scala 56:28]
  wire [64:0] _GEN_7; // @[Branch.scala 56:33]
  wire [64:0] pcadd; // @[Branch.scala 56:44]
  wire  _T_38; // @[Branch.scala 59:30]
  wire [5:0] bit_pos; // @[Cat.scala 29:58]
  wire  _T_41; // @[Branch.scala 62:32]
  wire [64:0] bpc; // @[Branch.scala 62:16]
  wire [63:0] _T_44; // @[Branch.scala 72:27]
  wire [3:0] _GEN_8; // @[Branch.scala 72:37]
  wire  _T_46; // @[Branch.scala 72:37]
  wire  _T_48; // @[Branch.scala 74:57]
  wire  _T_49; // @[Branch.scala 74:75]
  wire  _T_50; // @[Branch.scala 74:23]
  wire  _T_52; // @[Branch.scala 75:57]
  wire  _T_53; // @[Branch.scala 75:75]
  wire  _T_54; // @[Branch.scala 75:23]
  wire  _T_55; // @[Mux.scala 80:60]
  wire  _T_56; // @[Mux.scala 80:57]
  wire  _T_57; // @[Mux.scala 80:60]
  wire  _T_58; // @[Mux.scala 80:57]
  wire  _T_61; // @[Mux.scala 80:60]
  wire  _T_62; // @[Mux.scala 80:57]
  wire  _T_64; // @[Mux.scala 80:57]
  wire  _T_66; // @[Mux.scala 80:57]
  wire  _T_69; // @[Branch.scala 83:23]
  wire  _T_71; // @[Branch.scala 83:34]
  wire  _T_74; // @[Branch.scala 84:31]
  wire  _T_75; // @[Branch.scala 83:59]
  wire [63:0] _T_77; // @[Branch.scala 86:24]
  wire [64:0] _GEN_5; // @[Branch.scala 84:58]
  assign immS2 = {io_dinst_imm,2'h0}; // @[Cat.scala 29:58]
  assign _T_2 = immS2[15:0]; // @[Branch.scala 39:40]
  assign imm14S2 = {{48{_T_2[15]}},_T_2}; // @[Branch.scala 39:50]
  assign _T_5 = {io_dinst_imm,2'h0}; // @[Branch.scala 40:40]
  assign imm26S2 = {{36{_T_5[27]}},_T_5}; // @[Branch.scala 40:50]
  assign _T_8 = immS2[20:0]; // @[Branch.scala 41:40]
  assign imm19S2 = {{43{_T_8[20]}},_T_8}; // @[Branch.scala 41:50]
  assign _T_11 = io_dinst_imm[20:0]; // @[Branch.scala 42:45]
  assign imm21S0 = {{43{_T_11[20]}},_T_11}; // @[Branch.scala 42:55]
  assign _T_15 = {io_dinst_imm[20:0],12'h0}; // @[Branch.scala 43:62]
  assign imm21S12 = {{31{_T_15[32]}},_T_15}; // @[Branch.scala 43:72]
  assign _T_17 = io_dinst_op == 4'h1; // @[Branch.scala 49:52]
  assign _T_18 = _T_17 ? $signed(imm21S12) : $signed(imm21S0); // @[Branch.scala 49:39]
  assign _T_19 = 5'h18 == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_20 = _T_19 ? $signed(imm26S2) : $signed(imm21S0); // @[Mux.scala 80:57]
  assign _T_21 = 5'h19 == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_22 = _T_21 ? $signed(imm19S2) : $signed(_T_20); // @[Mux.scala 80:57]
  assign _T_23 = 5'h1b == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_24 = _T_23 ? $signed(imm19S2) : $signed(_T_22); // @[Mux.scala 80:57]
  assign _T_25 = 5'h1a == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_26 = _T_25 ? $signed(imm14S2) : $signed(_T_24); // @[Mux.scala 80:57]
  assign _T_27 = 5'h3 == io_dinst_itype; // @[Mux.scala 80:60]
  assign immSExt = _T_27 ? $signed(_T_18) : $signed(_T_26); // @[Mux.scala 80:57]
  assign _T_28 = io_dinst_itype == 5'h3; // @[Branch.scala 53:23]
  assign _T_30 = _T_28 & _T_17; // @[Branch.scala 53:35]
  assign _T_32 = {io_pc[63:12],12'h0}; // @[Cat.scala 29:58]
  assign pc = _T_30 ? _T_32 : io_pc; // @[Branch.scala 53:63]
  assign _T_33 = {1'b0,$signed(pc)}; // @[Branch.scala 56:28]
  assign _GEN_7 = {{1{immSExt[63]}},immSExt}; // @[Branch.scala 56:33]
  assign pcadd = $signed(_T_33) + $signed(_GEN_7); // @[Branch.scala 56:44]
  assign _T_38 = ~io_dinst_is32bit; // @[Branch.scala 59:30]
  assign bit_pos = {_T_38,io_dinst_imm[18:14]}; // @[Cat.scala 29:58]
  assign _T_41 = io_dinst_itype == 5'h1c; // @[Branch.scala 62:32]
  assign bpc = _T_41 ? {{1'd0}, io_rVal1} : pcadd; // @[Branch.scala 62:16]
  assign _T_44 = io_rVal2 >> bit_pos; // @[Branch.scala 72:27]
  assign _GEN_8 = {{3'd0}, _T_44[0]}; // @[Branch.scala 72:37]
  assign _T_46 = _GEN_8 == io_dinst_op; // @[Branch.scala 72:37]
  assign _T_48 = io_rVal2[31:0] == 32'h0; // @[Branch.scala 74:57]
  assign _T_49 = io_rVal2 == 64'h0; // @[Branch.scala 74:75]
  assign _T_50 = io_dinst_is32bit ? _T_48 : _T_49; // @[Branch.scala 74:23]
  assign _T_52 = io_rVal2[31:0] != 32'h0; // @[Branch.scala 75:57]
  assign _T_53 = io_rVal2 != 64'h0; // @[Branch.scala 75:75]
  assign _T_54 = io_dinst_is32bit ? _T_52 : _T_53; // @[Branch.scala 75:23]
  assign _T_55 = 4'h0 == io_dinst_op; // @[Mux.scala 80:60]
  assign _T_56 = _T_55 & _T_50; // @[Mux.scala 80:57]
  assign _T_57 = 4'h1 == io_dinst_op; // @[Mux.scala 80:60]
  assign _T_58 = _T_57 ? _T_54 : _T_56; // @[Mux.scala 80:57]
  assign _T_61 = 5'h1c == io_dinst_itype; // @[Mux.scala 80:60]
  assign _T_62 = _T_61 | _T_19; // @[Mux.scala 80:57]
  assign _T_64 = _T_21 ? io_cond : _T_62; // @[Mux.scala 80:57]
  assign _T_66 = _T_25 ? _T_46 : _T_64; // @[Mux.scala 80:57]
  assign _T_69 = io_dinst_itype == 5'h18; // @[Branch.scala 83:23]
  assign _T_71 = _T_69 & _T_17; // @[Branch.scala 83:34]
  assign _T_74 = _T_41 & _T_17; // @[Branch.scala 84:31]
  assign _T_75 = _T_71 | _T_74; // @[Branch.scala 83:59]
  assign _T_77 = io_pc + 64'h4; // @[Branch.scala 86:24]
  assign _GEN_5 = _T_75 ? {{1'd0}, _T_77} : pcadd; // @[Branch.scala 84:58]
  assign io_binst_valid = _T_23 ? _T_58 : _T_66; // @[Branch.scala 67:18]
  assign io_binst_bits_pc = bpc[63:0]; // @[Branch.scala 66:17]
  assign io_binst_bits_unalignedExcp = bpc[1:0] != 2'h0; // @[Branch.scala 66:17]
  assign io_pcrel_valid = _T_75 | _T_28; // @[Branch.scala 82:18 Branch.scala 87:20 Branch.scala 91:20]
  assign io_pcrel_bits_rd = _T_75 ? 5'h1e : io_dinst_rd_bits; // @[Branch.scala 93:17]
  assign io_pcrel_bits_res = _GEN_5[63:0]; // @[Branch.scala 93:17]
endmodule
