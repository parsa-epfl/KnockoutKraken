module PseudoBitmapLRU(
  input        clock,
  input        reset,
  input        io_idx_1_valid,
  input  [5:0] io_idx_1_bits,
  input        io_idx_2_valid,
  input  [5:0] io_idx_2_bits,
  output [5:0] io_lru_idx
);
  reg  bitmap_0; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_0;
  reg  bitmap_1; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_1;
  reg  bitmap_2; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_2;
  reg  bitmap_3; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_3;
  reg  bitmap_4; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_4;
  reg  bitmap_5; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_5;
  reg  bitmap_6; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_6;
  reg  bitmap_7; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_7;
  reg  bitmap_8; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_8;
  reg  bitmap_9; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_9;
  reg  bitmap_10; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_10;
  reg  bitmap_11; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_11;
  reg  bitmap_12; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_12;
  reg  bitmap_13; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_13;
  reg  bitmap_14; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_14;
  reg  bitmap_15; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_15;
  reg  bitmap_16; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_16;
  reg  bitmap_17; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_17;
  reg  bitmap_18; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_18;
  reg  bitmap_19; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_19;
  reg  bitmap_20; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_20;
  reg  bitmap_21; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_21;
  reg  bitmap_22; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_22;
  reg  bitmap_23; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_23;
  reg  bitmap_24; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_24;
  reg  bitmap_25; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_25;
  reg  bitmap_26; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_26;
  reg  bitmap_27; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_27;
  reg  bitmap_28; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_28;
  reg  bitmap_29; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_29;
  reg  bitmap_30; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_30;
  reg  bitmap_31; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_31;
  reg  bitmap_32; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_32;
  reg  bitmap_33; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_33;
  reg  bitmap_34; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_34;
  reg  bitmap_35; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_35;
  reg  bitmap_36; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_36;
  reg  bitmap_37; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_37;
  reg  bitmap_38; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_38;
  reg  bitmap_39; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_39;
  reg  bitmap_40; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_40;
  reg  bitmap_41; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_41;
  reg  bitmap_42; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_42;
  reg  bitmap_43; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_43;
  reg  bitmap_44; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_44;
  reg  bitmap_45; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_45;
  reg  bitmap_46; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_46;
  reg  bitmap_47; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_47;
  reg  bitmap_48; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_48;
  reg  bitmap_49; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_49;
  reg  bitmap_50; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_50;
  reg  bitmap_51; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_51;
  reg  bitmap_52; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_52;
  reg  bitmap_53; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_53;
  reg  bitmap_54; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_54;
  reg  bitmap_55; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_55;
  reg  bitmap_56; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_56;
  reg  bitmap_57; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_57;
  reg  bitmap_58; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_58;
  reg  bitmap_59; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_59;
  reg  bitmap_60; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_60;
  reg  bitmap_61; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_61;
  reg  bitmap_62; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_62;
  reg  bitmap_63; // @[ReplacementPolicy.scala 78:23]
  reg [31:0] _RAND_63;
  wire  _GEN_320; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_0; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_321; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_1; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_322; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_2; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_323; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_3; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_324; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_4; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_325; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_5; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_326; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_6; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_327; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_7; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_328; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_8; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_329; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_9; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_330; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_10; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_331; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_11; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_332; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_12; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_333; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_13; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_334; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_14; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_335; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_15; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_336; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_16; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_337; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_17; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_338; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_18; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_339; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_19; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_340; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_20; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_341; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_21; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_342; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_22; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_343; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_23; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_344; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_24; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_345; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_25; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_346; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_26; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_347; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_27; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_348; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_28; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_349; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_29; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_350; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_30; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_351; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_31; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_352; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_32; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_353; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_33; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_354; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_34; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_355; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_35; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_356; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_36; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_357; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_37; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_358; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_38; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_359; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_39; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_360; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_40; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_361; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_41; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_362; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_42; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_363; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_43; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_364; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_44; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_365; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_45; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_366; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_46; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_367; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_47; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_368; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_48; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_369; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_49; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_370; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_50; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_371; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_51; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_372; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_52; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_373; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_53; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_374; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_54; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_375; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_55; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_376; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_56; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_377; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_57; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_378; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_58; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_379; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_59; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_380; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_60; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_381; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_61; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_382; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_62; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_383; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_63; // @[ReplacementPolicy.scala 80:27]
  wire  _GEN_64; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_65; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_66; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_67; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_68; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_69; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_70; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_71; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_72; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_73; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_74; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_75; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_76; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_77; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_78; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_79; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_80; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_81; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_82; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_83; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_84; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_85; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_86; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_87; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_88; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_89; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_90; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_91; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_92; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_93; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_94; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_95; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_96; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_97; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_98; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_99; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_100; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_101; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_102; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_103; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_104; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_105; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_106; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_107; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_108; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_109; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_110; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_111; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_112; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_113; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_114; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_115; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_116; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_117; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_118; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_119; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_120; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_121; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_122; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_123; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_124; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_125; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_126; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_127; // @[ReplacementPolicy.scala 79:24]
  wire  _GEN_384; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_128; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_385; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_129; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_386; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_130; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_387; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_131; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_388; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_132; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_389; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_133; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_390; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_134; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_391; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_135; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_392; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_136; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_393; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_137; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_394; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_138; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_395; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_139; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_396; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_140; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_397; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_141; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_398; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_142; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_399; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_143; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_400; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_144; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_401; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_145; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_402; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_146; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_403; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_147; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_404; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_148; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_405; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_149; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_406; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_150; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_407; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_151; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_408; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_152; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_409; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_153; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_410; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_154; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_411; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_155; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_412; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_156; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_413; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_157; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_414; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_158; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_415; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_159; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_416; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_160; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_417; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_161; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_418; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_162; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_419; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_163; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_420; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_164; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_421; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_165; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_422; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_166; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_423; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_167; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_424; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_168; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_425; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_169; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_426; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_170; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_427; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_171; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_428; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_172; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_429; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_173; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_430; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_174; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_431; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_175; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_432; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_176; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_433; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_177; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_434; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_178; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_435; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_179; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_436; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_180; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_437; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_181; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_438; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_182; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_439; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_183; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_440; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_184; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_441; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_185; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_442; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_186; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_443; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_187; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_444; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_188; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_445; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_189; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_446; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_190; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_447; // @[ReplacementPolicy.scala 84:27]
  wire  _GEN_191; // @[ReplacementPolicy.scala 84:27]
  wire [7:0] _T_7; // @[ReplacementPolicy.scala 87:33]
  wire [15:0] _T_15; // @[ReplacementPolicy.scala 87:33]
  wire [7:0] _T_22; // @[ReplacementPolicy.scala 87:33]
  wire [31:0] _T_31; // @[ReplacementPolicy.scala 87:33]
  wire [7:0] _T_38; // @[ReplacementPolicy.scala 87:33]
  wire [15:0] _T_46; // @[ReplacementPolicy.scala 87:33]
  wire [7:0] _T_53; // @[ReplacementPolicy.scala 87:33]
  wire [31:0] _T_62; // @[ReplacementPolicy.scala 87:33]
  wire [63:0] bitmapU; // @[ReplacementPolicy.scala 87:33]
  wire  _T_66; // @[ReplacementPolicy.scala 88:31]
  wire [63:0] bitmapUNeg; // @[ReplacementPolicy.scala 92:47]
  wire [5:0] _T_132; // @[Mux.scala 47:69]
  wire [5:0] _T_133; // @[Mux.scala 47:69]
  wire [5:0] _T_134; // @[Mux.scala 47:69]
  wire [5:0] _T_135; // @[Mux.scala 47:69]
  wire [5:0] _T_136; // @[Mux.scala 47:69]
  wire [5:0] _T_137; // @[Mux.scala 47:69]
  wire [5:0] _T_138; // @[Mux.scala 47:69]
  wire [5:0] _T_139; // @[Mux.scala 47:69]
  wire [5:0] _T_140; // @[Mux.scala 47:69]
  wire [5:0] _T_141; // @[Mux.scala 47:69]
  wire [5:0] _T_142; // @[Mux.scala 47:69]
  wire [5:0] _T_143; // @[Mux.scala 47:69]
  wire [5:0] _T_144; // @[Mux.scala 47:69]
  wire [5:0] _T_145; // @[Mux.scala 47:69]
  wire [5:0] _T_146; // @[Mux.scala 47:69]
  wire [5:0] _T_147; // @[Mux.scala 47:69]
  wire [5:0] _T_148; // @[Mux.scala 47:69]
  wire [5:0] _T_149; // @[Mux.scala 47:69]
  wire [5:0] _T_150; // @[Mux.scala 47:69]
  wire [5:0] _T_151; // @[Mux.scala 47:69]
  wire [5:0] _T_152; // @[Mux.scala 47:69]
  wire [5:0] _T_153; // @[Mux.scala 47:69]
  wire [5:0] _T_154; // @[Mux.scala 47:69]
  wire [5:0] _T_155; // @[Mux.scala 47:69]
  wire [5:0] _T_156; // @[Mux.scala 47:69]
  wire [5:0] _T_157; // @[Mux.scala 47:69]
  wire [5:0] _T_158; // @[Mux.scala 47:69]
  wire [5:0] _T_159; // @[Mux.scala 47:69]
  wire [5:0] _T_160; // @[Mux.scala 47:69]
  wire [5:0] _T_161; // @[Mux.scala 47:69]
  wire [5:0] _T_162; // @[Mux.scala 47:69]
  wire [5:0] _T_163; // @[Mux.scala 47:69]
  wire [5:0] _T_164; // @[Mux.scala 47:69]
  wire [5:0] _T_165; // @[Mux.scala 47:69]
  wire [5:0] _T_166; // @[Mux.scala 47:69]
  wire [5:0] _T_167; // @[Mux.scala 47:69]
  wire [5:0] _T_168; // @[Mux.scala 47:69]
  wire [5:0] _T_169; // @[Mux.scala 47:69]
  wire [5:0] _T_170; // @[Mux.scala 47:69]
  wire [5:0] _T_171; // @[Mux.scala 47:69]
  wire [5:0] _T_172; // @[Mux.scala 47:69]
  wire [5:0] _T_173; // @[Mux.scala 47:69]
  wire [5:0] _T_174; // @[Mux.scala 47:69]
  wire [5:0] _T_175; // @[Mux.scala 47:69]
  wire [5:0] _T_176; // @[Mux.scala 47:69]
  wire [5:0] _T_177; // @[Mux.scala 47:69]
  wire [5:0] _T_178; // @[Mux.scala 47:69]
  wire [5:0] _T_179; // @[Mux.scala 47:69]
  wire [5:0] _T_180; // @[Mux.scala 47:69]
  wire [5:0] _T_181; // @[Mux.scala 47:69]
  wire [5:0] _T_182; // @[Mux.scala 47:69]
  wire [5:0] _T_183; // @[Mux.scala 47:69]
  wire [5:0] _T_184; // @[Mux.scala 47:69]
  wire [5:0] _T_185; // @[Mux.scala 47:69]
  wire [5:0] _T_186; // @[Mux.scala 47:69]
  wire [5:0] _T_187; // @[Mux.scala 47:69]
  wire [5:0] _T_188; // @[Mux.scala 47:69]
  wire [5:0] _T_189; // @[Mux.scala 47:69]
  wire [5:0] _T_190; // @[Mux.scala 47:69]
  wire [5:0] _T_191; // @[Mux.scala 47:69]
  wire [5:0] _T_192; // @[Mux.scala 47:69]
  wire [5:0] _T_193; // @[Mux.scala 47:69]
  assign _GEN_320 = 6'h0 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_0 = _GEN_320 | bitmap_0; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_321 = 6'h1 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_1 = _GEN_321 | bitmap_1; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_322 = 6'h2 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_2 = _GEN_322 | bitmap_2; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_323 = 6'h3 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_3 = _GEN_323 | bitmap_3; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_324 = 6'h4 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_4 = _GEN_324 | bitmap_4; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_325 = 6'h5 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_5 = _GEN_325 | bitmap_5; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_326 = 6'h6 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_6 = _GEN_326 | bitmap_6; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_327 = 6'h7 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_7 = _GEN_327 | bitmap_7; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_328 = 6'h8 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_8 = _GEN_328 | bitmap_8; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_329 = 6'h9 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_9 = _GEN_329 | bitmap_9; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_330 = 6'ha == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_10 = _GEN_330 | bitmap_10; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_331 = 6'hb == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_11 = _GEN_331 | bitmap_11; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_332 = 6'hc == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_12 = _GEN_332 | bitmap_12; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_333 = 6'hd == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_13 = _GEN_333 | bitmap_13; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_334 = 6'he == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_14 = _GEN_334 | bitmap_14; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_335 = 6'hf == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_15 = _GEN_335 | bitmap_15; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_336 = 6'h10 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_16 = _GEN_336 | bitmap_16; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_337 = 6'h11 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_17 = _GEN_337 | bitmap_17; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_338 = 6'h12 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_18 = _GEN_338 | bitmap_18; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_339 = 6'h13 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_19 = _GEN_339 | bitmap_19; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_340 = 6'h14 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_20 = _GEN_340 | bitmap_20; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_341 = 6'h15 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_21 = _GEN_341 | bitmap_21; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_342 = 6'h16 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_22 = _GEN_342 | bitmap_22; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_343 = 6'h17 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_23 = _GEN_343 | bitmap_23; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_344 = 6'h18 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_24 = _GEN_344 | bitmap_24; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_345 = 6'h19 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_25 = _GEN_345 | bitmap_25; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_346 = 6'h1a == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_26 = _GEN_346 | bitmap_26; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_347 = 6'h1b == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_27 = _GEN_347 | bitmap_27; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_348 = 6'h1c == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_28 = _GEN_348 | bitmap_28; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_349 = 6'h1d == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_29 = _GEN_349 | bitmap_29; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_350 = 6'h1e == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_30 = _GEN_350 | bitmap_30; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_351 = 6'h1f == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_31 = _GEN_351 | bitmap_31; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_352 = 6'h20 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_32 = _GEN_352 | bitmap_32; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_353 = 6'h21 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_33 = _GEN_353 | bitmap_33; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_354 = 6'h22 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_34 = _GEN_354 | bitmap_34; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_355 = 6'h23 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_35 = _GEN_355 | bitmap_35; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_356 = 6'h24 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_36 = _GEN_356 | bitmap_36; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_357 = 6'h25 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_37 = _GEN_357 | bitmap_37; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_358 = 6'h26 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_38 = _GEN_358 | bitmap_38; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_359 = 6'h27 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_39 = _GEN_359 | bitmap_39; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_360 = 6'h28 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_40 = _GEN_360 | bitmap_40; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_361 = 6'h29 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_41 = _GEN_361 | bitmap_41; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_362 = 6'h2a == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_42 = _GEN_362 | bitmap_42; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_363 = 6'h2b == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_43 = _GEN_363 | bitmap_43; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_364 = 6'h2c == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_44 = _GEN_364 | bitmap_44; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_365 = 6'h2d == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_45 = _GEN_365 | bitmap_45; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_366 = 6'h2e == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_46 = _GEN_366 | bitmap_46; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_367 = 6'h2f == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_47 = _GEN_367 | bitmap_47; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_368 = 6'h30 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_48 = _GEN_368 | bitmap_48; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_369 = 6'h31 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_49 = _GEN_369 | bitmap_49; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_370 = 6'h32 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_50 = _GEN_370 | bitmap_50; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_371 = 6'h33 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_51 = _GEN_371 | bitmap_51; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_372 = 6'h34 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_52 = _GEN_372 | bitmap_52; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_373 = 6'h35 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_53 = _GEN_373 | bitmap_53; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_374 = 6'h36 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_54 = _GEN_374 | bitmap_54; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_375 = 6'h37 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_55 = _GEN_375 | bitmap_55; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_376 = 6'h38 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_56 = _GEN_376 | bitmap_56; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_377 = 6'h39 == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_57 = _GEN_377 | bitmap_57; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_378 = 6'h3a == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_58 = _GEN_378 | bitmap_58; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_379 = 6'h3b == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_59 = _GEN_379 | bitmap_59; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_380 = 6'h3c == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_60 = _GEN_380 | bitmap_60; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_381 = 6'h3d == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_61 = _GEN_381 | bitmap_61; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_382 = 6'h3e == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_62 = _GEN_382 | bitmap_62; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_383 = 6'h3f == io_idx_1_bits; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_63 = _GEN_383 | bitmap_63; // @[ReplacementPolicy.scala 80:27]
  assign _GEN_64 = io_idx_1_valid ? _GEN_0 : bitmap_0; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_65 = io_idx_1_valid ? _GEN_1 : bitmap_1; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_66 = io_idx_1_valid ? _GEN_2 : bitmap_2; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_67 = io_idx_1_valid ? _GEN_3 : bitmap_3; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_68 = io_idx_1_valid ? _GEN_4 : bitmap_4; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_69 = io_idx_1_valid ? _GEN_5 : bitmap_5; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_70 = io_idx_1_valid ? _GEN_6 : bitmap_6; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_71 = io_idx_1_valid ? _GEN_7 : bitmap_7; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_72 = io_idx_1_valid ? _GEN_8 : bitmap_8; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_73 = io_idx_1_valid ? _GEN_9 : bitmap_9; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_74 = io_idx_1_valid ? _GEN_10 : bitmap_10; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_75 = io_idx_1_valid ? _GEN_11 : bitmap_11; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_76 = io_idx_1_valid ? _GEN_12 : bitmap_12; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_77 = io_idx_1_valid ? _GEN_13 : bitmap_13; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_78 = io_idx_1_valid ? _GEN_14 : bitmap_14; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_79 = io_idx_1_valid ? _GEN_15 : bitmap_15; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_80 = io_idx_1_valid ? _GEN_16 : bitmap_16; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_81 = io_idx_1_valid ? _GEN_17 : bitmap_17; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_82 = io_idx_1_valid ? _GEN_18 : bitmap_18; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_83 = io_idx_1_valid ? _GEN_19 : bitmap_19; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_84 = io_idx_1_valid ? _GEN_20 : bitmap_20; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_85 = io_idx_1_valid ? _GEN_21 : bitmap_21; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_86 = io_idx_1_valid ? _GEN_22 : bitmap_22; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_87 = io_idx_1_valid ? _GEN_23 : bitmap_23; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_88 = io_idx_1_valid ? _GEN_24 : bitmap_24; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_89 = io_idx_1_valid ? _GEN_25 : bitmap_25; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_90 = io_idx_1_valid ? _GEN_26 : bitmap_26; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_91 = io_idx_1_valid ? _GEN_27 : bitmap_27; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_92 = io_idx_1_valid ? _GEN_28 : bitmap_28; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_93 = io_idx_1_valid ? _GEN_29 : bitmap_29; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_94 = io_idx_1_valid ? _GEN_30 : bitmap_30; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_95 = io_idx_1_valid ? _GEN_31 : bitmap_31; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_96 = io_idx_1_valid ? _GEN_32 : bitmap_32; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_97 = io_idx_1_valid ? _GEN_33 : bitmap_33; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_98 = io_idx_1_valid ? _GEN_34 : bitmap_34; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_99 = io_idx_1_valid ? _GEN_35 : bitmap_35; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_100 = io_idx_1_valid ? _GEN_36 : bitmap_36; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_101 = io_idx_1_valid ? _GEN_37 : bitmap_37; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_102 = io_idx_1_valid ? _GEN_38 : bitmap_38; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_103 = io_idx_1_valid ? _GEN_39 : bitmap_39; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_104 = io_idx_1_valid ? _GEN_40 : bitmap_40; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_105 = io_idx_1_valid ? _GEN_41 : bitmap_41; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_106 = io_idx_1_valid ? _GEN_42 : bitmap_42; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_107 = io_idx_1_valid ? _GEN_43 : bitmap_43; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_108 = io_idx_1_valid ? _GEN_44 : bitmap_44; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_109 = io_idx_1_valid ? _GEN_45 : bitmap_45; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_110 = io_idx_1_valid ? _GEN_46 : bitmap_46; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_111 = io_idx_1_valid ? _GEN_47 : bitmap_47; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_112 = io_idx_1_valid ? _GEN_48 : bitmap_48; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_113 = io_idx_1_valid ? _GEN_49 : bitmap_49; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_114 = io_idx_1_valid ? _GEN_50 : bitmap_50; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_115 = io_idx_1_valid ? _GEN_51 : bitmap_51; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_116 = io_idx_1_valid ? _GEN_52 : bitmap_52; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_117 = io_idx_1_valid ? _GEN_53 : bitmap_53; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_118 = io_idx_1_valid ? _GEN_54 : bitmap_54; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_119 = io_idx_1_valid ? _GEN_55 : bitmap_55; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_120 = io_idx_1_valid ? _GEN_56 : bitmap_56; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_121 = io_idx_1_valid ? _GEN_57 : bitmap_57; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_122 = io_idx_1_valid ? _GEN_58 : bitmap_58; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_123 = io_idx_1_valid ? _GEN_59 : bitmap_59; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_124 = io_idx_1_valid ? _GEN_60 : bitmap_60; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_125 = io_idx_1_valid ? _GEN_61 : bitmap_61; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_126 = io_idx_1_valid ? _GEN_62 : bitmap_62; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_127 = io_idx_1_valid ? _GEN_63 : bitmap_63; // @[ReplacementPolicy.scala 79:24]
  assign _GEN_384 = 6'h0 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_128 = _GEN_384 | _GEN_64; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_385 = 6'h1 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_129 = _GEN_385 | _GEN_65; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_386 = 6'h2 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_130 = _GEN_386 | _GEN_66; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_387 = 6'h3 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_131 = _GEN_387 | _GEN_67; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_388 = 6'h4 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_132 = _GEN_388 | _GEN_68; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_389 = 6'h5 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_133 = _GEN_389 | _GEN_69; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_390 = 6'h6 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_134 = _GEN_390 | _GEN_70; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_391 = 6'h7 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_135 = _GEN_391 | _GEN_71; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_392 = 6'h8 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_136 = _GEN_392 | _GEN_72; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_393 = 6'h9 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_137 = _GEN_393 | _GEN_73; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_394 = 6'ha == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_138 = _GEN_394 | _GEN_74; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_395 = 6'hb == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_139 = _GEN_395 | _GEN_75; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_396 = 6'hc == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_140 = _GEN_396 | _GEN_76; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_397 = 6'hd == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_141 = _GEN_397 | _GEN_77; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_398 = 6'he == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_142 = _GEN_398 | _GEN_78; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_399 = 6'hf == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_143 = _GEN_399 | _GEN_79; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_400 = 6'h10 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_144 = _GEN_400 | _GEN_80; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_401 = 6'h11 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_145 = _GEN_401 | _GEN_81; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_402 = 6'h12 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_146 = _GEN_402 | _GEN_82; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_403 = 6'h13 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_147 = _GEN_403 | _GEN_83; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_404 = 6'h14 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_148 = _GEN_404 | _GEN_84; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_405 = 6'h15 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_149 = _GEN_405 | _GEN_85; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_406 = 6'h16 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_150 = _GEN_406 | _GEN_86; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_407 = 6'h17 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_151 = _GEN_407 | _GEN_87; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_408 = 6'h18 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_152 = _GEN_408 | _GEN_88; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_409 = 6'h19 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_153 = _GEN_409 | _GEN_89; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_410 = 6'h1a == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_154 = _GEN_410 | _GEN_90; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_411 = 6'h1b == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_155 = _GEN_411 | _GEN_91; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_412 = 6'h1c == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_156 = _GEN_412 | _GEN_92; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_413 = 6'h1d == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_157 = _GEN_413 | _GEN_93; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_414 = 6'h1e == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_158 = _GEN_414 | _GEN_94; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_415 = 6'h1f == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_159 = _GEN_415 | _GEN_95; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_416 = 6'h20 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_160 = _GEN_416 | _GEN_96; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_417 = 6'h21 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_161 = _GEN_417 | _GEN_97; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_418 = 6'h22 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_162 = _GEN_418 | _GEN_98; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_419 = 6'h23 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_163 = _GEN_419 | _GEN_99; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_420 = 6'h24 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_164 = _GEN_420 | _GEN_100; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_421 = 6'h25 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_165 = _GEN_421 | _GEN_101; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_422 = 6'h26 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_166 = _GEN_422 | _GEN_102; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_423 = 6'h27 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_167 = _GEN_423 | _GEN_103; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_424 = 6'h28 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_168 = _GEN_424 | _GEN_104; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_425 = 6'h29 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_169 = _GEN_425 | _GEN_105; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_426 = 6'h2a == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_170 = _GEN_426 | _GEN_106; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_427 = 6'h2b == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_171 = _GEN_427 | _GEN_107; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_428 = 6'h2c == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_172 = _GEN_428 | _GEN_108; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_429 = 6'h2d == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_173 = _GEN_429 | _GEN_109; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_430 = 6'h2e == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_174 = _GEN_430 | _GEN_110; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_431 = 6'h2f == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_175 = _GEN_431 | _GEN_111; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_432 = 6'h30 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_176 = _GEN_432 | _GEN_112; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_433 = 6'h31 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_177 = _GEN_433 | _GEN_113; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_434 = 6'h32 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_178 = _GEN_434 | _GEN_114; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_435 = 6'h33 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_179 = _GEN_435 | _GEN_115; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_436 = 6'h34 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_180 = _GEN_436 | _GEN_116; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_437 = 6'h35 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_181 = _GEN_437 | _GEN_117; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_438 = 6'h36 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_182 = _GEN_438 | _GEN_118; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_439 = 6'h37 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_183 = _GEN_439 | _GEN_119; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_440 = 6'h38 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_184 = _GEN_440 | _GEN_120; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_441 = 6'h39 == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_185 = _GEN_441 | _GEN_121; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_442 = 6'h3a == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_186 = _GEN_442 | _GEN_122; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_443 = 6'h3b == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_187 = _GEN_443 | _GEN_123; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_444 = 6'h3c == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_188 = _GEN_444 | _GEN_124; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_445 = 6'h3d == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_189 = _GEN_445 | _GEN_125; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_446 = 6'h3e == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_190 = _GEN_446 | _GEN_126; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_447 = 6'h3f == io_idx_2_bits; // @[ReplacementPolicy.scala 84:27]
  assign _GEN_191 = _GEN_447 | _GEN_127; // @[ReplacementPolicy.scala 84:27]
  assign _T_7 = {bitmap_7,bitmap_6,bitmap_5,bitmap_4,bitmap_3,bitmap_2,bitmap_1,bitmap_0}; // @[ReplacementPolicy.scala 87:33]
  assign _T_15 = {bitmap_15,bitmap_14,bitmap_13,bitmap_12,bitmap_11,bitmap_10,bitmap_9,bitmap_8,_T_7}; // @[ReplacementPolicy.scala 87:33]
  assign _T_22 = {bitmap_23,bitmap_22,bitmap_21,bitmap_20,bitmap_19,bitmap_18,bitmap_17,bitmap_16}; // @[ReplacementPolicy.scala 87:33]
  assign _T_31 = {bitmap_31,bitmap_30,bitmap_29,bitmap_28,bitmap_27,bitmap_26,bitmap_25,bitmap_24,_T_22,_T_15}; // @[ReplacementPolicy.scala 87:33]
  assign _T_38 = {bitmap_39,bitmap_38,bitmap_37,bitmap_36,bitmap_35,bitmap_34,bitmap_33,bitmap_32}; // @[ReplacementPolicy.scala 87:33]
  assign _T_46 = {bitmap_47,bitmap_46,bitmap_45,bitmap_44,bitmap_43,bitmap_42,bitmap_41,bitmap_40,_T_38}; // @[ReplacementPolicy.scala 87:33]
  assign _T_53 = {bitmap_55,bitmap_54,bitmap_53,bitmap_52,bitmap_51,bitmap_50,bitmap_49,bitmap_48}; // @[ReplacementPolicy.scala 87:33]
  assign _T_62 = {bitmap_63,bitmap_62,bitmap_61,bitmap_60,bitmap_59,bitmap_58,bitmap_57,bitmap_56,_T_53,_T_46}; // @[ReplacementPolicy.scala 87:33]
  assign bitmapU = {_T_62,_T_31}; // @[ReplacementPolicy.scala 87:33]
  assign _T_66 = bitmapU[62:0] == 63'h3fffffffffffffff; // @[ReplacementPolicy.scala 88:31]
  assign bitmapUNeg = ~bitmapU; // @[ReplacementPolicy.scala 92:47]
  assign _T_132 = bitmapUNeg[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  assign _T_133 = bitmapUNeg[61] ? 6'h3d : _T_132; // @[Mux.scala 47:69]
  assign _T_134 = bitmapUNeg[60] ? 6'h3c : _T_133; // @[Mux.scala 47:69]
  assign _T_135 = bitmapUNeg[59] ? 6'h3b : _T_134; // @[Mux.scala 47:69]
  assign _T_136 = bitmapUNeg[58] ? 6'h3a : _T_135; // @[Mux.scala 47:69]
  assign _T_137 = bitmapUNeg[57] ? 6'h39 : _T_136; // @[Mux.scala 47:69]
  assign _T_138 = bitmapUNeg[56] ? 6'h38 : _T_137; // @[Mux.scala 47:69]
  assign _T_139 = bitmapUNeg[55] ? 6'h37 : _T_138; // @[Mux.scala 47:69]
  assign _T_140 = bitmapUNeg[54] ? 6'h36 : _T_139; // @[Mux.scala 47:69]
  assign _T_141 = bitmapUNeg[53] ? 6'h35 : _T_140; // @[Mux.scala 47:69]
  assign _T_142 = bitmapUNeg[52] ? 6'h34 : _T_141; // @[Mux.scala 47:69]
  assign _T_143 = bitmapUNeg[51] ? 6'h33 : _T_142; // @[Mux.scala 47:69]
  assign _T_144 = bitmapUNeg[50] ? 6'h32 : _T_143; // @[Mux.scala 47:69]
  assign _T_145 = bitmapUNeg[49] ? 6'h31 : _T_144; // @[Mux.scala 47:69]
  assign _T_146 = bitmapUNeg[48] ? 6'h30 : _T_145; // @[Mux.scala 47:69]
  assign _T_147 = bitmapUNeg[47] ? 6'h2f : _T_146; // @[Mux.scala 47:69]
  assign _T_148 = bitmapUNeg[46] ? 6'h2e : _T_147; // @[Mux.scala 47:69]
  assign _T_149 = bitmapUNeg[45] ? 6'h2d : _T_148; // @[Mux.scala 47:69]
  assign _T_150 = bitmapUNeg[44] ? 6'h2c : _T_149; // @[Mux.scala 47:69]
  assign _T_151 = bitmapUNeg[43] ? 6'h2b : _T_150; // @[Mux.scala 47:69]
  assign _T_152 = bitmapUNeg[42] ? 6'h2a : _T_151; // @[Mux.scala 47:69]
  assign _T_153 = bitmapUNeg[41] ? 6'h29 : _T_152; // @[Mux.scala 47:69]
  assign _T_154 = bitmapUNeg[40] ? 6'h28 : _T_153; // @[Mux.scala 47:69]
  assign _T_155 = bitmapUNeg[39] ? 6'h27 : _T_154; // @[Mux.scala 47:69]
  assign _T_156 = bitmapUNeg[38] ? 6'h26 : _T_155; // @[Mux.scala 47:69]
  assign _T_157 = bitmapUNeg[37] ? 6'h25 : _T_156; // @[Mux.scala 47:69]
  assign _T_158 = bitmapUNeg[36] ? 6'h24 : _T_157; // @[Mux.scala 47:69]
  assign _T_159 = bitmapUNeg[35] ? 6'h23 : _T_158; // @[Mux.scala 47:69]
  assign _T_160 = bitmapUNeg[34] ? 6'h22 : _T_159; // @[Mux.scala 47:69]
  assign _T_161 = bitmapUNeg[33] ? 6'h21 : _T_160; // @[Mux.scala 47:69]
  assign _T_162 = bitmapUNeg[32] ? 6'h20 : _T_161; // @[Mux.scala 47:69]
  assign _T_163 = bitmapUNeg[31] ? 6'h1f : _T_162; // @[Mux.scala 47:69]
  assign _T_164 = bitmapUNeg[30] ? 6'h1e : _T_163; // @[Mux.scala 47:69]
  assign _T_165 = bitmapUNeg[29] ? 6'h1d : _T_164; // @[Mux.scala 47:69]
  assign _T_166 = bitmapUNeg[28] ? 6'h1c : _T_165; // @[Mux.scala 47:69]
  assign _T_167 = bitmapUNeg[27] ? 6'h1b : _T_166; // @[Mux.scala 47:69]
  assign _T_168 = bitmapUNeg[26] ? 6'h1a : _T_167; // @[Mux.scala 47:69]
  assign _T_169 = bitmapUNeg[25] ? 6'h19 : _T_168; // @[Mux.scala 47:69]
  assign _T_170 = bitmapUNeg[24] ? 6'h18 : _T_169; // @[Mux.scala 47:69]
  assign _T_171 = bitmapUNeg[23] ? 6'h17 : _T_170; // @[Mux.scala 47:69]
  assign _T_172 = bitmapUNeg[22] ? 6'h16 : _T_171; // @[Mux.scala 47:69]
  assign _T_173 = bitmapUNeg[21] ? 6'h15 : _T_172; // @[Mux.scala 47:69]
  assign _T_174 = bitmapUNeg[20] ? 6'h14 : _T_173; // @[Mux.scala 47:69]
  assign _T_175 = bitmapUNeg[19] ? 6'h13 : _T_174; // @[Mux.scala 47:69]
  assign _T_176 = bitmapUNeg[18] ? 6'h12 : _T_175; // @[Mux.scala 47:69]
  assign _T_177 = bitmapUNeg[17] ? 6'h11 : _T_176; // @[Mux.scala 47:69]
  assign _T_178 = bitmapUNeg[16] ? 6'h10 : _T_177; // @[Mux.scala 47:69]
  assign _T_179 = bitmapUNeg[15] ? 6'hf : _T_178; // @[Mux.scala 47:69]
  assign _T_180 = bitmapUNeg[14] ? 6'he : _T_179; // @[Mux.scala 47:69]
  assign _T_181 = bitmapUNeg[13] ? 6'hd : _T_180; // @[Mux.scala 47:69]
  assign _T_182 = bitmapUNeg[12] ? 6'hc : _T_181; // @[Mux.scala 47:69]
  assign _T_183 = bitmapUNeg[11] ? 6'hb : _T_182; // @[Mux.scala 47:69]
  assign _T_184 = bitmapUNeg[10] ? 6'ha : _T_183; // @[Mux.scala 47:69]
  assign _T_185 = bitmapUNeg[9] ? 6'h9 : _T_184; // @[Mux.scala 47:69]
  assign _T_186 = bitmapUNeg[8] ? 6'h8 : _T_185; // @[Mux.scala 47:69]
  assign _T_187 = bitmapUNeg[7] ? 6'h7 : _T_186; // @[Mux.scala 47:69]
  assign _T_188 = bitmapUNeg[6] ? 6'h6 : _T_187; // @[Mux.scala 47:69]
  assign _T_189 = bitmapUNeg[5] ? 6'h5 : _T_188; // @[Mux.scala 47:69]
  assign _T_190 = bitmapUNeg[4] ? 6'h4 : _T_189; // @[Mux.scala 47:69]
  assign _T_191 = bitmapUNeg[3] ? 6'h3 : _T_190; // @[Mux.scala 47:69]
  assign _T_192 = bitmapUNeg[2] ? 6'h2 : _T_191; // @[Mux.scala 47:69]
  assign _T_193 = bitmapUNeg[1] ? 6'h1 : _T_192; // @[Mux.scala 47:69]
  assign io_lru_idx = bitmapUNeg[0] ? 6'h0 : _T_193; // @[ReplacementPolicy.scala 93:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  bitmap_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  bitmap_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  bitmap_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  bitmap_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  bitmap_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  bitmap_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  bitmap_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  bitmap_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  bitmap_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  bitmap_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  bitmap_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  bitmap_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  bitmap_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  bitmap_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  bitmap_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  bitmap_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  bitmap_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  bitmap_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  bitmap_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  bitmap_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  bitmap_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  bitmap_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  bitmap_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  bitmap_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  bitmap_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  bitmap_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  bitmap_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  bitmap_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  bitmap_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  bitmap_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  bitmap_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  bitmap_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  bitmap_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  bitmap_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  bitmap_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  bitmap_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  bitmap_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  bitmap_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  bitmap_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  bitmap_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  bitmap_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  bitmap_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  bitmap_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  bitmap_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  bitmap_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  bitmap_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  bitmap_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  bitmap_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  bitmap_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  bitmap_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  bitmap_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  bitmap_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  bitmap_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  bitmap_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  bitmap_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  bitmap_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  bitmap_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  bitmap_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  bitmap_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  bitmap_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  bitmap_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  bitmap_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  bitmap_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      bitmap_0 <= 1'h0;
    end else if (_T_66) begin
      bitmap_0 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_0 <= _GEN_128;
    end else if (io_idx_1_valid) begin
      bitmap_0 <= _GEN_0;
    end
    if (reset) begin
      bitmap_1 <= 1'h0;
    end else if (_T_66) begin
      bitmap_1 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_1 <= _GEN_129;
    end else if (io_idx_1_valid) begin
      bitmap_1 <= _GEN_1;
    end
    if (reset) begin
      bitmap_2 <= 1'h0;
    end else if (_T_66) begin
      bitmap_2 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_2 <= _GEN_130;
    end else if (io_idx_1_valid) begin
      bitmap_2 <= _GEN_2;
    end
    if (reset) begin
      bitmap_3 <= 1'h0;
    end else if (_T_66) begin
      bitmap_3 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_3 <= _GEN_131;
    end else if (io_idx_1_valid) begin
      bitmap_3 <= _GEN_3;
    end
    if (reset) begin
      bitmap_4 <= 1'h0;
    end else if (_T_66) begin
      bitmap_4 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_4 <= _GEN_132;
    end else if (io_idx_1_valid) begin
      bitmap_4 <= _GEN_4;
    end
    if (reset) begin
      bitmap_5 <= 1'h0;
    end else if (_T_66) begin
      bitmap_5 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_5 <= _GEN_133;
    end else if (io_idx_1_valid) begin
      bitmap_5 <= _GEN_5;
    end
    if (reset) begin
      bitmap_6 <= 1'h0;
    end else if (_T_66) begin
      bitmap_6 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_6 <= _GEN_134;
    end else if (io_idx_1_valid) begin
      bitmap_6 <= _GEN_6;
    end
    if (reset) begin
      bitmap_7 <= 1'h0;
    end else if (_T_66) begin
      bitmap_7 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_7 <= _GEN_135;
    end else if (io_idx_1_valid) begin
      bitmap_7 <= _GEN_7;
    end
    if (reset) begin
      bitmap_8 <= 1'h0;
    end else if (_T_66) begin
      bitmap_8 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_8 <= _GEN_136;
    end else if (io_idx_1_valid) begin
      bitmap_8 <= _GEN_8;
    end
    if (reset) begin
      bitmap_9 <= 1'h0;
    end else if (_T_66) begin
      bitmap_9 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_9 <= _GEN_137;
    end else if (io_idx_1_valid) begin
      bitmap_9 <= _GEN_9;
    end
    if (reset) begin
      bitmap_10 <= 1'h0;
    end else if (_T_66) begin
      bitmap_10 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_10 <= _GEN_138;
    end else if (io_idx_1_valid) begin
      bitmap_10 <= _GEN_10;
    end
    if (reset) begin
      bitmap_11 <= 1'h0;
    end else if (_T_66) begin
      bitmap_11 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_11 <= _GEN_139;
    end else if (io_idx_1_valid) begin
      bitmap_11 <= _GEN_11;
    end
    if (reset) begin
      bitmap_12 <= 1'h0;
    end else if (_T_66) begin
      bitmap_12 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_12 <= _GEN_140;
    end else if (io_idx_1_valid) begin
      bitmap_12 <= _GEN_12;
    end
    if (reset) begin
      bitmap_13 <= 1'h0;
    end else if (_T_66) begin
      bitmap_13 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_13 <= _GEN_141;
    end else if (io_idx_1_valid) begin
      bitmap_13 <= _GEN_13;
    end
    if (reset) begin
      bitmap_14 <= 1'h0;
    end else if (_T_66) begin
      bitmap_14 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_14 <= _GEN_142;
    end else if (io_idx_1_valid) begin
      bitmap_14 <= _GEN_14;
    end
    if (reset) begin
      bitmap_15 <= 1'h0;
    end else if (_T_66) begin
      bitmap_15 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_15 <= _GEN_143;
    end else if (io_idx_1_valid) begin
      bitmap_15 <= _GEN_15;
    end
    if (reset) begin
      bitmap_16 <= 1'h0;
    end else if (_T_66) begin
      bitmap_16 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_16 <= _GEN_144;
    end else if (io_idx_1_valid) begin
      bitmap_16 <= _GEN_16;
    end
    if (reset) begin
      bitmap_17 <= 1'h0;
    end else if (_T_66) begin
      bitmap_17 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_17 <= _GEN_145;
    end else if (io_idx_1_valid) begin
      bitmap_17 <= _GEN_17;
    end
    if (reset) begin
      bitmap_18 <= 1'h0;
    end else if (_T_66) begin
      bitmap_18 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_18 <= _GEN_146;
    end else if (io_idx_1_valid) begin
      bitmap_18 <= _GEN_18;
    end
    if (reset) begin
      bitmap_19 <= 1'h0;
    end else if (_T_66) begin
      bitmap_19 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_19 <= _GEN_147;
    end else if (io_idx_1_valid) begin
      bitmap_19 <= _GEN_19;
    end
    if (reset) begin
      bitmap_20 <= 1'h0;
    end else if (_T_66) begin
      bitmap_20 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_20 <= _GEN_148;
    end else if (io_idx_1_valid) begin
      bitmap_20 <= _GEN_20;
    end
    if (reset) begin
      bitmap_21 <= 1'h0;
    end else if (_T_66) begin
      bitmap_21 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_21 <= _GEN_149;
    end else if (io_idx_1_valid) begin
      bitmap_21 <= _GEN_21;
    end
    if (reset) begin
      bitmap_22 <= 1'h0;
    end else if (_T_66) begin
      bitmap_22 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_22 <= _GEN_150;
    end else if (io_idx_1_valid) begin
      bitmap_22 <= _GEN_22;
    end
    if (reset) begin
      bitmap_23 <= 1'h0;
    end else if (_T_66) begin
      bitmap_23 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_23 <= _GEN_151;
    end else if (io_idx_1_valid) begin
      bitmap_23 <= _GEN_23;
    end
    if (reset) begin
      bitmap_24 <= 1'h0;
    end else if (_T_66) begin
      bitmap_24 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_24 <= _GEN_152;
    end else if (io_idx_1_valid) begin
      bitmap_24 <= _GEN_24;
    end
    if (reset) begin
      bitmap_25 <= 1'h0;
    end else if (_T_66) begin
      bitmap_25 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_25 <= _GEN_153;
    end else if (io_idx_1_valid) begin
      bitmap_25 <= _GEN_25;
    end
    if (reset) begin
      bitmap_26 <= 1'h0;
    end else if (_T_66) begin
      bitmap_26 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_26 <= _GEN_154;
    end else if (io_idx_1_valid) begin
      bitmap_26 <= _GEN_26;
    end
    if (reset) begin
      bitmap_27 <= 1'h0;
    end else if (_T_66) begin
      bitmap_27 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_27 <= _GEN_155;
    end else if (io_idx_1_valid) begin
      bitmap_27 <= _GEN_27;
    end
    if (reset) begin
      bitmap_28 <= 1'h0;
    end else if (_T_66) begin
      bitmap_28 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_28 <= _GEN_156;
    end else if (io_idx_1_valid) begin
      bitmap_28 <= _GEN_28;
    end
    if (reset) begin
      bitmap_29 <= 1'h0;
    end else if (_T_66) begin
      bitmap_29 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_29 <= _GEN_157;
    end else if (io_idx_1_valid) begin
      bitmap_29 <= _GEN_29;
    end
    if (reset) begin
      bitmap_30 <= 1'h0;
    end else if (_T_66) begin
      bitmap_30 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_30 <= _GEN_158;
    end else if (io_idx_1_valid) begin
      bitmap_30 <= _GEN_30;
    end
    if (reset) begin
      bitmap_31 <= 1'h0;
    end else if (_T_66) begin
      bitmap_31 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_31 <= _GEN_159;
    end else if (io_idx_1_valid) begin
      bitmap_31 <= _GEN_31;
    end
    if (reset) begin
      bitmap_32 <= 1'h0;
    end else if (_T_66) begin
      bitmap_32 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_32 <= _GEN_160;
    end else if (io_idx_1_valid) begin
      bitmap_32 <= _GEN_32;
    end
    if (reset) begin
      bitmap_33 <= 1'h0;
    end else if (_T_66) begin
      bitmap_33 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_33 <= _GEN_161;
    end else if (io_idx_1_valid) begin
      bitmap_33 <= _GEN_33;
    end
    if (reset) begin
      bitmap_34 <= 1'h0;
    end else if (_T_66) begin
      bitmap_34 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_34 <= _GEN_162;
    end else if (io_idx_1_valid) begin
      bitmap_34 <= _GEN_34;
    end
    if (reset) begin
      bitmap_35 <= 1'h0;
    end else if (_T_66) begin
      bitmap_35 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_35 <= _GEN_163;
    end else if (io_idx_1_valid) begin
      bitmap_35 <= _GEN_35;
    end
    if (reset) begin
      bitmap_36 <= 1'h0;
    end else if (_T_66) begin
      bitmap_36 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_36 <= _GEN_164;
    end else if (io_idx_1_valid) begin
      bitmap_36 <= _GEN_36;
    end
    if (reset) begin
      bitmap_37 <= 1'h0;
    end else if (_T_66) begin
      bitmap_37 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_37 <= _GEN_165;
    end else if (io_idx_1_valid) begin
      bitmap_37 <= _GEN_37;
    end
    if (reset) begin
      bitmap_38 <= 1'h0;
    end else if (_T_66) begin
      bitmap_38 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_38 <= _GEN_166;
    end else if (io_idx_1_valid) begin
      bitmap_38 <= _GEN_38;
    end
    if (reset) begin
      bitmap_39 <= 1'h0;
    end else if (_T_66) begin
      bitmap_39 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_39 <= _GEN_167;
    end else if (io_idx_1_valid) begin
      bitmap_39 <= _GEN_39;
    end
    if (reset) begin
      bitmap_40 <= 1'h0;
    end else if (_T_66) begin
      bitmap_40 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_40 <= _GEN_168;
    end else if (io_idx_1_valid) begin
      bitmap_40 <= _GEN_40;
    end
    if (reset) begin
      bitmap_41 <= 1'h0;
    end else if (_T_66) begin
      bitmap_41 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_41 <= _GEN_169;
    end else if (io_idx_1_valid) begin
      bitmap_41 <= _GEN_41;
    end
    if (reset) begin
      bitmap_42 <= 1'h0;
    end else if (_T_66) begin
      bitmap_42 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_42 <= _GEN_170;
    end else if (io_idx_1_valid) begin
      bitmap_42 <= _GEN_42;
    end
    if (reset) begin
      bitmap_43 <= 1'h0;
    end else if (_T_66) begin
      bitmap_43 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_43 <= _GEN_171;
    end else if (io_idx_1_valid) begin
      bitmap_43 <= _GEN_43;
    end
    if (reset) begin
      bitmap_44 <= 1'h0;
    end else if (_T_66) begin
      bitmap_44 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_44 <= _GEN_172;
    end else if (io_idx_1_valid) begin
      bitmap_44 <= _GEN_44;
    end
    if (reset) begin
      bitmap_45 <= 1'h0;
    end else if (_T_66) begin
      bitmap_45 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_45 <= _GEN_173;
    end else if (io_idx_1_valid) begin
      bitmap_45 <= _GEN_45;
    end
    if (reset) begin
      bitmap_46 <= 1'h0;
    end else if (_T_66) begin
      bitmap_46 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_46 <= _GEN_174;
    end else if (io_idx_1_valid) begin
      bitmap_46 <= _GEN_46;
    end
    if (reset) begin
      bitmap_47 <= 1'h0;
    end else if (_T_66) begin
      bitmap_47 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_47 <= _GEN_175;
    end else if (io_idx_1_valid) begin
      bitmap_47 <= _GEN_47;
    end
    if (reset) begin
      bitmap_48 <= 1'h0;
    end else if (_T_66) begin
      bitmap_48 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_48 <= _GEN_176;
    end else if (io_idx_1_valid) begin
      bitmap_48 <= _GEN_48;
    end
    if (reset) begin
      bitmap_49 <= 1'h0;
    end else if (_T_66) begin
      bitmap_49 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_49 <= _GEN_177;
    end else if (io_idx_1_valid) begin
      bitmap_49 <= _GEN_49;
    end
    if (reset) begin
      bitmap_50 <= 1'h0;
    end else if (_T_66) begin
      bitmap_50 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_50 <= _GEN_178;
    end else if (io_idx_1_valid) begin
      bitmap_50 <= _GEN_50;
    end
    if (reset) begin
      bitmap_51 <= 1'h0;
    end else if (_T_66) begin
      bitmap_51 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_51 <= _GEN_179;
    end else if (io_idx_1_valid) begin
      bitmap_51 <= _GEN_51;
    end
    if (reset) begin
      bitmap_52 <= 1'h0;
    end else if (_T_66) begin
      bitmap_52 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_52 <= _GEN_180;
    end else if (io_idx_1_valid) begin
      bitmap_52 <= _GEN_52;
    end
    if (reset) begin
      bitmap_53 <= 1'h0;
    end else if (_T_66) begin
      bitmap_53 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_53 <= _GEN_181;
    end else if (io_idx_1_valid) begin
      bitmap_53 <= _GEN_53;
    end
    if (reset) begin
      bitmap_54 <= 1'h0;
    end else if (_T_66) begin
      bitmap_54 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_54 <= _GEN_182;
    end else if (io_idx_1_valid) begin
      bitmap_54 <= _GEN_54;
    end
    if (reset) begin
      bitmap_55 <= 1'h0;
    end else if (_T_66) begin
      bitmap_55 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_55 <= _GEN_183;
    end else if (io_idx_1_valid) begin
      bitmap_55 <= _GEN_55;
    end
    if (reset) begin
      bitmap_56 <= 1'h0;
    end else if (_T_66) begin
      bitmap_56 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_56 <= _GEN_184;
    end else if (io_idx_1_valid) begin
      bitmap_56 <= _GEN_56;
    end
    if (reset) begin
      bitmap_57 <= 1'h0;
    end else if (_T_66) begin
      bitmap_57 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_57 <= _GEN_185;
    end else if (io_idx_1_valid) begin
      bitmap_57 <= _GEN_57;
    end
    if (reset) begin
      bitmap_58 <= 1'h0;
    end else if (_T_66) begin
      bitmap_58 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_58 <= _GEN_186;
    end else if (io_idx_1_valid) begin
      bitmap_58 <= _GEN_58;
    end
    if (reset) begin
      bitmap_59 <= 1'h0;
    end else if (_T_66) begin
      bitmap_59 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_59 <= _GEN_187;
    end else if (io_idx_1_valid) begin
      bitmap_59 <= _GEN_59;
    end
    if (reset) begin
      bitmap_60 <= 1'h0;
    end else if (_T_66) begin
      bitmap_60 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_60 <= _GEN_188;
    end else if (io_idx_1_valid) begin
      bitmap_60 <= _GEN_60;
    end
    if (reset) begin
      bitmap_61 <= 1'h0;
    end else if (_T_66) begin
      bitmap_61 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_61 <= _GEN_189;
    end else if (io_idx_1_valid) begin
      bitmap_61 <= _GEN_61;
    end
    if (reset) begin
      bitmap_62 <= 1'h0;
    end else if (_T_66) begin
      bitmap_62 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_62 <= _GEN_190;
    end else if (io_idx_1_valid) begin
      bitmap_62 <= _GEN_62;
    end
    if (reset) begin
      bitmap_63 <= 1'h0;
    end else if (_T_66) begin
      bitmap_63 <= 1'h0;
    end else if (io_idx_2_valid) begin
      bitmap_63 <= _GEN_191;
    end else if (io_idx_1_valid) begin
      bitmap_63 <= _GEN_63;
    end
  end
endmodule
