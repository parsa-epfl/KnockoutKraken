module BranchUnit( // @[:@2856.2]
  input  [25:0] io_dinst_imm_bits, // @[:@2859.4]
  input  [3:0]  io_dinst_cond_bits, // @[:@2859.4]
  input  [2:0]  io_dinst_itype, // @[:@2859.4]
  input  [2:0]  io_dinst_op, // @[:@2859.4]
  input  [3:0]  io_nzcv, // @[:@2859.4]
  output        io_binst_valid, // @[:@2859.4]
  output [63:0] io_binst_bits_offset // @[:@2859.4]
);
  wire [3:0] cond_io_cond; // @[branch.scala 59:20:@2867.4]
  wire [3:0] cond_io_nzcv; // @[branch.scala 59:20:@2867.4]
  wire  cond_io_res; // @[branch.scala 59:20:@2867.4]
  wire [25:0] _T_99; // @[branch.scala 55:37:@2863.4]
  wire [63:0] signExtended; // @[branch.scala 54:26:@2862.4 branch.scala 55:16:@2864.4]
  wire  _T_101; // @[branch.scala 62:24:@2872.4]
  wire  _T_102; // @[branch.scala 62:54:@2873.4]
  wire  _T_103; // @[branch.scala 62:36:@2874.4]
  wire  _T_104; // @[branch.scala 63:22:@2876.6]
  wire  _T_105; // @[branch.scala 65:28:@2881.8]
  wire  _GEN_1; // @[branch.scala 63:36:@2877.6]
  CondUnit cond ( // @[branch.scala 59:20:@2867.4]
    .io_cond(cond_io_cond),
    .io_nzcv(cond_io_nzcv),
    .io_res(cond_io_res)
  );
  assign _T_99 = $signed(io_dinst_imm_bits); // @[branch.scala 55:37:@2863.4]
  assign signExtended = {{38{_T_99[25]}},_T_99}; // @[branch.scala 54:26:@2862.4 branch.scala 55:16:@2864.4]
  assign _T_101 = io_dinst_itype == 3'h2; // @[branch.scala 62:24:@2872.4]
  assign _T_102 = io_dinst_itype == 3'h3; // @[branch.scala 62:54:@2873.4]
  assign _T_103 = _T_101 | _T_102; // @[branch.scala 62:36:@2874.4]
  assign _T_104 = io_dinst_op == 3'h1; // @[branch.scala 63:22:@2876.6]
  assign _T_105 = io_dinst_op == 3'h0; // @[branch.scala 65:28:@2881.8]
  assign _GEN_1 = _T_104 ? cond_io_res : _T_105; // @[branch.scala 63:36:@2877.6]
  assign io_binst_valid = _T_103 ? _GEN_1 : 1'h0; // @[branch.scala 51:18:@2861.4 branch.scala 64:22:@2878.8 branch.scala 66:22:@2883.10]
  assign io_binst_bits_offset = $unsigned(signExtended); // @[branch.scala 56:24:@2866.4]
  assign cond_io_cond = io_dinst_cond_bits; // @[branch.scala 60:16:@2870.4]
  assign cond_io_nzcv = io_nzcv; // @[branch.scala 61:16:@2871.4]
endmodule
