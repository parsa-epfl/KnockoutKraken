module CondUnit( // @[:@2594.2]
  input  [3:0] io_cond, // @[:@2597.4]
  input  [3:0] io_nzcv, // @[:@2597.4]
  output       io_res // @[:@2597.4]
);
  wire [2:0] _T_13; // @[branch.scala 23:21:@2601.4]
  wire  _T_15; // @[branch.scala 23:27:@2602.4]
  wire  _T_16; // @[branch.scala 23:60:@2604.6]
  wire  _T_21; // @[branch.scala 24:27:@2610.6]
  wire  _T_22; // @[branch.scala 24:60:@2612.8]
  wire  _T_27; // @[branch.scala 25:27:@2618.8]
  wire  _T_28; // @[branch.scala 25:60:@2620.10]
  wire  _T_33; // @[branch.scala 26:27:@2626.10]
  wire  _T_34; // @[branch.scala 26:60:@2628.12]
  wire  _T_39; // @[branch.scala 27:27:@2634.12]
  wire  _T_45; // @[branch.scala 28:27:@2642.14]
  wire  _T_51; // @[branch.scala 29:27:@2650.16]
  wire  _T_57; // @[branch.scala 30:27:@2658.18]
  wire  _GEN_1; // @[branch.scala 29:41:@2651.16]
  wire  _GEN_2; // @[branch.scala 28:41:@2643.14]
  wire  _GEN_3; // @[branch.scala 27:41:@2635.12]
  wire  _GEN_4; // @[branch.scala 26:41:@2627.10]
  wire  _GEN_5; // @[branch.scala 25:41:@2619.8]
  wire  _GEN_6; // @[branch.scala 24:41:@2611.6]
  wire  result; // @[branch.scala 23:41:@2603.4]
  wire  _T_59; // @[branch.scala 32:15:@2662.4]
  wire  _T_63; // @[branch.scala 32:38:@2664.4]
  wire  _T_64; // @[branch.scala 32:27:@2665.4]
  wire  _T_66; // @[branch.scala 33:15:@2667.6]
  assign _T_13 = io_cond[3:1]; // @[branch.scala 23:21:@2601.4]
  assign _T_15 = _T_13 == 3'h0; // @[branch.scala 23:27:@2602.4]
  assign _T_16 = io_nzcv[2]; // @[branch.scala 23:60:@2604.6]
  assign _T_21 = _T_13 == 3'h1; // @[branch.scala 24:27:@2610.6]
  assign _T_22 = io_nzcv[1]; // @[branch.scala 24:60:@2612.8]
  assign _T_27 = _T_13 == 3'h2; // @[branch.scala 25:27:@2618.8]
  assign _T_28 = io_nzcv[3]; // @[branch.scala 25:60:@2620.10]
  assign _T_33 = _T_13 == 3'h3; // @[branch.scala 26:27:@2626.10]
  assign _T_34 = io_nzcv[0]; // @[branch.scala 26:60:@2628.12]
  assign _T_39 = _T_13 == 3'h4; // @[branch.scala 27:27:@2634.12]
  assign _T_45 = _T_13 == 3'h5; // @[branch.scala 28:27:@2642.14]
  assign _T_51 = _T_13 == 3'h6; // @[branch.scala 29:27:@2650.16]
  assign _T_57 = _T_13 == 3'h7; // @[branch.scala 30:27:@2658.18]
  assign _GEN_1 = _T_51 ? _T_28 : _T_57; // @[branch.scala 29:41:@2651.16]
  assign _GEN_2 = _T_45 ? _T_28 : _GEN_1; // @[branch.scala 28:41:@2643.14]
  assign _GEN_3 = _T_39 ? _T_22 : _GEN_2; // @[branch.scala 27:41:@2635.12]
  assign _GEN_4 = _T_33 ? _T_34 : _GEN_3; // @[branch.scala 26:41:@2627.10]
  assign _GEN_5 = _T_27 ? _T_28 : _GEN_4; // @[branch.scala 25:41:@2619.8]
  assign _GEN_6 = _T_21 ? _T_22 : _GEN_5; // @[branch.scala 24:41:@2611.6]
  assign result = _T_15 ? _T_16 : _GEN_6; // @[branch.scala 23:41:@2603.4]
  assign _T_59 = io_cond[0]; // @[branch.scala 32:15:@2662.4]
  assign _T_63 = io_cond != 4'hf; // @[branch.scala 32:38:@2664.4]
  assign _T_64 = _T_59 & _T_63; // @[branch.scala 32:27:@2665.4]
  assign _T_66 = result == 1'h0; // @[branch.scala 33:15:@2667.6]
  assign io_res = _T_64 ? _T_66 : result; // @[branch.scala 33:12:@2668.6 branch.scala 35:12:@2671.6]
endmodule
