module TLBUnit( // @[:@452.2]
  input         clock, // @[:@453.4]
  input         reset, // @[:@454.4]
  input  [63:0] io_vaddrFill, // @[:@455.4]
  input         io_fill, // @[:@455.4]
  input         io_vaddr_valid, // @[:@455.4]
  input  [63:0] io_vaddr_bits, // @[:@455.4]
  output        io_hit, // @[:@455.4]
  output        io_paddr_valid, // @[:@455.4]
  output [63:0] io_paddr_bits // @[:@455.4]
);
  wire [53:0] vpage; // @[TLB.scala 20:29:@457.4]
  wire [4:0] vpageTLB; // @[TLB.scala 21:23:@458.4]
  wire [48:0] vpageTAG; // @[TLB.scala 22:24:@459.4]
  wire [53:0] vpageFill; // @[TLB.scala 24:32:@460.4]
  wire [4:0] vpageFillTLB; // @[TLB.scala 25:31:@461.4]
  wire [48:0] vpageFillTAG; // @[TLB.scala 26:32:@462.4]
  reg  tlb_0_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_0;
  reg [48:0] tlb_0_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_1;
  reg  tlb_1_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_2;
  reg [48:0] tlb_1_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_3;
  reg  tlb_2_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_4;
  reg [48:0] tlb_2_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_5;
  reg  tlb_3_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_6;
  reg [48:0] tlb_3_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_7;
  reg  tlb_4_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_8;
  reg [48:0] tlb_4_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_9;
  reg  tlb_5_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_10;
  reg [48:0] tlb_5_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_11;
  reg  tlb_6_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_12;
  reg [48:0] tlb_6_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_13;
  reg  tlb_7_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_14;
  reg [48:0] tlb_7_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_15;
  reg  tlb_8_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_16;
  reg [48:0] tlb_8_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_17;
  reg  tlb_9_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_18;
  reg [48:0] tlb_9_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_19;
  reg  tlb_10_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_20;
  reg [48:0] tlb_10_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_21;
  reg  tlb_11_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_22;
  reg [48:0] tlb_11_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_23;
  reg  tlb_12_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_24;
  reg [48:0] tlb_12_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_25;
  reg  tlb_13_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_26;
  reg [48:0] tlb_13_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_27;
  reg  tlb_14_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_28;
  reg [48:0] tlb_14_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_29;
  reg  tlb_15_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_30;
  reg [48:0] tlb_15_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_31;
  reg  tlb_16_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_32;
  reg [48:0] tlb_16_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_33;
  reg  tlb_17_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_34;
  reg [48:0] tlb_17_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_35;
  reg  tlb_18_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_36;
  reg [48:0] tlb_18_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_37;
  reg  tlb_19_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_38;
  reg [48:0] tlb_19_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_39;
  reg  tlb_20_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_40;
  reg [48:0] tlb_20_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_41;
  reg  tlb_21_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_42;
  reg [48:0] tlb_21_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_43;
  reg  tlb_22_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_44;
  reg [48:0] tlb_22_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_45;
  reg  tlb_23_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_46;
  reg [48:0] tlb_23_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_47;
  reg  tlb_24_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_48;
  reg [48:0] tlb_24_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_49;
  reg  tlb_25_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_50;
  reg [48:0] tlb_25_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_51;
  reg  tlb_26_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_52;
  reg [48:0] tlb_26_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_53;
  reg  tlb_27_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_54;
  reg [48:0] tlb_27_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_55;
  reg  tlb_28_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_56;
  reg [48:0] tlb_28_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_57;
  reg  tlb_29_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_58;
  reg [48:0] tlb_29_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_59;
  reg  tlb_30_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_60;
  reg [48:0] tlb_30_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_61;
  reg  tlb_31_valid; // @[TLB.scala 35:20:@531.4]
  reg [31:0] _RAND_62;
  reg [48:0] tlb_31_bits; // @[TLB.scala 35:20:@531.4]
  reg [63:0] _RAND_63;
  wire [48:0] _GEN_0; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_1; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_2; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_3; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_4; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_5; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_6; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_7; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_8; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_9; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_10; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_11; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_12; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_13; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_14; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_15; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_16; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_17; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_18; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_19; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_20; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_21; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_22; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_23; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_24; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_25; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_26; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_27; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_28; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_29; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_30; // @[TLB.scala 37:28:@533.6]
  wire [48:0] _GEN_31; // @[TLB.scala 37:28:@533.6]
  wire  _GEN_32; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_33; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_34; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_35; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_36; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_37; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_38; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_39; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_40; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_41; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_42; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_43; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_44; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_45; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_46; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_47; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_48; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_49; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_50; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_51; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_52; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_53; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_54; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_55; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_56; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_57; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_58; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_59; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_60; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_61; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_62; // @[TLB.scala 38:29:@534.6]
  wire  _GEN_63; // @[TLB.scala 38:29:@534.6]
  wire [48:0] _GEN_64; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_65; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_66; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_67; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_68; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_69; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_70; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_71; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_72; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_73; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_74; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_75; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_76; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_77; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_78; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_79; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_80; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_81; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_82; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_83; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_84; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_85; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_86; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_87; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_88; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_89; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_90; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_91; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_92; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_93; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_94; // @[TLB.scala 36:17:@532.4]
  wire [48:0] _GEN_95; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_96; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_97; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_98; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_99; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_100; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_101; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_102; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_103; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_104; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_105; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_106; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_107; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_108; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_109; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_110; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_111; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_112; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_113; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_114; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_115; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_116; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_117; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_118; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_119; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_120; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_121; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_122; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_123; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_124; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_125; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_126; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_127; // @[TLB.scala 36:17:@532.4]
  wire  _GEN_130; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_131; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_132; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_133; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_134; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_135; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_136; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_137; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_138; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_139; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_140; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_141; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_142; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_143; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_144; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_145; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_146; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_147; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_148; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_149; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_150; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_151; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_152; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_153; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_154; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_155; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_156; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_157; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_158; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_159; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_160; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_161; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_162; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_163; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_164; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_165; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_166; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_167; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_168; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_169; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_170; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_171; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_172; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_173; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_174; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_175; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_176; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_177; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_178; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_179; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_180; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_181; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_182; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_183; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_184; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_185; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_186; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_187; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_188; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_189; // @[TLB.scala 41:56:@536.4]
  wire  _GEN_190; // @[TLB.scala 41:56:@536.4]
  wire [48:0] _GEN_191; // @[TLB.scala 41:56:@536.4]
  wire  _T_616; // @[TLB.scala 42:55:@539.4]
  assign vpage = io_vaddr_bits[63:10]; // @[TLB.scala 20:29:@457.4]
  assign vpageTLB = vpage[4:0]; // @[TLB.scala 21:23:@458.4]
  assign vpageTAG = vpage[53:5]; // @[TLB.scala 22:24:@459.4]
  assign vpageFill = io_vaddrFill[63:10]; // @[TLB.scala 24:32:@460.4]
  assign vpageFillTLB = vpageFill[4:0]; // @[TLB.scala 25:31:@461.4]
  assign vpageFillTAG = vpageFill[53:5]; // @[TLB.scala 26:32:@462.4]
  assign _GEN_0 = 5'h0 == vpageFillTLB ? vpageFillTAG : tlb_0_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_1 = 5'h1 == vpageFillTLB ? vpageFillTAG : tlb_1_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_2 = 5'h2 == vpageFillTLB ? vpageFillTAG : tlb_2_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_3 = 5'h3 == vpageFillTLB ? vpageFillTAG : tlb_3_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_4 = 5'h4 == vpageFillTLB ? vpageFillTAG : tlb_4_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_5 = 5'h5 == vpageFillTLB ? vpageFillTAG : tlb_5_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_6 = 5'h6 == vpageFillTLB ? vpageFillTAG : tlb_6_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_7 = 5'h7 == vpageFillTLB ? vpageFillTAG : tlb_7_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_8 = 5'h8 == vpageFillTLB ? vpageFillTAG : tlb_8_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_9 = 5'h9 == vpageFillTLB ? vpageFillTAG : tlb_9_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_10 = 5'ha == vpageFillTLB ? vpageFillTAG : tlb_10_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_11 = 5'hb == vpageFillTLB ? vpageFillTAG : tlb_11_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_12 = 5'hc == vpageFillTLB ? vpageFillTAG : tlb_12_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_13 = 5'hd == vpageFillTLB ? vpageFillTAG : tlb_13_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_14 = 5'he == vpageFillTLB ? vpageFillTAG : tlb_14_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_15 = 5'hf == vpageFillTLB ? vpageFillTAG : tlb_15_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_16 = 5'h10 == vpageFillTLB ? vpageFillTAG : tlb_16_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_17 = 5'h11 == vpageFillTLB ? vpageFillTAG : tlb_17_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_18 = 5'h12 == vpageFillTLB ? vpageFillTAG : tlb_18_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_19 = 5'h13 == vpageFillTLB ? vpageFillTAG : tlb_19_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_20 = 5'h14 == vpageFillTLB ? vpageFillTAG : tlb_20_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_21 = 5'h15 == vpageFillTLB ? vpageFillTAG : tlb_21_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_22 = 5'h16 == vpageFillTLB ? vpageFillTAG : tlb_22_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_23 = 5'h17 == vpageFillTLB ? vpageFillTAG : tlb_23_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_24 = 5'h18 == vpageFillTLB ? vpageFillTAG : tlb_24_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_25 = 5'h19 == vpageFillTLB ? vpageFillTAG : tlb_25_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_26 = 5'h1a == vpageFillTLB ? vpageFillTAG : tlb_26_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_27 = 5'h1b == vpageFillTLB ? vpageFillTAG : tlb_27_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_28 = 5'h1c == vpageFillTLB ? vpageFillTAG : tlb_28_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_29 = 5'h1d == vpageFillTLB ? vpageFillTAG : tlb_29_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_30 = 5'h1e == vpageFillTLB ? vpageFillTAG : tlb_30_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_31 = 5'h1f == vpageFillTLB ? vpageFillTAG : tlb_31_bits; // @[TLB.scala 37:28:@533.6]
  assign _GEN_32 = 5'h0 == vpageFillTLB ? 1'h1 : tlb_0_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_33 = 5'h1 == vpageFillTLB ? 1'h1 : tlb_1_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_34 = 5'h2 == vpageFillTLB ? 1'h1 : tlb_2_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_35 = 5'h3 == vpageFillTLB ? 1'h1 : tlb_3_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_36 = 5'h4 == vpageFillTLB ? 1'h1 : tlb_4_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_37 = 5'h5 == vpageFillTLB ? 1'h1 : tlb_5_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_38 = 5'h6 == vpageFillTLB ? 1'h1 : tlb_6_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_39 = 5'h7 == vpageFillTLB ? 1'h1 : tlb_7_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_40 = 5'h8 == vpageFillTLB ? 1'h1 : tlb_8_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_41 = 5'h9 == vpageFillTLB ? 1'h1 : tlb_9_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_42 = 5'ha == vpageFillTLB ? 1'h1 : tlb_10_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_43 = 5'hb == vpageFillTLB ? 1'h1 : tlb_11_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_44 = 5'hc == vpageFillTLB ? 1'h1 : tlb_12_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_45 = 5'hd == vpageFillTLB ? 1'h1 : tlb_13_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_46 = 5'he == vpageFillTLB ? 1'h1 : tlb_14_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_47 = 5'hf == vpageFillTLB ? 1'h1 : tlb_15_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_48 = 5'h10 == vpageFillTLB ? 1'h1 : tlb_16_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_49 = 5'h11 == vpageFillTLB ? 1'h1 : tlb_17_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_50 = 5'h12 == vpageFillTLB ? 1'h1 : tlb_18_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_51 = 5'h13 == vpageFillTLB ? 1'h1 : tlb_19_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_52 = 5'h14 == vpageFillTLB ? 1'h1 : tlb_20_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_53 = 5'h15 == vpageFillTLB ? 1'h1 : tlb_21_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_54 = 5'h16 == vpageFillTLB ? 1'h1 : tlb_22_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_55 = 5'h17 == vpageFillTLB ? 1'h1 : tlb_23_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_56 = 5'h18 == vpageFillTLB ? 1'h1 : tlb_24_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_57 = 5'h19 == vpageFillTLB ? 1'h1 : tlb_25_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_58 = 5'h1a == vpageFillTLB ? 1'h1 : tlb_26_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_59 = 5'h1b == vpageFillTLB ? 1'h1 : tlb_27_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_60 = 5'h1c == vpageFillTLB ? 1'h1 : tlb_28_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_61 = 5'h1d == vpageFillTLB ? 1'h1 : tlb_29_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_62 = 5'h1e == vpageFillTLB ? 1'h1 : tlb_30_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_63 = 5'h1f == vpageFillTLB ? 1'h1 : tlb_31_valid; // @[TLB.scala 38:29:@534.6]
  assign _GEN_64 = io_fill ? _GEN_0 : tlb_0_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_65 = io_fill ? _GEN_1 : tlb_1_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_66 = io_fill ? _GEN_2 : tlb_2_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_67 = io_fill ? _GEN_3 : tlb_3_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_68 = io_fill ? _GEN_4 : tlb_4_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_69 = io_fill ? _GEN_5 : tlb_5_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_70 = io_fill ? _GEN_6 : tlb_6_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_71 = io_fill ? _GEN_7 : tlb_7_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_72 = io_fill ? _GEN_8 : tlb_8_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_73 = io_fill ? _GEN_9 : tlb_9_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_74 = io_fill ? _GEN_10 : tlb_10_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_75 = io_fill ? _GEN_11 : tlb_11_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_76 = io_fill ? _GEN_12 : tlb_12_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_77 = io_fill ? _GEN_13 : tlb_13_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_78 = io_fill ? _GEN_14 : tlb_14_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_79 = io_fill ? _GEN_15 : tlb_15_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_80 = io_fill ? _GEN_16 : tlb_16_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_81 = io_fill ? _GEN_17 : tlb_17_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_82 = io_fill ? _GEN_18 : tlb_18_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_83 = io_fill ? _GEN_19 : tlb_19_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_84 = io_fill ? _GEN_20 : tlb_20_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_85 = io_fill ? _GEN_21 : tlb_21_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_86 = io_fill ? _GEN_22 : tlb_22_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_87 = io_fill ? _GEN_23 : tlb_23_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_88 = io_fill ? _GEN_24 : tlb_24_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_89 = io_fill ? _GEN_25 : tlb_25_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_90 = io_fill ? _GEN_26 : tlb_26_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_91 = io_fill ? _GEN_27 : tlb_27_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_92 = io_fill ? _GEN_28 : tlb_28_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_93 = io_fill ? _GEN_29 : tlb_29_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_94 = io_fill ? _GEN_30 : tlb_30_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_95 = io_fill ? _GEN_31 : tlb_31_bits; // @[TLB.scala 36:17:@532.4]
  assign _GEN_96 = io_fill ? _GEN_32 : tlb_0_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_97 = io_fill ? _GEN_33 : tlb_1_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_98 = io_fill ? _GEN_34 : tlb_2_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_99 = io_fill ? _GEN_35 : tlb_3_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_100 = io_fill ? _GEN_36 : tlb_4_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_101 = io_fill ? _GEN_37 : tlb_5_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_102 = io_fill ? _GEN_38 : tlb_6_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_103 = io_fill ? _GEN_39 : tlb_7_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_104 = io_fill ? _GEN_40 : tlb_8_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_105 = io_fill ? _GEN_41 : tlb_9_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_106 = io_fill ? _GEN_42 : tlb_10_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_107 = io_fill ? _GEN_43 : tlb_11_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_108 = io_fill ? _GEN_44 : tlb_12_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_109 = io_fill ? _GEN_45 : tlb_13_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_110 = io_fill ? _GEN_46 : tlb_14_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_111 = io_fill ? _GEN_47 : tlb_15_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_112 = io_fill ? _GEN_48 : tlb_16_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_113 = io_fill ? _GEN_49 : tlb_17_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_114 = io_fill ? _GEN_50 : tlb_18_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_115 = io_fill ? _GEN_51 : tlb_19_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_116 = io_fill ? _GEN_52 : tlb_20_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_117 = io_fill ? _GEN_53 : tlb_21_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_118 = io_fill ? _GEN_54 : tlb_22_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_119 = io_fill ? _GEN_55 : tlb_23_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_120 = io_fill ? _GEN_56 : tlb_24_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_121 = io_fill ? _GEN_57 : tlb_25_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_122 = io_fill ? _GEN_58 : tlb_26_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_123 = io_fill ? _GEN_59 : tlb_27_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_124 = io_fill ? _GEN_60 : tlb_28_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_125 = io_fill ? _GEN_61 : tlb_29_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_126 = io_fill ? _GEN_62 : tlb_30_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_127 = io_fill ? _GEN_63 : tlb_31_valid; // @[TLB.scala 36:17:@532.4]
  assign _GEN_130 = 5'h1 == vpageTLB ? tlb_1_valid : tlb_0_valid; // @[TLB.scala 41:56:@536.4]
  assign _GEN_131 = 5'h1 == vpageTLB ? tlb_1_bits : tlb_0_bits; // @[TLB.scala 41:56:@536.4]
  assign _GEN_132 = 5'h2 == vpageTLB ? tlb_2_valid : _GEN_130; // @[TLB.scala 41:56:@536.4]
  assign _GEN_133 = 5'h2 == vpageTLB ? tlb_2_bits : _GEN_131; // @[TLB.scala 41:56:@536.4]
  assign _GEN_134 = 5'h3 == vpageTLB ? tlb_3_valid : _GEN_132; // @[TLB.scala 41:56:@536.4]
  assign _GEN_135 = 5'h3 == vpageTLB ? tlb_3_bits : _GEN_133; // @[TLB.scala 41:56:@536.4]
  assign _GEN_136 = 5'h4 == vpageTLB ? tlb_4_valid : _GEN_134; // @[TLB.scala 41:56:@536.4]
  assign _GEN_137 = 5'h4 == vpageTLB ? tlb_4_bits : _GEN_135; // @[TLB.scala 41:56:@536.4]
  assign _GEN_138 = 5'h5 == vpageTLB ? tlb_5_valid : _GEN_136; // @[TLB.scala 41:56:@536.4]
  assign _GEN_139 = 5'h5 == vpageTLB ? tlb_5_bits : _GEN_137; // @[TLB.scala 41:56:@536.4]
  assign _GEN_140 = 5'h6 == vpageTLB ? tlb_6_valid : _GEN_138; // @[TLB.scala 41:56:@536.4]
  assign _GEN_141 = 5'h6 == vpageTLB ? tlb_6_bits : _GEN_139; // @[TLB.scala 41:56:@536.4]
  assign _GEN_142 = 5'h7 == vpageTLB ? tlb_7_valid : _GEN_140; // @[TLB.scala 41:56:@536.4]
  assign _GEN_143 = 5'h7 == vpageTLB ? tlb_7_bits : _GEN_141; // @[TLB.scala 41:56:@536.4]
  assign _GEN_144 = 5'h8 == vpageTLB ? tlb_8_valid : _GEN_142; // @[TLB.scala 41:56:@536.4]
  assign _GEN_145 = 5'h8 == vpageTLB ? tlb_8_bits : _GEN_143; // @[TLB.scala 41:56:@536.4]
  assign _GEN_146 = 5'h9 == vpageTLB ? tlb_9_valid : _GEN_144; // @[TLB.scala 41:56:@536.4]
  assign _GEN_147 = 5'h9 == vpageTLB ? tlb_9_bits : _GEN_145; // @[TLB.scala 41:56:@536.4]
  assign _GEN_148 = 5'ha == vpageTLB ? tlb_10_valid : _GEN_146; // @[TLB.scala 41:56:@536.4]
  assign _GEN_149 = 5'ha == vpageTLB ? tlb_10_bits : _GEN_147; // @[TLB.scala 41:56:@536.4]
  assign _GEN_150 = 5'hb == vpageTLB ? tlb_11_valid : _GEN_148; // @[TLB.scala 41:56:@536.4]
  assign _GEN_151 = 5'hb == vpageTLB ? tlb_11_bits : _GEN_149; // @[TLB.scala 41:56:@536.4]
  assign _GEN_152 = 5'hc == vpageTLB ? tlb_12_valid : _GEN_150; // @[TLB.scala 41:56:@536.4]
  assign _GEN_153 = 5'hc == vpageTLB ? tlb_12_bits : _GEN_151; // @[TLB.scala 41:56:@536.4]
  assign _GEN_154 = 5'hd == vpageTLB ? tlb_13_valid : _GEN_152; // @[TLB.scala 41:56:@536.4]
  assign _GEN_155 = 5'hd == vpageTLB ? tlb_13_bits : _GEN_153; // @[TLB.scala 41:56:@536.4]
  assign _GEN_156 = 5'he == vpageTLB ? tlb_14_valid : _GEN_154; // @[TLB.scala 41:56:@536.4]
  assign _GEN_157 = 5'he == vpageTLB ? tlb_14_bits : _GEN_155; // @[TLB.scala 41:56:@536.4]
  assign _GEN_158 = 5'hf == vpageTLB ? tlb_15_valid : _GEN_156; // @[TLB.scala 41:56:@536.4]
  assign _GEN_159 = 5'hf == vpageTLB ? tlb_15_bits : _GEN_157; // @[TLB.scala 41:56:@536.4]
  assign _GEN_160 = 5'h10 == vpageTLB ? tlb_16_valid : _GEN_158; // @[TLB.scala 41:56:@536.4]
  assign _GEN_161 = 5'h10 == vpageTLB ? tlb_16_bits : _GEN_159; // @[TLB.scala 41:56:@536.4]
  assign _GEN_162 = 5'h11 == vpageTLB ? tlb_17_valid : _GEN_160; // @[TLB.scala 41:56:@536.4]
  assign _GEN_163 = 5'h11 == vpageTLB ? tlb_17_bits : _GEN_161; // @[TLB.scala 41:56:@536.4]
  assign _GEN_164 = 5'h12 == vpageTLB ? tlb_18_valid : _GEN_162; // @[TLB.scala 41:56:@536.4]
  assign _GEN_165 = 5'h12 == vpageTLB ? tlb_18_bits : _GEN_163; // @[TLB.scala 41:56:@536.4]
  assign _GEN_166 = 5'h13 == vpageTLB ? tlb_19_valid : _GEN_164; // @[TLB.scala 41:56:@536.4]
  assign _GEN_167 = 5'h13 == vpageTLB ? tlb_19_bits : _GEN_165; // @[TLB.scala 41:56:@536.4]
  assign _GEN_168 = 5'h14 == vpageTLB ? tlb_20_valid : _GEN_166; // @[TLB.scala 41:56:@536.4]
  assign _GEN_169 = 5'h14 == vpageTLB ? tlb_20_bits : _GEN_167; // @[TLB.scala 41:56:@536.4]
  assign _GEN_170 = 5'h15 == vpageTLB ? tlb_21_valid : _GEN_168; // @[TLB.scala 41:56:@536.4]
  assign _GEN_171 = 5'h15 == vpageTLB ? tlb_21_bits : _GEN_169; // @[TLB.scala 41:56:@536.4]
  assign _GEN_172 = 5'h16 == vpageTLB ? tlb_22_valid : _GEN_170; // @[TLB.scala 41:56:@536.4]
  assign _GEN_173 = 5'h16 == vpageTLB ? tlb_22_bits : _GEN_171; // @[TLB.scala 41:56:@536.4]
  assign _GEN_174 = 5'h17 == vpageTLB ? tlb_23_valid : _GEN_172; // @[TLB.scala 41:56:@536.4]
  assign _GEN_175 = 5'h17 == vpageTLB ? tlb_23_bits : _GEN_173; // @[TLB.scala 41:56:@536.4]
  assign _GEN_176 = 5'h18 == vpageTLB ? tlb_24_valid : _GEN_174; // @[TLB.scala 41:56:@536.4]
  assign _GEN_177 = 5'h18 == vpageTLB ? tlb_24_bits : _GEN_175; // @[TLB.scala 41:56:@536.4]
  assign _GEN_178 = 5'h19 == vpageTLB ? tlb_25_valid : _GEN_176; // @[TLB.scala 41:56:@536.4]
  assign _GEN_179 = 5'h19 == vpageTLB ? tlb_25_bits : _GEN_177; // @[TLB.scala 41:56:@536.4]
  assign _GEN_180 = 5'h1a == vpageTLB ? tlb_26_valid : _GEN_178; // @[TLB.scala 41:56:@536.4]
  assign _GEN_181 = 5'h1a == vpageTLB ? tlb_26_bits : _GEN_179; // @[TLB.scala 41:56:@536.4]
  assign _GEN_182 = 5'h1b == vpageTLB ? tlb_27_valid : _GEN_180; // @[TLB.scala 41:56:@536.4]
  assign _GEN_183 = 5'h1b == vpageTLB ? tlb_27_bits : _GEN_181; // @[TLB.scala 41:56:@536.4]
  assign _GEN_184 = 5'h1c == vpageTLB ? tlb_28_valid : _GEN_182; // @[TLB.scala 41:56:@536.4]
  assign _GEN_185 = 5'h1c == vpageTLB ? tlb_28_bits : _GEN_183; // @[TLB.scala 41:56:@536.4]
  assign _GEN_186 = 5'h1d == vpageTLB ? tlb_29_valid : _GEN_184; // @[TLB.scala 41:56:@536.4]
  assign _GEN_187 = 5'h1d == vpageTLB ? tlb_29_bits : _GEN_185; // @[TLB.scala 41:56:@536.4]
  assign _GEN_188 = 5'h1e == vpageTLB ? tlb_30_valid : _GEN_186; // @[TLB.scala 41:56:@536.4]
  assign _GEN_189 = 5'h1e == vpageTLB ? tlb_30_bits : _GEN_187; // @[TLB.scala 41:56:@536.4]
  assign _GEN_190 = 5'h1f == vpageTLB ? tlb_31_valid : _GEN_188; // @[TLB.scala 41:56:@536.4]
  assign _GEN_191 = 5'h1f == vpageTLB ? tlb_31_bits : _GEN_189; // @[TLB.scala 41:56:@536.4]
  assign _T_616 = _GEN_191 == vpageTAG; // @[TLB.scala 42:55:@539.4]
  assign io_hit = _GEN_190 & _T_616; // @[TLB.scala 42:10:@541.4]
  assign io_paddr_valid = io_vaddr_valid; // @[TLB.scala 43:18:@542.4]
  assign io_paddr_bits = io_vaddr_bits >> 2'h2; // @[TLB.scala 44:17:@544.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tlb_0_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  tlb_0_bits = _RAND_1[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tlb_1_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  tlb_1_bits = _RAND_3[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  tlb_2_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  tlb_2_bits = _RAND_5[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  tlb_3_valid = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  tlb_3_bits = _RAND_7[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tlb_4_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  tlb_4_bits = _RAND_9[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tlb_5_valid = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  tlb_5_bits = _RAND_11[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  tlb_6_valid = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  tlb_6_bits = _RAND_13[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  tlb_7_valid = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  tlb_7_bits = _RAND_15[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  tlb_8_valid = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{`RANDOM}};
  tlb_8_bits = _RAND_17[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  tlb_9_valid = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  tlb_9_bits = _RAND_19[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  tlb_10_valid = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  tlb_10_bits = _RAND_21[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  tlb_11_valid = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{`RANDOM}};
  tlb_11_bits = _RAND_23[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  tlb_12_valid = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  tlb_12_bits = _RAND_25[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  tlb_13_valid = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  tlb_13_bits = _RAND_27[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  tlb_14_valid = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  tlb_14_bits = _RAND_29[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  tlb_15_valid = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  tlb_15_bits = _RAND_31[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  tlb_16_valid = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  tlb_16_bits = _RAND_33[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  tlb_17_valid = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  tlb_17_bits = _RAND_35[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  tlb_18_valid = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  tlb_18_bits = _RAND_37[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  tlb_19_valid = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  tlb_19_bits = _RAND_39[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  tlb_20_valid = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{`RANDOM}};
  tlb_20_bits = _RAND_41[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  tlb_21_valid = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  tlb_21_bits = _RAND_43[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  tlb_22_valid = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  tlb_22_bits = _RAND_45[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  tlb_23_valid = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  tlb_23_bits = _RAND_47[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  tlb_24_valid = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  tlb_24_bits = _RAND_49[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  tlb_25_valid = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {2{`RANDOM}};
  tlb_25_bits = _RAND_51[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  tlb_26_valid = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {2{`RANDOM}};
  tlb_26_bits = _RAND_53[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  tlb_27_valid = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  tlb_27_bits = _RAND_55[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  tlb_28_valid = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  tlb_28_bits = _RAND_57[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  tlb_29_valid = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {2{`RANDOM}};
  tlb_29_bits = _RAND_59[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  tlb_30_valid = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {2{`RANDOM}};
  tlb_30_bits = _RAND_61[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  tlb_31_valid = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {2{`RANDOM}};
  tlb_31_bits = _RAND_63[48:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      tlb_0_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h0 == vpageFillTLB) begin
          tlb_0_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_0_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h0 == vpageFillTLB) begin
          tlb_0_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_1_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h1 == vpageFillTLB) begin
          tlb_1_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_1_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h1 == vpageFillTLB) begin
          tlb_1_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_2_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h2 == vpageFillTLB) begin
          tlb_2_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_2_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h2 == vpageFillTLB) begin
          tlb_2_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_3_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h3 == vpageFillTLB) begin
          tlb_3_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_3_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h3 == vpageFillTLB) begin
          tlb_3_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_4_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h4 == vpageFillTLB) begin
          tlb_4_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_4_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h4 == vpageFillTLB) begin
          tlb_4_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_5_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h5 == vpageFillTLB) begin
          tlb_5_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_5_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h5 == vpageFillTLB) begin
          tlb_5_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_6_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h6 == vpageFillTLB) begin
          tlb_6_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_6_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h6 == vpageFillTLB) begin
          tlb_6_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_7_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h7 == vpageFillTLB) begin
          tlb_7_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_7_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h7 == vpageFillTLB) begin
          tlb_7_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_8_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h8 == vpageFillTLB) begin
          tlb_8_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_8_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h8 == vpageFillTLB) begin
          tlb_8_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_9_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h9 == vpageFillTLB) begin
          tlb_9_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_9_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h9 == vpageFillTLB) begin
          tlb_9_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_10_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'ha == vpageFillTLB) begin
          tlb_10_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_10_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'ha == vpageFillTLB) begin
          tlb_10_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_11_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'hb == vpageFillTLB) begin
          tlb_11_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_11_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'hb == vpageFillTLB) begin
          tlb_11_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_12_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'hc == vpageFillTLB) begin
          tlb_12_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_12_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'hc == vpageFillTLB) begin
          tlb_12_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_13_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'hd == vpageFillTLB) begin
          tlb_13_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_13_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'hd == vpageFillTLB) begin
          tlb_13_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_14_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'he == vpageFillTLB) begin
          tlb_14_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_14_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'he == vpageFillTLB) begin
          tlb_14_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_15_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'hf == vpageFillTLB) begin
          tlb_15_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_15_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'hf == vpageFillTLB) begin
          tlb_15_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_16_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h10 == vpageFillTLB) begin
          tlb_16_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_16_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h10 == vpageFillTLB) begin
          tlb_16_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_17_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h11 == vpageFillTLB) begin
          tlb_17_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_17_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h11 == vpageFillTLB) begin
          tlb_17_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_18_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h12 == vpageFillTLB) begin
          tlb_18_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_18_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h12 == vpageFillTLB) begin
          tlb_18_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_19_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h13 == vpageFillTLB) begin
          tlb_19_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_19_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h13 == vpageFillTLB) begin
          tlb_19_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_20_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h14 == vpageFillTLB) begin
          tlb_20_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_20_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h14 == vpageFillTLB) begin
          tlb_20_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_21_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h15 == vpageFillTLB) begin
          tlb_21_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_21_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h15 == vpageFillTLB) begin
          tlb_21_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_22_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h16 == vpageFillTLB) begin
          tlb_22_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_22_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h16 == vpageFillTLB) begin
          tlb_22_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_23_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h17 == vpageFillTLB) begin
          tlb_23_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_23_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h17 == vpageFillTLB) begin
          tlb_23_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_24_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h18 == vpageFillTLB) begin
          tlb_24_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_24_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h18 == vpageFillTLB) begin
          tlb_24_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_25_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h19 == vpageFillTLB) begin
          tlb_25_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_25_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h19 == vpageFillTLB) begin
          tlb_25_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_26_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h1a == vpageFillTLB) begin
          tlb_26_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_26_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h1a == vpageFillTLB) begin
          tlb_26_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_27_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h1b == vpageFillTLB) begin
          tlb_27_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_27_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h1b == vpageFillTLB) begin
          tlb_27_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_28_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h1c == vpageFillTLB) begin
          tlb_28_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_28_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h1c == vpageFillTLB) begin
          tlb_28_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_29_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h1d == vpageFillTLB) begin
          tlb_29_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_29_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h1d == vpageFillTLB) begin
          tlb_29_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_30_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h1e == vpageFillTLB) begin
          tlb_30_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_30_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h1e == vpageFillTLB) begin
          tlb_30_bits <= vpageFillTAG;
        end
      end
    end
    if (reset) begin
      tlb_31_valid <= 1'h0;
    end else begin
      if (io_fill) begin
        if (5'h1f == vpageFillTLB) begin
          tlb_31_valid <= 1'h1;
        end
      end
    end
    if (reset) begin
      tlb_31_bits <= 49'h0;
    end else begin
      if (io_fill) begin
        if (5'h1f == vpageFillTLB) begin
          tlb_31_bits <= vpageFillTAG;
        end
      end
    end
  end
endmodule
