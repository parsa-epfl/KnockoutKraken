module CondUnit( // @[:@2776.2]
  input  [3:0] io_cond, // @[:@2779.4]
  input  [3:0] io_nzcv, // @[:@2779.4]
  output       io_res // @[:@2779.4]
);
  wire [2:0] _T_13; // @[branch.scala 22:21:@2783.4]
  wire  _T_15; // @[branch.scala 22:27:@2784.4]
  wire  _T_16; // @[branch.scala 22:60:@2786.6]
  wire  _T_21; // @[branch.scala 23:27:@2792.6]
  wire  _T_22; // @[branch.scala 23:60:@2794.8]
  wire  _T_27; // @[branch.scala 24:27:@2800.8]
  wire  _T_28; // @[branch.scala 24:60:@2802.10]
  wire  _T_33; // @[branch.scala 25:27:@2808.10]
  wire  _T_34; // @[branch.scala 25:60:@2810.12]
  wire  _T_39; // @[branch.scala 26:27:@2816.12]
  wire  _T_45; // @[branch.scala 27:27:@2824.14]
  wire  _T_51; // @[branch.scala 28:27:@2832.16]
  wire  _T_57; // @[branch.scala 29:27:@2840.18]
  wire  _GEN_1; // @[branch.scala 28:41:@2833.16]
  wire  _GEN_2; // @[branch.scala 27:41:@2825.14]
  wire  _GEN_3; // @[branch.scala 26:41:@2817.12]
  wire  _GEN_4; // @[branch.scala 25:41:@2809.10]
  wire  _GEN_5; // @[branch.scala 24:41:@2801.8]
  wire  _GEN_6; // @[branch.scala 23:41:@2793.6]
  wire  result; // @[branch.scala 22:41:@2785.4]
  wire  _T_59; // @[branch.scala 31:15:@2844.4]
  wire  _T_63; // @[branch.scala 31:38:@2846.4]
  wire  _T_64; // @[branch.scala 31:27:@2847.4]
  wire  _T_66; // @[branch.scala 32:15:@2849.6]
  assign _T_13 = io_cond[3:1]; // @[branch.scala 22:21:@2783.4]
  assign _T_15 = _T_13 == 3'h0; // @[branch.scala 22:27:@2784.4]
  assign _T_16 = io_nzcv[2]; // @[branch.scala 22:60:@2786.6]
  assign _T_21 = _T_13 == 3'h1; // @[branch.scala 23:27:@2792.6]
  assign _T_22 = io_nzcv[1]; // @[branch.scala 23:60:@2794.8]
  assign _T_27 = _T_13 == 3'h2; // @[branch.scala 24:27:@2800.8]
  assign _T_28 = io_nzcv[3]; // @[branch.scala 24:60:@2802.10]
  assign _T_33 = _T_13 == 3'h3; // @[branch.scala 25:27:@2808.10]
  assign _T_34 = io_nzcv[0]; // @[branch.scala 25:60:@2810.12]
  assign _T_39 = _T_13 == 3'h4; // @[branch.scala 26:27:@2816.12]
  assign _T_45 = _T_13 == 3'h5; // @[branch.scala 27:27:@2824.14]
  assign _T_51 = _T_13 == 3'h6; // @[branch.scala 28:27:@2832.16]
  assign _T_57 = _T_13 == 3'h7; // @[branch.scala 29:27:@2840.18]
  assign _GEN_1 = _T_51 ? _T_28 : _T_57; // @[branch.scala 28:41:@2833.16]
  assign _GEN_2 = _T_45 ? _T_28 : _GEN_1; // @[branch.scala 27:41:@2825.14]
  assign _GEN_3 = _T_39 ? _T_22 : _GEN_2; // @[branch.scala 26:41:@2817.12]
  assign _GEN_4 = _T_33 ? _T_34 : _GEN_3; // @[branch.scala 25:41:@2809.10]
  assign _GEN_5 = _T_27 ? _T_28 : _GEN_4; // @[branch.scala 24:41:@2801.8]
  assign _GEN_6 = _T_21 ? _T_22 : _GEN_5; // @[branch.scala 23:41:@2793.6]
  assign result = _T_15 ? _T_16 : _GEN_6; // @[branch.scala 22:41:@2785.4]
  assign _T_59 = io_cond[0]; // @[branch.scala 31:15:@2844.4]
  assign _T_63 = io_cond != 4'hf; // @[branch.scala 31:38:@2846.4]
  assign _T_64 = _T_59 & _T_63; // @[branch.scala 31:27:@2847.4]
  assign _T_66 = result == 1'h0; // @[branch.scala 32:15:@2849.6]
  assign io_res = _T_64 ? _T_66 : result; // @[branch.scala 32:12:@2850.6 branch.scala 34:12:@2853.6]
endmodule
