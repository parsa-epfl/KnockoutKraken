module TLBUnit(
  input         clock,
  input         reset,
  input         io_fillTLB_valid,
  input         io_fillTLB_bits_tlbEntry_wrEn,
  input  [51:0] io_fillTLB_bits_tlbEntry_tag,
  input  [5:0]  io_fillTLB_bits_tlbIdx,
  input         io_iPort_vaddr_valid,
  input  [63:0] io_iPort_vaddr_bits,
  output [63:0] io_iPort_paddr,
  output        io_iPort_miss_valid,
  output [63:0] io_iPort_miss_bits_vaddr,
  output [5:0]  io_iPort_miss_bits_tlbIdx,
  input         io_dPort_vaddr_valid,
  input  [63:0] io_dPort_vaddr_bits,
  output [63:0] io_dPort_paddr,
  output        io_dPort_miss_valid,
  output [63:0] io_dPort_miss_bits_vaddr,
  output [5:0]  io_dPort_miss_bits_tlbIdx
);
  reg [53:0] tlb [0:63]; // @[TLB.scala 53:16]
  reg [63:0] _RAND_0;
  wire [53:0] tlb__T_4_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_4_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_16_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_16_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_28_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_28_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_40_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_40_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_52_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_52_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_64_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_64_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_76_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_76_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_88_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_88_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_100_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_100_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_112_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_112_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_124_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_124_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_136_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_136_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_148_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_148_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_160_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_160_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_172_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_172_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_184_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_184_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_196_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_196_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_208_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_208_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_220_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_220_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_232_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_232_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_244_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_244_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_256_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_256_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_268_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_268_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_280_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_280_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_292_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_292_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_304_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_304_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_316_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_316_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_328_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_328_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_340_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_340_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_352_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_352_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_364_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_364_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_376_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_376_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_388_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_388_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_400_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_400_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_412_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_412_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_424_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_424_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_436_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_436_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_448_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_448_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_460_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_460_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_472_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_472_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_484_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_484_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_496_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_496_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_508_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_508_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_520_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_520_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_532_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_532_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_544_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_544_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_556_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_556_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_568_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_568_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_580_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_580_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_592_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_592_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_604_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_604_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_616_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_616_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_628_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_628_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_640_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_640_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_652_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_652_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_664_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_664_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_676_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_676_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_688_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_688_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_700_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_700_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_712_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_712_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_724_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_724_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_736_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_736_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_748_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_748_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_760_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_760_addr; // @[TLB.scala 53:16]
  wire [53:0] tlb__T_788_data; // @[TLB.scala 53:16]
  wire [5:0] tlb__T_788_addr; // @[TLB.scala 53:16]
  wire  tlb__T_788_mask; // @[TLB.scala 53:16]
  wire  tlb__T_788_en; // @[TLB.scala 53:16]
  wire  lru_clock; // @[TLB.scala 81:19]
  wire  lru_reset; // @[TLB.scala 81:19]
  wire  lru_io_idx_1_valid; // @[TLB.scala 81:19]
  wire [5:0] lru_io_idx_1_bits; // @[TLB.scala 81:19]
  wire  lru_io_idx_2_valid; // @[TLB.scala 81:19]
  wire [5:0] lru_io_idx_2_bits; // @[TLB.scala 81:19]
  wire [5:0] lru_io_lru_idx; // @[TLB.scala 81:19]
  wire [1:0] _T; // @[TLB.scala 53:60]
  wire [51:0] iPortTagIn; // @[TLB.scala 12:9]
  wire [51:0] dPortTagIn; // @[TLB.scala 12:9]
  wire [53:0] _T_6;
  wire  _T_10; // @[TLB.scala 68:25]
  wire  _T_13; // @[TLB.scala 73:25]
  wire  _GEN_7; // @[TLB.scala 67:26]
  wire  _GEN_10; // @[TLB.scala 67:26]
  wire [53:0] _T_18;
  wire  _T_22; // @[TLB.scala 68:25]
  wire [5:0] _GEN_12; // @[TLB.scala 68:41]
  wire  _GEN_13; // @[TLB.scala 68:41]
  wire  _T_25; // @[TLB.scala 73:25]
  wire [5:0] _GEN_15; // @[TLB.scala 73:41]
  wire  _GEN_16; // @[TLB.scala 73:41]
  wire [5:0] _GEN_18; // @[TLB.scala 67:26]
  wire  _GEN_19; // @[TLB.scala 67:26]
  wire [5:0] _GEN_21; // @[TLB.scala 67:26]
  wire  _GEN_22; // @[TLB.scala 67:26]
  wire [53:0] _T_30;
  wire  _T_34; // @[TLB.scala 68:25]
  wire [5:0] _GEN_24; // @[TLB.scala 68:41]
  wire  _GEN_25; // @[TLB.scala 68:41]
  wire  _T_37; // @[TLB.scala 73:25]
  wire [5:0] _GEN_27; // @[TLB.scala 73:41]
  wire  _GEN_28; // @[TLB.scala 73:41]
  wire [5:0] _GEN_30; // @[TLB.scala 67:26]
  wire  _GEN_31; // @[TLB.scala 67:26]
  wire [5:0] _GEN_33; // @[TLB.scala 67:26]
  wire  _GEN_34; // @[TLB.scala 67:26]
  wire [53:0] _T_42;
  wire  _T_46; // @[TLB.scala 68:25]
  wire [5:0] _GEN_36; // @[TLB.scala 68:41]
  wire  _GEN_37; // @[TLB.scala 68:41]
  wire  _T_49; // @[TLB.scala 73:25]
  wire [5:0] _GEN_39; // @[TLB.scala 73:41]
  wire  _GEN_40; // @[TLB.scala 73:41]
  wire [5:0] _GEN_42; // @[TLB.scala 67:26]
  wire  _GEN_43; // @[TLB.scala 67:26]
  wire [5:0] _GEN_45; // @[TLB.scala 67:26]
  wire  _GEN_46; // @[TLB.scala 67:26]
  wire [53:0] _T_54;
  wire  _T_58; // @[TLB.scala 68:25]
  wire [5:0] _GEN_48; // @[TLB.scala 68:41]
  wire  _GEN_49; // @[TLB.scala 68:41]
  wire  _T_61; // @[TLB.scala 73:25]
  wire [5:0] _GEN_51; // @[TLB.scala 73:41]
  wire  _GEN_52; // @[TLB.scala 73:41]
  wire [5:0] _GEN_54; // @[TLB.scala 67:26]
  wire  _GEN_55; // @[TLB.scala 67:26]
  wire [5:0] _GEN_57; // @[TLB.scala 67:26]
  wire  _GEN_58; // @[TLB.scala 67:26]
  wire [53:0] _T_66;
  wire  _T_70; // @[TLB.scala 68:25]
  wire [5:0] _GEN_60; // @[TLB.scala 68:41]
  wire  _GEN_61; // @[TLB.scala 68:41]
  wire  _T_73; // @[TLB.scala 73:25]
  wire [5:0] _GEN_63; // @[TLB.scala 73:41]
  wire  _GEN_64; // @[TLB.scala 73:41]
  wire [5:0] _GEN_66; // @[TLB.scala 67:26]
  wire  _GEN_67; // @[TLB.scala 67:26]
  wire [5:0] _GEN_69; // @[TLB.scala 67:26]
  wire  _GEN_70; // @[TLB.scala 67:26]
  wire [53:0] _T_78;
  wire  _T_82; // @[TLB.scala 68:25]
  wire [5:0] _GEN_72; // @[TLB.scala 68:41]
  wire  _GEN_73; // @[TLB.scala 68:41]
  wire  _T_85; // @[TLB.scala 73:25]
  wire [5:0] _GEN_75; // @[TLB.scala 73:41]
  wire  _GEN_76; // @[TLB.scala 73:41]
  wire [5:0] _GEN_78; // @[TLB.scala 67:26]
  wire  _GEN_79; // @[TLB.scala 67:26]
  wire [5:0] _GEN_81; // @[TLB.scala 67:26]
  wire  _GEN_82; // @[TLB.scala 67:26]
  wire [53:0] _T_90;
  wire  _T_94; // @[TLB.scala 68:25]
  wire [5:0] _GEN_84; // @[TLB.scala 68:41]
  wire  _GEN_85; // @[TLB.scala 68:41]
  wire  _T_97; // @[TLB.scala 73:25]
  wire [5:0] _GEN_87; // @[TLB.scala 73:41]
  wire  _GEN_88; // @[TLB.scala 73:41]
  wire [5:0] _GEN_90; // @[TLB.scala 67:26]
  wire  _GEN_91; // @[TLB.scala 67:26]
  wire [5:0] _GEN_93; // @[TLB.scala 67:26]
  wire  _GEN_94; // @[TLB.scala 67:26]
  wire [53:0] _T_102;
  wire  _T_106; // @[TLB.scala 68:25]
  wire [5:0] _GEN_96; // @[TLB.scala 68:41]
  wire  _GEN_97; // @[TLB.scala 68:41]
  wire  _T_109; // @[TLB.scala 73:25]
  wire [5:0] _GEN_99; // @[TLB.scala 73:41]
  wire  _GEN_100; // @[TLB.scala 73:41]
  wire [5:0] _GEN_102; // @[TLB.scala 67:26]
  wire  _GEN_103; // @[TLB.scala 67:26]
  wire [5:0] _GEN_105; // @[TLB.scala 67:26]
  wire  _GEN_106; // @[TLB.scala 67:26]
  wire [53:0] _T_114;
  wire  _T_118; // @[TLB.scala 68:25]
  wire [5:0] _GEN_108; // @[TLB.scala 68:41]
  wire  _GEN_109; // @[TLB.scala 68:41]
  wire  _T_121; // @[TLB.scala 73:25]
  wire [5:0] _GEN_111; // @[TLB.scala 73:41]
  wire  _GEN_112; // @[TLB.scala 73:41]
  wire [5:0] _GEN_114; // @[TLB.scala 67:26]
  wire  _GEN_115; // @[TLB.scala 67:26]
  wire [5:0] _GEN_117; // @[TLB.scala 67:26]
  wire  _GEN_118; // @[TLB.scala 67:26]
  wire [53:0] _T_126;
  wire  _T_130; // @[TLB.scala 68:25]
  wire [5:0] _GEN_120; // @[TLB.scala 68:41]
  wire  _GEN_121; // @[TLB.scala 68:41]
  wire  _T_133; // @[TLB.scala 73:25]
  wire [5:0] _GEN_123; // @[TLB.scala 73:41]
  wire  _GEN_124; // @[TLB.scala 73:41]
  wire [5:0] _GEN_126; // @[TLB.scala 67:26]
  wire  _GEN_127; // @[TLB.scala 67:26]
  wire [5:0] _GEN_129; // @[TLB.scala 67:26]
  wire  _GEN_130; // @[TLB.scala 67:26]
  wire [53:0] _T_138;
  wire  _T_142; // @[TLB.scala 68:25]
  wire [5:0] _GEN_132; // @[TLB.scala 68:41]
  wire  _GEN_133; // @[TLB.scala 68:41]
  wire  _T_145; // @[TLB.scala 73:25]
  wire [5:0] _GEN_135; // @[TLB.scala 73:41]
  wire  _GEN_136; // @[TLB.scala 73:41]
  wire [5:0] _GEN_138; // @[TLB.scala 67:26]
  wire  _GEN_139; // @[TLB.scala 67:26]
  wire [5:0] _GEN_141; // @[TLB.scala 67:26]
  wire  _GEN_142; // @[TLB.scala 67:26]
  wire [53:0] _T_150;
  wire  _T_154; // @[TLB.scala 68:25]
  wire [5:0] _GEN_144; // @[TLB.scala 68:41]
  wire  _GEN_145; // @[TLB.scala 68:41]
  wire  _T_157; // @[TLB.scala 73:25]
  wire [5:0] _GEN_147; // @[TLB.scala 73:41]
  wire  _GEN_148; // @[TLB.scala 73:41]
  wire [5:0] _GEN_150; // @[TLB.scala 67:26]
  wire  _GEN_151; // @[TLB.scala 67:26]
  wire [5:0] _GEN_153; // @[TLB.scala 67:26]
  wire  _GEN_154; // @[TLB.scala 67:26]
  wire [53:0] _T_162;
  wire  _T_166; // @[TLB.scala 68:25]
  wire [5:0] _GEN_156; // @[TLB.scala 68:41]
  wire  _GEN_157; // @[TLB.scala 68:41]
  wire  _T_169; // @[TLB.scala 73:25]
  wire [5:0] _GEN_159; // @[TLB.scala 73:41]
  wire  _GEN_160; // @[TLB.scala 73:41]
  wire [5:0] _GEN_162; // @[TLB.scala 67:26]
  wire  _GEN_163; // @[TLB.scala 67:26]
  wire [5:0] _GEN_165; // @[TLB.scala 67:26]
  wire  _GEN_166; // @[TLB.scala 67:26]
  wire [53:0] _T_174;
  wire  _T_178; // @[TLB.scala 68:25]
  wire [5:0] _GEN_168; // @[TLB.scala 68:41]
  wire  _GEN_169; // @[TLB.scala 68:41]
  wire  _T_181; // @[TLB.scala 73:25]
  wire [5:0] _GEN_171; // @[TLB.scala 73:41]
  wire  _GEN_172; // @[TLB.scala 73:41]
  wire [5:0] _GEN_174; // @[TLB.scala 67:26]
  wire  _GEN_175; // @[TLB.scala 67:26]
  wire [5:0] _GEN_177; // @[TLB.scala 67:26]
  wire  _GEN_178; // @[TLB.scala 67:26]
  wire [53:0] _T_186;
  wire  _T_190; // @[TLB.scala 68:25]
  wire [5:0] _GEN_180; // @[TLB.scala 68:41]
  wire  _GEN_181; // @[TLB.scala 68:41]
  wire  _T_193; // @[TLB.scala 73:25]
  wire [5:0] _GEN_183; // @[TLB.scala 73:41]
  wire  _GEN_184; // @[TLB.scala 73:41]
  wire [5:0] _GEN_186; // @[TLB.scala 67:26]
  wire  _GEN_187; // @[TLB.scala 67:26]
  wire [5:0] _GEN_189; // @[TLB.scala 67:26]
  wire  _GEN_190; // @[TLB.scala 67:26]
  wire [53:0] _T_198;
  wire  _T_202; // @[TLB.scala 68:25]
  wire [5:0] _GEN_192; // @[TLB.scala 68:41]
  wire  _GEN_193; // @[TLB.scala 68:41]
  wire  _T_205; // @[TLB.scala 73:25]
  wire [5:0] _GEN_195; // @[TLB.scala 73:41]
  wire  _GEN_196; // @[TLB.scala 73:41]
  wire [5:0] _GEN_198; // @[TLB.scala 67:26]
  wire  _GEN_199; // @[TLB.scala 67:26]
  wire [5:0] _GEN_201; // @[TLB.scala 67:26]
  wire  _GEN_202; // @[TLB.scala 67:26]
  wire [53:0] _T_210;
  wire  _T_214; // @[TLB.scala 68:25]
  wire [5:0] _GEN_204; // @[TLB.scala 68:41]
  wire  _GEN_205; // @[TLB.scala 68:41]
  wire  _T_217; // @[TLB.scala 73:25]
  wire [5:0] _GEN_207; // @[TLB.scala 73:41]
  wire  _GEN_208; // @[TLB.scala 73:41]
  wire [5:0] _GEN_210; // @[TLB.scala 67:26]
  wire  _GEN_211; // @[TLB.scala 67:26]
  wire [5:0] _GEN_213; // @[TLB.scala 67:26]
  wire  _GEN_214; // @[TLB.scala 67:26]
  wire [53:0] _T_222;
  wire  _T_226; // @[TLB.scala 68:25]
  wire [5:0] _GEN_216; // @[TLB.scala 68:41]
  wire  _GEN_217; // @[TLB.scala 68:41]
  wire  _T_229; // @[TLB.scala 73:25]
  wire [5:0] _GEN_219; // @[TLB.scala 73:41]
  wire  _GEN_220; // @[TLB.scala 73:41]
  wire [5:0] _GEN_222; // @[TLB.scala 67:26]
  wire  _GEN_223; // @[TLB.scala 67:26]
  wire [5:0] _GEN_225; // @[TLB.scala 67:26]
  wire  _GEN_226; // @[TLB.scala 67:26]
  wire [53:0] _T_234;
  wire  _T_238; // @[TLB.scala 68:25]
  wire [5:0] _GEN_228; // @[TLB.scala 68:41]
  wire  _GEN_229; // @[TLB.scala 68:41]
  wire  _T_241; // @[TLB.scala 73:25]
  wire [5:0] _GEN_231; // @[TLB.scala 73:41]
  wire  _GEN_232; // @[TLB.scala 73:41]
  wire [5:0] _GEN_234; // @[TLB.scala 67:26]
  wire  _GEN_235; // @[TLB.scala 67:26]
  wire [5:0] _GEN_237; // @[TLB.scala 67:26]
  wire  _GEN_238; // @[TLB.scala 67:26]
  wire [53:0] _T_246;
  wire  _T_250; // @[TLB.scala 68:25]
  wire [5:0] _GEN_240; // @[TLB.scala 68:41]
  wire  _GEN_241; // @[TLB.scala 68:41]
  wire  _T_253; // @[TLB.scala 73:25]
  wire [5:0] _GEN_243; // @[TLB.scala 73:41]
  wire  _GEN_244; // @[TLB.scala 73:41]
  wire [5:0] _GEN_246; // @[TLB.scala 67:26]
  wire  _GEN_247; // @[TLB.scala 67:26]
  wire [5:0] _GEN_249; // @[TLB.scala 67:26]
  wire  _GEN_250; // @[TLB.scala 67:26]
  wire [53:0] _T_258;
  wire  _T_262; // @[TLB.scala 68:25]
  wire [5:0] _GEN_252; // @[TLB.scala 68:41]
  wire  _GEN_253; // @[TLB.scala 68:41]
  wire  _T_265; // @[TLB.scala 73:25]
  wire [5:0] _GEN_255; // @[TLB.scala 73:41]
  wire  _GEN_256; // @[TLB.scala 73:41]
  wire [5:0] _GEN_258; // @[TLB.scala 67:26]
  wire  _GEN_259; // @[TLB.scala 67:26]
  wire [5:0] _GEN_261; // @[TLB.scala 67:26]
  wire  _GEN_262; // @[TLB.scala 67:26]
  wire [53:0] _T_270;
  wire  _T_274; // @[TLB.scala 68:25]
  wire [5:0] _GEN_264; // @[TLB.scala 68:41]
  wire  _GEN_265; // @[TLB.scala 68:41]
  wire  _T_277; // @[TLB.scala 73:25]
  wire [5:0] _GEN_267; // @[TLB.scala 73:41]
  wire  _GEN_268; // @[TLB.scala 73:41]
  wire [5:0] _GEN_270; // @[TLB.scala 67:26]
  wire  _GEN_271; // @[TLB.scala 67:26]
  wire [5:0] _GEN_273; // @[TLB.scala 67:26]
  wire  _GEN_274; // @[TLB.scala 67:26]
  wire [53:0] _T_282;
  wire  _T_286; // @[TLB.scala 68:25]
  wire [5:0] _GEN_276; // @[TLB.scala 68:41]
  wire  _GEN_277; // @[TLB.scala 68:41]
  wire  _T_289; // @[TLB.scala 73:25]
  wire [5:0] _GEN_279; // @[TLB.scala 73:41]
  wire  _GEN_280; // @[TLB.scala 73:41]
  wire [5:0] _GEN_282; // @[TLB.scala 67:26]
  wire  _GEN_283; // @[TLB.scala 67:26]
  wire [5:0] _GEN_285; // @[TLB.scala 67:26]
  wire  _GEN_286; // @[TLB.scala 67:26]
  wire [53:0] _T_294;
  wire  _T_298; // @[TLB.scala 68:25]
  wire [5:0] _GEN_288; // @[TLB.scala 68:41]
  wire  _GEN_289; // @[TLB.scala 68:41]
  wire  _T_301; // @[TLB.scala 73:25]
  wire [5:0] _GEN_291; // @[TLB.scala 73:41]
  wire  _GEN_292; // @[TLB.scala 73:41]
  wire [5:0] _GEN_294; // @[TLB.scala 67:26]
  wire  _GEN_295; // @[TLB.scala 67:26]
  wire [5:0] _GEN_297; // @[TLB.scala 67:26]
  wire  _GEN_298; // @[TLB.scala 67:26]
  wire [53:0] _T_306;
  wire  _T_310; // @[TLB.scala 68:25]
  wire [5:0] _GEN_300; // @[TLB.scala 68:41]
  wire  _GEN_301; // @[TLB.scala 68:41]
  wire  _T_313; // @[TLB.scala 73:25]
  wire [5:0] _GEN_303; // @[TLB.scala 73:41]
  wire  _GEN_304; // @[TLB.scala 73:41]
  wire [5:0] _GEN_306; // @[TLB.scala 67:26]
  wire  _GEN_307; // @[TLB.scala 67:26]
  wire [5:0] _GEN_309; // @[TLB.scala 67:26]
  wire  _GEN_310; // @[TLB.scala 67:26]
  wire [53:0] _T_318;
  wire  _T_322; // @[TLB.scala 68:25]
  wire [5:0] _GEN_312; // @[TLB.scala 68:41]
  wire  _GEN_313; // @[TLB.scala 68:41]
  wire  _T_325; // @[TLB.scala 73:25]
  wire [5:0] _GEN_315; // @[TLB.scala 73:41]
  wire  _GEN_316; // @[TLB.scala 73:41]
  wire [5:0] _GEN_318; // @[TLB.scala 67:26]
  wire  _GEN_319; // @[TLB.scala 67:26]
  wire [5:0] _GEN_321; // @[TLB.scala 67:26]
  wire  _GEN_322; // @[TLB.scala 67:26]
  wire [53:0] _T_330;
  wire  _T_334; // @[TLB.scala 68:25]
  wire [5:0] _GEN_324; // @[TLB.scala 68:41]
  wire  _GEN_325; // @[TLB.scala 68:41]
  wire  _T_337; // @[TLB.scala 73:25]
  wire [5:0] _GEN_327; // @[TLB.scala 73:41]
  wire  _GEN_328; // @[TLB.scala 73:41]
  wire [5:0] _GEN_330; // @[TLB.scala 67:26]
  wire  _GEN_331; // @[TLB.scala 67:26]
  wire [5:0] _GEN_333; // @[TLB.scala 67:26]
  wire  _GEN_334; // @[TLB.scala 67:26]
  wire [53:0] _T_342;
  wire  _T_346; // @[TLB.scala 68:25]
  wire [5:0] _GEN_336; // @[TLB.scala 68:41]
  wire  _GEN_337; // @[TLB.scala 68:41]
  wire  _T_349; // @[TLB.scala 73:25]
  wire [5:0] _GEN_339; // @[TLB.scala 73:41]
  wire  _GEN_340; // @[TLB.scala 73:41]
  wire [5:0] _GEN_342; // @[TLB.scala 67:26]
  wire  _GEN_343; // @[TLB.scala 67:26]
  wire [5:0] _GEN_345; // @[TLB.scala 67:26]
  wire  _GEN_346; // @[TLB.scala 67:26]
  wire [53:0] _T_354;
  wire  _T_358; // @[TLB.scala 68:25]
  wire [5:0] _GEN_348; // @[TLB.scala 68:41]
  wire  _GEN_349; // @[TLB.scala 68:41]
  wire  _T_361; // @[TLB.scala 73:25]
  wire [5:0] _GEN_351; // @[TLB.scala 73:41]
  wire  _GEN_352; // @[TLB.scala 73:41]
  wire [5:0] _GEN_354; // @[TLB.scala 67:26]
  wire  _GEN_355; // @[TLB.scala 67:26]
  wire [5:0] _GEN_357; // @[TLB.scala 67:26]
  wire  _GEN_358; // @[TLB.scala 67:26]
  wire [53:0] _T_366;
  wire  _T_370; // @[TLB.scala 68:25]
  wire [5:0] _GEN_360; // @[TLB.scala 68:41]
  wire  _GEN_361; // @[TLB.scala 68:41]
  wire  _T_373; // @[TLB.scala 73:25]
  wire [5:0] _GEN_363; // @[TLB.scala 73:41]
  wire  _GEN_364; // @[TLB.scala 73:41]
  wire [5:0] _GEN_366; // @[TLB.scala 67:26]
  wire  _GEN_367; // @[TLB.scala 67:26]
  wire [5:0] _GEN_369; // @[TLB.scala 67:26]
  wire  _GEN_370; // @[TLB.scala 67:26]
  wire [53:0] _T_378;
  wire  _T_382; // @[TLB.scala 68:25]
  wire [5:0] _GEN_372; // @[TLB.scala 68:41]
  wire  _GEN_373; // @[TLB.scala 68:41]
  wire  _T_385; // @[TLB.scala 73:25]
  wire [5:0] _GEN_375; // @[TLB.scala 73:41]
  wire  _GEN_376; // @[TLB.scala 73:41]
  wire [5:0] _GEN_378; // @[TLB.scala 67:26]
  wire  _GEN_379; // @[TLB.scala 67:26]
  wire [5:0] _GEN_381; // @[TLB.scala 67:26]
  wire  _GEN_382; // @[TLB.scala 67:26]
  wire [53:0] _T_390;
  wire  _T_394; // @[TLB.scala 68:25]
  wire [5:0] _GEN_384; // @[TLB.scala 68:41]
  wire  _GEN_385; // @[TLB.scala 68:41]
  wire  _T_397; // @[TLB.scala 73:25]
  wire [5:0] _GEN_387; // @[TLB.scala 73:41]
  wire  _GEN_388; // @[TLB.scala 73:41]
  wire [5:0] _GEN_390; // @[TLB.scala 67:26]
  wire  _GEN_391; // @[TLB.scala 67:26]
  wire [5:0] _GEN_393; // @[TLB.scala 67:26]
  wire  _GEN_394; // @[TLB.scala 67:26]
  wire [53:0] _T_402;
  wire  _T_406; // @[TLB.scala 68:25]
  wire [5:0] _GEN_396; // @[TLB.scala 68:41]
  wire  _GEN_397; // @[TLB.scala 68:41]
  wire  _T_409; // @[TLB.scala 73:25]
  wire [5:0] _GEN_399; // @[TLB.scala 73:41]
  wire  _GEN_400; // @[TLB.scala 73:41]
  wire [5:0] _GEN_402; // @[TLB.scala 67:26]
  wire  _GEN_403; // @[TLB.scala 67:26]
  wire [5:0] _GEN_405; // @[TLB.scala 67:26]
  wire  _GEN_406; // @[TLB.scala 67:26]
  wire [53:0] _T_414;
  wire  _T_418; // @[TLB.scala 68:25]
  wire [5:0] _GEN_408; // @[TLB.scala 68:41]
  wire  _GEN_409; // @[TLB.scala 68:41]
  wire  _T_421; // @[TLB.scala 73:25]
  wire [5:0] _GEN_411; // @[TLB.scala 73:41]
  wire  _GEN_412; // @[TLB.scala 73:41]
  wire [5:0] _GEN_414; // @[TLB.scala 67:26]
  wire  _GEN_415; // @[TLB.scala 67:26]
  wire [5:0] _GEN_417; // @[TLB.scala 67:26]
  wire  _GEN_418; // @[TLB.scala 67:26]
  wire [53:0] _T_426;
  wire  _T_430; // @[TLB.scala 68:25]
  wire [5:0] _GEN_420; // @[TLB.scala 68:41]
  wire  _GEN_421; // @[TLB.scala 68:41]
  wire  _T_433; // @[TLB.scala 73:25]
  wire [5:0] _GEN_423; // @[TLB.scala 73:41]
  wire  _GEN_424; // @[TLB.scala 73:41]
  wire [5:0] _GEN_426; // @[TLB.scala 67:26]
  wire  _GEN_427; // @[TLB.scala 67:26]
  wire [5:0] _GEN_429; // @[TLB.scala 67:26]
  wire  _GEN_430; // @[TLB.scala 67:26]
  wire [53:0] _T_438;
  wire  _T_442; // @[TLB.scala 68:25]
  wire [5:0] _GEN_432; // @[TLB.scala 68:41]
  wire  _GEN_433; // @[TLB.scala 68:41]
  wire  _T_445; // @[TLB.scala 73:25]
  wire [5:0] _GEN_435; // @[TLB.scala 73:41]
  wire  _GEN_436; // @[TLB.scala 73:41]
  wire [5:0] _GEN_438; // @[TLB.scala 67:26]
  wire  _GEN_439; // @[TLB.scala 67:26]
  wire [5:0] _GEN_441; // @[TLB.scala 67:26]
  wire  _GEN_442; // @[TLB.scala 67:26]
  wire [53:0] _T_450;
  wire  _T_454; // @[TLB.scala 68:25]
  wire [5:0] _GEN_444; // @[TLB.scala 68:41]
  wire  _GEN_445; // @[TLB.scala 68:41]
  wire  _T_457; // @[TLB.scala 73:25]
  wire [5:0] _GEN_447; // @[TLB.scala 73:41]
  wire  _GEN_448; // @[TLB.scala 73:41]
  wire [5:0] _GEN_450; // @[TLB.scala 67:26]
  wire  _GEN_451; // @[TLB.scala 67:26]
  wire [5:0] _GEN_453; // @[TLB.scala 67:26]
  wire  _GEN_454; // @[TLB.scala 67:26]
  wire [53:0] _T_462;
  wire  _T_466; // @[TLB.scala 68:25]
  wire [5:0] _GEN_456; // @[TLB.scala 68:41]
  wire  _GEN_457; // @[TLB.scala 68:41]
  wire  _T_469; // @[TLB.scala 73:25]
  wire [5:0] _GEN_459; // @[TLB.scala 73:41]
  wire  _GEN_460; // @[TLB.scala 73:41]
  wire [5:0] _GEN_462; // @[TLB.scala 67:26]
  wire  _GEN_463; // @[TLB.scala 67:26]
  wire [5:0] _GEN_465; // @[TLB.scala 67:26]
  wire  _GEN_466; // @[TLB.scala 67:26]
  wire [53:0] _T_474;
  wire  _T_478; // @[TLB.scala 68:25]
  wire [5:0] _GEN_468; // @[TLB.scala 68:41]
  wire  _GEN_469; // @[TLB.scala 68:41]
  wire  _T_481; // @[TLB.scala 73:25]
  wire [5:0] _GEN_471; // @[TLB.scala 73:41]
  wire  _GEN_472; // @[TLB.scala 73:41]
  wire [5:0] _GEN_474; // @[TLB.scala 67:26]
  wire  _GEN_475; // @[TLB.scala 67:26]
  wire [5:0] _GEN_477; // @[TLB.scala 67:26]
  wire  _GEN_478; // @[TLB.scala 67:26]
  wire [53:0] _T_486;
  wire  _T_490; // @[TLB.scala 68:25]
  wire [5:0] _GEN_480; // @[TLB.scala 68:41]
  wire  _GEN_481; // @[TLB.scala 68:41]
  wire  _T_493; // @[TLB.scala 73:25]
  wire [5:0] _GEN_483; // @[TLB.scala 73:41]
  wire  _GEN_484; // @[TLB.scala 73:41]
  wire [5:0] _GEN_486; // @[TLB.scala 67:26]
  wire  _GEN_487; // @[TLB.scala 67:26]
  wire [5:0] _GEN_489; // @[TLB.scala 67:26]
  wire  _GEN_490; // @[TLB.scala 67:26]
  wire [53:0] _T_498;
  wire  _T_502; // @[TLB.scala 68:25]
  wire [5:0] _GEN_492; // @[TLB.scala 68:41]
  wire  _GEN_493; // @[TLB.scala 68:41]
  wire  _T_505; // @[TLB.scala 73:25]
  wire [5:0] _GEN_495; // @[TLB.scala 73:41]
  wire  _GEN_496; // @[TLB.scala 73:41]
  wire [5:0] _GEN_498; // @[TLB.scala 67:26]
  wire  _GEN_499; // @[TLB.scala 67:26]
  wire [5:0] _GEN_501; // @[TLB.scala 67:26]
  wire  _GEN_502; // @[TLB.scala 67:26]
  wire [53:0] _T_510;
  wire  _T_514; // @[TLB.scala 68:25]
  wire [5:0] _GEN_504; // @[TLB.scala 68:41]
  wire  _GEN_505; // @[TLB.scala 68:41]
  wire  _T_517; // @[TLB.scala 73:25]
  wire [5:0] _GEN_507; // @[TLB.scala 73:41]
  wire  _GEN_508; // @[TLB.scala 73:41]
  wire [5:0] _GEN_510; // @[TLB.scala 67:26]
  wire  _GEN_511; // @[TLB.scala 67:26]
  wire [5:0] _GEN_513; // @[TLB.scala 67:26]
  wire  _GEN_514; // @[TLB.scala 67:26]
  wire [53:0] _T_522;
  wire  _T_526; // @[TLB.scala 68:25]
  wire [5:0] _GEN_516; // @[TLB.scala 68:41]
  wire  _GEN_517; // @[TLB.scala 68:41]
  wire  _T_529; // @[TLB.scala 73:25]
  wire [5:0] _GEN_519; // @[TLB.scala 73:41]
  wire  _GEN_520; // @[TLB.scala 73:41]
  wire [5:0] _GEN_522; // @[TLB.scala 67:26]
  wire  _GEN_523; // @[TLB.scala 67:26]
  wire [5:0] _GEN_525; // @[TLB.scala 67:26]
  wire  _GEN_526; // @[TLB.scala 67:26]
  wire [53:0] _T_534;
  wire  _T_538; // @[TLB.scala 68:25]
  wire [5:0] _GEN_528; // @[TLB.scala 68:41]
  wire  _GEN_529; // @[TLB.scala 68:41]
  wire  _T_541; // @[TLB.scala 73:25]
  wire [5:0] _GEN_531; // @[TLB.scala 73:41]
  wire  _GEN_532; // @[TLB.scala 73:41]
  wire [5:0] _GEN_534; // @[TLB.scala 67:26]
  wire  _GEN_535; // @[TLB.scala 67:26]
  wire [5:0] _GEN_537; // @[TLB.scala 67:26]
  wire  _GEN_538; // @[TLB.scala 67:26]
  wire [53:0] _T_546;
  wire  _T_550; // @[TLB.scala 68:25]
  wire [5:0] _GEN_540; // @[TLB.scala 68:41]
  wire  _GEN_541; // @[TLB.scala 68:41]
  wire  _T_553; // @[TLB.scala 73:25]
  wire [5:0] _GEN_543; // @[TLB.scala 73:41]
  wire  _GEN_544; // @[TLB.scala 73:41]
  wire [5:0] _GEN_546; // @[TLB.scala 67:26]
  wire  _GEN_547; // @[TLB.scala 67:26]
  wire [5:0] _GEN_549; // @[TLB.scala 67:26]
  wire  _GEN_550; // @[TLB.scala 67:26]
  wire [53:0] _T_558;
  wire  _T_562; // @[TLB.scala 68:25]
  wire [5:0] _GEN_552; // @[TLB.scala 68:41]
  wire  _GEN_553; // @[TLB.scala 68:41]
  wire  _T_565; // @[TLB.scala 73:25]
  wire [5:0] _GEN_555; // @[TLB.scala 73:41]
  wire  _GEN_556; // @[TLB.scala 73:41]
  wire [5:0] _GEN_558; // @[TLB.scala 67:26]
  wire  _GEN_559; // @[TLB.scala 67:26]
  wire [5:0] _GEN_561; // @[TLB.scala 67:26]
  wire  _GEN_562; // @[TLB.scala 67:26]
  wire [53:0] _T_570;
  wire  _T_574; // @[TLB.scala 68:25]
  wire [5:0] _GEN_564; // @[TLB.scala 68:41]
  wire  _GEN_565; // @[TLB.scala 68:41]
  wire  _T_577; // @[TLB.scala 73:25]
  wire [5:0] _GEN_567; // @[TLB.scala 73:41]
  wire  _GEN_568; // @[TLB.scala 73:41]
  wire [5:0] _GEN_570; // @[TLB.scala 67:26]
  wire  _GEN_571; // @[TLB.scala 67:26]
  wire [5:0] _GEN_573; // @[TLB.scala 67:26]
  wire  _GEN_574; // @[TLB.scala 67:26]
  wire [53:0] _T_582;
  wire  _T_586; // @[TLB.scala 68:25]
  wire [5:0] _GEN_576; // @[TLB.scala 68:41]
  wire  _GEN_577; // @[TLB.scala 68:41]
  wire  _T_589; // @[TLB.scala 73:25]
  wire [5:0] _GEN_579; // @[TLB.scala 73:41]
  wire  _GEN_580; // @[TLB.scala 73:41]
  wire [5:0] _GEN_582; // @[TLB.scala 67:26]
  wire  _GEN_583; // @[TLB.scala 67:26]
  wire [5:0] _GEN_585; // @[TLB.scala 67:26]
  wire  _GEN_586; // @[TLB.scala 67:26]
  wire [53:0] _T_594;
  wire  _T_598; // @[TLB.scala 68:25]
  wire [5:0] _GEN_588; // @[TLB.scala 68:41]
  wire  _GEN_589; // @[TLB.scala 68:41]
  wire  _T_601; // @[TLB.scala 73:25]
  wire [5:0] _GEN_591; // @[TLB.scala 73:41]
  wire  _GEN_592; // @[TLB.scala 73:41]
  wire [5:0] _GEN_594; // @[TLB.scala 67:26]
  wire  _GEN_595; // @[TLB.scala 67:26]
  wire [5:0] _GEN_597; // @[TLB.scala 67:26]
  wire  _GEN_598; // @[TLB.scala 67:26]
  wire [53:0] _T_606;
  wire  _T_610; // @[TLB.scala 68:25]
  wire [5:0] _GEN_600; // @[TLB.scala 68:41]
  wire  _GEN_601; // @[TLB.scala 68:41]
  wire  _T_613; // @[TLB.scala 73:25]
  wire [5:0] _GEN_603; // @[TLB.scala 73:41]
  wire  _GEN_604; // @[TLB.scala 73:41]
  wire [5:0] _GEN_606; // @[TLB.scala 67:26]
  wire  _GEN_607; // @[TLB.scala 67:26]
  wire [5:0] _GEN_609; // @[TLB.scala 67:26]
  wire  _GEN_610; // @[TLB.scala 67:26]
  wire [53:0] _T_618;
  wire  _T_622; // @[TLB.scala 68:25]
  wire [5:0] _GEN_612; // @[TLB.scala 68:41]
  wire  _GEN_613; // @[TLB.scala 68:41]
  wire  _T_625; // @[TLB.scala 73:25]
  wire [5:0] _GEN_615; // @[TLB.scala 73:41]
  wire  _GEN_616; // @[TLB.scala 73:41]
  wire [5:0] _GEN_618; // @[TLB.scala 67:26]
  wire  _GEN_619; // @[TLB.scala 67:26]
  wire [5:0] _GEN_621; // @[TLB.scala 67:26]
  wire  _GEN_622; // @[TLB.scala 67:26]
  wire [53:0] _T_630;
  wire  _T_634; // @[TLB.scala 68:25]
  wire [5:0] _GEN_624; // @[TLB.scala 68:41]
  wire  _GEN_625; // @[TLB.scala 68:41]
  wire  _T_637; // @[TLB.scala 73:25]
  wire [5:0] _GEN_627; // @[TLB.scala 73:41]
  wire  _GEN_628; // @[TLB.scala 73:41]
  wire [5:0] _GEN_630; // @[TLB.scala 67:26]
  wire  _GEN_631; // @[TLB.scala 67:26]
  wire [5:0] _GEN_633; // @[TLB.scala 67:26]
  wire  _GEN_634; // @[TLB.scala 67:26]
  wire [53:0] _T_642;
  wire  _T_646; // @[TLB.scala 68:25]
  wire [5:0] _GEN_636; // @[TLB.scala 68:41]
  wire  _GEN_637; // @[TLB.scala 68:41]
  wire  _T_649; // @[TLB.scala 73:25]
  wire [5:0] _GEN_639; // @[TLB.scala 73:41]
  wire  _GEN_640; // @[TLB.scala 73:41]
  wire [5:0] _GEN_642; // @[TLB.scala 67:26]
  wire  _GEN_643; // @[TLB.scala 67:26]
  wire [5:0] _GEN_645; // @[TLB.scala 67:26]
  wire  _GEN_646; // @[TLB.scala 67:26]
  wire [53:0] _T_654;
  wire  _T_658; // @[TLB.scala 68:25]
  wire [5:0] _GEN_648; // @[TLB.scala 68:41]
  wire  _GEN_649; // @[TLB.scala 68:41]
  wire  _T_661; // @[TLB.scala 73:25]
  wire [5:0] _GEN_651; // @[TLB.scala 73:41]
  wire  _GEN_652; // @[TLB.scala 73:41]
  wire [5:0] _GEN_654; // @[TLB.scala 67:26]
  wire  _GEN_655; // @[TLB.scala 67:26]
  wire [5:0] _GEN_657; // @[TLB.scala 67:26]
  wire  _GEN_658; // @[TLB.scala 67:26]
  wire [53:0] _T_666;
  wire  _T_670; // @[TLB.scala 68:25]
  wire [5:0] _GEN_660; // @[TLB.scala 68:41]
  wire  _GEN_661; // @[TLB.scala 68:41]
  wire  _T_673; // @[TLB.scala 73:25]
  wire [5:0] _GEN_663; // @[TLB.scala 73:41]
  wire  _GEN_664; // @[TLB.scala 73:41]
  wire [5:0] _GEN_666; // @[TLB.scala 67:26]
  wire  _GEN_667; // @[TLB.scala 67:26]
  wire [5:0] _GEN_669; // @[TLB.scala 67:26]
  wire  _GEN_670; // @[TLB.scala 67:26]
  wire [53:0] _T_678;
  wire  _T_682; // @[TLB.scala 68:25]
  wire [5:0] _GEN_672; // @[TLB.scala 68:41]
  wire  _GEN_673; // @[TLB.scala 68:41]
  wire  _T_685; // @[TLB.scala 73:25]
  wire [5:0] _GEN_675; // @[TLB.scala 73:41]
  wire  _GEN_676; // @[TLB.scala 73:41]
  wire [5:0] _GEN_678; // @[TLB.scala 67:26]
  wire  _GEN_679; // @[TLB.scala 67:26]
  wire [5:0] _GEN_681; // @[TLB.scala 67:26]
  wire  _GEN_682; // @[TLB.scala 67:26]
  wire [53:0] _T_690;
  wire  _T_694; // @[TLB.scala 68:25]
  wire [5:0] _GEN_684; // @[TLB.scala 68:41]
  wire  _GEN_685; // @[TLB.scala 68:41]
  wire  _T_697; // @[TLB.scala 73:25]
  wire [5:0] _GEN_687; // @[TLB.scala 73:41]
  wire  _GEN_688; // @[TLB.scala 73:41]
  wire [5:0] _GEN_690; // @[TLB.scala 67:26]
  wire  _GEN_691; // @[TLB.scala 67:26]
  wire [5:0] _GEN_693; // @[TLB.scala 67:26]
  wire  _GEN_694; // @[TLB.scala 67:26]
  wire [53:0] _T_702;
  wire  _T_706; // @[TLB.scala 68:25]
  wire [5:0] _GEN_696; // @[TLB.scala 68:41]
  wire  _GEN_697; // @[TLB.scala 68:41]
  wire  _T_709; // @[TLB.scala 73:25]
  wire [5:0] _GEN_699; // @[TLB.scala 73:41]
  wire  _GEN_700; // @[TLB.scala 73:41]
  wire [5:0] _GEN_702; // @[TLB.scala 67:26]
  wire  _GEN_703; // @[TLB.scala 67:26]
  wire [5:0] _GEN_705; // @[TLB.scala 67:26]
  wire  _GEN_706; // @[TLB.scala 67:26]
  wire [53:0] _T_714;
  wire  _T_718; // @[TLB.scala 68:25]
  wire [5:0] _GEN_708; // @[TLB.scala 68:41]
  wire  _GEN_709; // @[TLB.scala 68:41]
  wire  _T_721; // @[TLB.scala 73:25]
  wire [5:0] _GEN_711; // @[TLB.scala 73:41]
  wire  _GEN_712; // @[TLB.scala 73:41]
  wire [5:0] _GEN_714; // @[TLB.scala 67:26]
  wire  _GEN_715; // @[TLB.scala 67:26]
  wire [5:0] _GEN_717; // @[TLB.scala 67:26]
  wire  _GEN_718; // @[TLB.scala 67:26]
  wire [53:0] _T_726;
  wire  _T_730; // @[TLB.scala 68:25]
  wire [5:0] _GEN_720; // @[TLB.scala 68:41]
  wire  _GEN_721; // @[TLB.scala 68:41]
  wire  _T_733; // @[TLB.scala 73:25]
  wire [5:0] _GEN_723; // @[TLB.scala 73:41]
  wire  _GEN_724; // @[TLB.scala 73:41]
  wire [5:0] _GEN_726; // @[TLB.scala 67:26]
  wire  _GEN_727; // @[TLB.scala 67:26]
  wire [5:0] _GEN_729; // @[TLB.scala 67:26]
  wire  _GEN_730; // @[TLB.scala 67:26]
  wire [53:0] _T_738;
  wire  _T_742; // @[TLB.scala 68:25]
  wire [5:0] _GEN_732; // @[TLB.scala 68:41]
  wire  _GEN_733; // @[TLB.scala 68:41]
  wire  _T_745; // @[TLB.scala 73:25]
  wire [5:0] _GEN_735; // @[TLB.scala 73:41]
  wire  _GEN_736; // @[TLB.scala 73:41]
  wire [5:0] _GEN_738; // @[TLB.scala 67:26]
  wire  _GEN_739; // @[TLB.scala 67:26]
  wire [5:0] _GEN_741; // @[TLB.scala 67:26]
  wire  _GEN_742; // @[TLB.scala 67:26]
  wire [53:0] _T_750;
  wire  _T_754; // @[TLB.scala 68:25]
  wire [5:0] _GEN_744; // @[TLB.scala 68:41]
  wire  _GEN_745; // @[TLB.scala 68:41]
  wire  _T_757; // @[TLB.scala 73:25]
  wire [5:0] _GEN_747; // @[TLB.scala 73:41]
  wire  _GEN_748; // @[TLB.scala 73:41]
  wire [5:0] _GEN_750; // @[TLB.scala 67:26]
  wire  _GEN_751; // @[TLB.scala 67:26]
  wire [5:0] _GEN_753; // @[TLB.scala 67:26]
  wire  _GEN_754; // @[TLB.scala 67:26]
  wire [53:0] _T_762;
  wire  _T_766; // @[TLB.scala 68:25]
  wire [5:0] _GEN_756; // @[TLB.scala 68:41]
  wire  _GEN_757; // @[TLB.scala 68:41]
  wire  _T_769; // @[TLB.scala 73:25]
  wire [5:0] _GEN_759; // @[TLB.scala 73:41]
  wire  _GEN_760; // @[TLB.scala 73:41]
  wire [5:0] iPortIdx; // @[TLB.scala 67:26]
  wire  iPortHit; // @[TLB.scala 67:26]
  wire [5:0] dPortIdx; // @[TLB.scala 67:26]
  wire  dPortHit; // @[TLB.scala 67:26]
  wire [63:0] _T_774; // @[TLB.scala 87:56]
  wire [14:0] _T_776; // @[Cat.scala 29:58]
  wire [63:0] _T_777; // @[TLB.scala 88:56]
  wire [14:0] _T_779; // @[Cat.scala 29:58]
  wire  _T_781; // @[TLB.scala 90:28]
  wire [5:0] pseudoLRU_idx2; // @[Cat.scala 29:58]
  wire  _T_784; // @[TLB.scala 95:26]
  wire  _T_786; // @[TLB.scala 96:26]
  PseudoBitmapLRU lru ( // @[TLB.scala 81:19]
    .clock(lru_clock),
    .reset(lru_reset),
    .io_idx_1_valid(lru_io_idx_1_valid),
    .io_idx_1_bits(lru_io_idx_1_bits),
    .io_idx_2_valid(lru_io_idx_2_valid),
    .io_idx_2_bits(lru_io_idx_2_bits),
    .io_lru_idx(lru_io_lru_idx)
  );
  assign tlb__T_4_addr = 6'h0;
  assign tlb__T_4_data = tlb[tlb__T_4_addr]; // @[TLB.scala 53:16]
  assign tlb__T_16_addr = 6'h1;
  assign tlb__T_16_data = tlb[tlb__T_16_addr]; // @[TLB.scala 53:16]
  assign tlb__T_28_addr = 6'h2;
  assign tlb__T_28_data = tlb[tlb__T_28_addr]; // @[TLB.scala 53:16]
  assign tlb__T_40_addr = 6'h3;
  assign tlb__T_40_data = tlb[tlb__T_40_addr]; // @[TLB.scala 53:16]
  assign tlb__T_52_addr = 6'h4;
  assign tlb__T_52_data = tlb[tlb__T_52_addr]; // @[TLB.scala 53:16]
  assign tlb__T_64_addr = 6'h5;
  assign tlb__T_64_data = tlb[tlb__T_64_addr]; // @[TLB.scala 53:16]
  assign tlb__T_76_addr = 6'h6;
  assign tlb__T_76_data = tlb[tlb__T_76_addr]; // @[TLB.scala 53:16]
  assign tlb__T_88_addr = 6'h7;
  assign tlb__T_88_data = tlb[tlb__T_88_addr]; // @[TLB.scala 53:16]
  assign tlb__T_100_addr = 6'h8;
  assign tlb__T_100_data = tlb[tlb__T_100_addr]; // @[TLB.scala 53:16]
  assign tlb__T_112_addr = 6'h9;
  assign tlb__T_112_data = tlb[tlb__T_112_addr]; // @[TLB.scala 53:16]
  assign tlb__T_124_addr = 6'ha;
  assign tlb__T_124_data = tlb[tlb__T_124_addr]; // @[TLB.scala 53:16]
  assign tlb__T_136_addr = 6'hb;
  assign tlb__T_136_data = tlb[tlb__T_136_addr]; // @[TLB.scala 53:16]
  assign tlb__T_148_addr = 6'hc;
  assign tlb__T_148_data = tlb[tlb__T_148_addr]; // @[TLB.scala 53:16]
  assign tlb__T_160_addr = 6'hd;
  assign tlb__T_160_data = tlb[tlb__T_160_addr]; // @[TLB.scala 53:16]
  assign tlb__T_172_addr = 6'he;
  assign tlb__T_172_data = tlb[tlb__T_172_addr]; // @[TLB.scala 53:16]
  assign tlb__T_184_addr = 6'hf;
  assign tlb__T_184_data = tlb[tlb__T_184_addr]; // @[TLB.scala 53:16]
  assign tlb__T_196_addr = 6'h10;
  assign tlb__T_196_data = tlb[tlb__T_196_addr]; // @[TLB.scala 53:16]
  assign tlb__T_208_addr = 6'h11;
  assign tlb__T_208_data = tlb[tlb__T_208_addr]; // @[TLB.scala 53:16]
  assign tlb__T_220_addr = 6'h12;
  assign tlb__T_220_data = tlb[tlb__T_220_addr]; // @[TLB.scala 53:16]
  assign tlb__T_232_addr = 6'h13;
  assign tlb__T_232_data = tlb[tlb__T_232_addr]; // @[TLB.scala 53:16]
  assign tlb__T_244_addr = 6'h14;
  assign tlb__T_244_data = tlb[tlb__T_244_addr]; // @[TLB.scala 53:16]
  assign tlb__T_256_addr = 6'h15;
  assign tlb__T_256_data = tlb[tlb__T_256_addr]; // @[TLB.scala 53:16]
  assign tlb__T_268_addr = 6'h16;
  assign tlb__T_268_data = tlb[tlb__T_268_addr]; // @[TLB.scala 53:16]
  assign tlb__T_280_addr = 6'h17;
  assign tlb__T_280_data = tlb[tlb__T_280_addr]; // @[TLB.scala 53:16]
  assign tlb__T_292_addr = 6'h18;
  assign tlb__T_292_data = tlb[tlb__T_292_addr]; // @[TLB.scala 53:16]
  assign tlb__T_304_addr = 6'h19;
  assign tlb__T_304_data = tlb[tlb__T_304_addr]; // @[TLB.scala 53:16]
  assign tlb__T_316_addr = 6'h1a;
  assign tlb__T_316_data = tlb[tlb__T_316_addr]; // @[TLB.scala 53:16]
  assign tlb__T_328_addr = 6'h1b;
  assign tlb__T_328_data = tlb[tlb__T_328_addr]; // @[TLB.scala 53:16]
  assign tlb__T_340_addr = 6'h1c;
  assign tlb__T_340_data = tlb[tlb__T_340_addr]; // @[TLB.scala 53:16]
  assign tlb__T_352_addr = 6'h1d;
  assign tlb__T_352_data = tlb[tlb__T_352_addr]; // @[TLB.scala 53:16]
  assign tlb__T_364_addr = 6'h1e;
  assign tlb__T_364_data = tlb[tlb__T_364_addr]; // @[TLB.scala 53:16]
  assign tlb__T_376_addr = 6'h1f;
  assign tlb__T_376_data = tlb[tlb__T_376_addr]; // @[TLB.scala 53:16]
  assign tlb__T_388_addr = 6'h20;
  assign tlb__T_388_data = tlb[tlb__T_388_addr]; // @[TLB.scala 53:16]
  assign tlb__T_400_addr = 6'h21;
  assign tlb__T_400_data = tlb[tlb__T_400_addr]; // @[TLB.scala 53:16]
  assign tlb__T_412_addr = 6'h22;
  assign tlb__T_412_data = tlb[tlb__T_412_addr]; // @[TLB.scala 53:16]
  assign tlb__T_424_addr = 6'h23;
  assign tlb__T_424_data = tlb[tlb__T_424_addr]; // @[TLB.scala 53:16]
  assign tlb__T_436_addr = 6'h24;
  assign tlb__T_436_data = tlb[tlb__T_436_addr]; // @[TLB.scala 53:16]
  assign tlb__T_448_addr = 6'h25;
  assign tlb__T_448_data = tlb[tlb__T_448_addr]; // @[TLB.scala 53:16]
  assign tlb__T_460_addr = 6'h26;
  assign tlb__T_460_data = tlb[tlb__T_460_addr]; // @[TLB.scala 53:16]
  assign tlb__T_472_addr = 6'h27;
  assign tlb__T_472_data = tlb[tlb__T_472_addr]; // @[TLB.scala 53:16]
  assign tlb__T_484_addr = 6'h28;
  assign tlb__T_484_data = tlb[tlb__T_484_addr]; // @[TLB.scala 53:16]
  assign tlb__T_496_addr = 6'h29;
  assign tlb__T_496_data = tlb[tlb__T_496_addr]; // @[TLB.scala 53:16]
  assign tlb__T_508_addr = 6'h2a;
  assign tlb__T_508_data = tlb[tlb__T_508_addr]; // @[TLB.scala 53:16]
  assign tlb__T_520_addr = 6'h2b;
  assign tlb__T_520_data = tlb[tlb__T_520_addr]; // @[TLB.scala 53:16]
  assign tlb__T_532_addr = 6'h2c;
  assign tlb__T_532_data = tlb[tlb__T_532_addr]; // @[TLB.scala 53:16]
  assign tlb__T_544_addr = 6'h2d;
  assign tlb__T_544_data = tlb[tlb__T_544_addr]; // @[TLB.scala 53:16]
  assign tlb__T_556_addr = 6'h2e;
  assign tlb__T_556_data = tlb[tlb__T_556_addr]; // @[TLB.scala 53:16]
  assign tlb__T_568_addr = 6'h2f;
  assign tlb__T_568_data = tlb[tlb__T_568_addr]; // @[TLB.scala 53:16]
  assign tlb__T_580_addr = 6'h30;
  assign tlb__T_580_data = tlb[tlb__T_580_addr]; // @[TLB.scala 53:16]
  assign tlb__T_592_addr = 6'h31;
  assign tlb__T_592_data = tlb[tlb__T_592_addr]; // @[TLB.scala 53:16]
  assign tlb__T_604_addr = 6'h32;
  assign tlb__T_604_data = tlb[tlb__T_604_addr]; // @[TLB.scala 53:16]
  assign tlb__T_616_addr = 6'h33;
  assign tlb__T_616_data = tlb[tlb__T_616_addr]; // @[TLB.scala 53:16]
  assign tlb__T_628_addr = 6'h34;
  assign tlb__T_628_data = tlb[tlb__T_628_addr]; // @[TLB.scala 53:16]
  assign tlb__T_640_addr = 6'h35;
  assign tlb__T_640_data = tlb[tlb__T_640_addr]; // @[TLB.scala 53:16]
  assign tlb__T_652_addr = 6'h36;
  assign tlb__T_652_data = tlb[tlb__T_652_addr]; // @[TLB.scala 53:16]
  assign tlb__T_664_addr = 6'h37;
  assign tlb__T_664_data = tlb[tlb__T_664_addr]; // @[TLB.scala 53:16]
  assign tlb__T_676_addr = 6'h38;
  assign tlb__T_676_data = tlb[tlb__T_676_addr]; // @[TLB.scala 53:16]
  assign tlb__T_688_addr = 6'h39;
  assign tlb__T_688_data = tlb[tlb__T_688_addr]; // @[TLB.scala 53:16]
  assign tlb__T_700_addr = 6'h3a;
  assign tlb__T_700_data = tlb[tlb__T_700_addr]; // @[TLB.scala 53:16]
  assign tlb__T_712_addr = 6'h3b;
  assign tlb__T_712_data = tlb[tlb__T_712_addr]; // @[TLB.scala 53:16]
  assign tlb__T_724_addr = 6'h3c;
  assign tlb__T_724_data = tlb[tlb__T_724_addr]; // @[TLB.scala 53:16]
  assign tlb__T_736_addr = 6'h3d;
  assign tlb__T_736_data = tlb[tlb__T_736_addr]; // @[TLB.scala 53:16]
  assign tlb__T_748_addr = 6'h3e;
  assign tlb__T_748_data = tlb[tlb__T_748_addr]; // @[TLB.scala 53:16]
  assign tlb__T_760_addr = 6'h3f;
  assign tlb__T_760_data = tlb[tlb__T_760_addr]; // @[TLB.scala 53:16]
  assign tlb__T_788_data = {_T,io_fillTLB_bits_tlbEntry_tag};
  assign tlb__T_788_addr = io_fillTLB_bits_tlbIdx;
  assign tlb__T_788_mask = 1'h1;
  assign tlb__T_788_en = io_fillTLB_valid;
  assign _T = {1'h1,io_fillTLB_bits_tlbEntry_wrEn}; // @[TLB.scala 53:60]
  assign iPortTagIn = io_iPort_vaddr_bits[63:12]; // @[TLB.scala 12:9]
  assign dPortTagIn = io_dPort_vaddr_bits[63:12]; // @[TLB.scala 12:9]
  assign _T_6 = tlb__T_4_data;
  assign _T_10 = _T_6[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _T_13 = _T_6[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_7 = _T_6[53] & _T_10; // @[TLB.scala 67:26]
  assign _GEN_10 = _T_6[53] & _T_13; // @[TLB.scala 67:26]
  assign _T_18 = tlb__T_16_data;
  assign _T_22 = _T_18[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_12 = _T_22 ? 6'h1 : 6'h0; // @[TLB.scala 68:41]
  assign _GEN_13 = _T_22 | _GEN_7; // @[TLB.scala 68:41]
  assign _T_25 = _T_18[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_15 = _T_25 ? 6'h1 : 6'h0; // @[TLB.scala 73:41]
  assign _GEN_16 = _T_25 | _GEN_10; // @[TLB.scala 73:41]
  assign _GEN_18 = _T_18[53] ? _GEN_12 : 6'h0; // @[TLB.scala 67:26]
  assign _GEN_19 = _T_18[53] ? _GEN_13 : _GEN_7; // @[TLB.scala 67:26]
  assign _GEN_21 = _T_18[53] ? _GEN_15 : 6'h0; // @[TLB.scala 67:26]
  assign _GEN_22 = _T_18[53] ? _GEN_16 : _GEN_10; // @[TLB.scala 67:26]
  assign _T_30 = tlb__T_28_data;
  assign _T_34 = _T_30[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_24 = _T_34 ? 6'h2 : _GEN_18; // @[TLB.scala 68:41]
  assign _GEN_25 = _T_34 | _GEN_19; // @[TLB.scala 68:41]
  assign _T_37 = _T_30[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_27 = _T_37 ? 6'h2 : _GEN_21; // @[TLB.scala 73:41]
  assign _GEN_28 = _T_37 | _GEN_22; // @[TLB.scala 73:41]
  assign _GEN_30 = _T_30[53] ? _GEN_24 : _GEN_18; // @[TLB.scala 67:26]
  assign _GEN_31 = _T_30[53] ? _GEN_25 : _GEN_19; // @[TLB.scala 67:26]
  assign _GEN_33 = _T_30[53] ? _GEN_27 : _GEN_21; // @[TLB.scala 67:26]
  assign _GEN_34 = _T_30[53] ? _GEN_28 : _GEN_22; // @[TLB.scala 67:26]
  assign _T_42 = tlb__T_40_data;
  assign _T_46 = _T_42[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_36 = _T_46 ? 6'h3 : _GEN_30; // @[TLB.scala 68:41]
  assign _GEN_37 = _T_46 | _GEN_31; // @[TLB.scala 68:41]
  assign _T_49 = _T_42[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_39 = _T_49 ? 6'h3 : _GEN_33; // @[TLB.scala 73:41]
  assign _GEN_40 = _T_49 | _GEN_34; // @[TLB.scala 73:41]
  assign _GEN_42 = _T_42[53] ? _GEN_36 : _GEN_30; // @[TLB.scala 67:26]
  assign _GEN_43 = _T_42[53] ? _GEN_37 : _GEN_31; // @[TLB.scala 67:26]
  assign _GEN_45 = _T_42[53] ? _GEN_39 : _GEN_33; // @[TLB.scala 67:26]
  assign _GEN_46 = _T_42[53] ? _GEN_40 : _GEN_34; // @[TLB.scala 67:26]
  assign _T_54 = tlb__T_52_data;
  assign _T_58 = _T_54[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_48 = _T_58 ? 6'h4 : _GEN_42; // @[TLB.scala 68:41]
  assign _GEN_49 = _T_58 | _GEN_43; // @[TLB.scala 68:41]
  assign _T_61 = _T_54[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_51 = _T_61 ? 6'h4 : _GEN_45; // @[TLB.scala 73:41]
  assign _GEN_52 = _T_61 | _GEN_46; // @[TLB.scala 73:41]
  assign _GEN_54 = _T_54[53] ? _GEN_48 : _GEN_42; // @[TLB.scala 67:26]
  assign _GEN_55 = _T_54[53] ? _GEN_49 : _GEN_43; // @[TLB.scala 67:26]
  assign _GEN_57 = _T_54[53] ? _GEN_51 : _GEN_45; // @[TLB.scala 67:26]
  assign _GEN_58 = _T_54[53] ? _GEN_52 : _GEN_46; // @[TLB.scala 67:26]
  assign _T_66 = tlb__T_64_data;
  assign _T_70 = _T_66[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_60 = _T_70 ? 6'h5 : _GEN_54; // @[TLB.scala 68:41]
  assign _GEN_61 = _T_70 | _GEN_55; // @[TLB.scala 68:41]
  assign _T_73 = _T_66[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_63 = _T_73 ? 6'h5 : _GEN_57; // @[TLB.scala 73:41]
  assign _GEN_64 = _T_73 | _GEN_58; // @[TLB.scala 73:41]
  assign _GEN_66 = _T_66[53] ? _GEN_60 : _GEN_54; // @[TLB.scala 67:26]
  assign _GEN_67 = _T_66[53] ? _GEN_61 : _GEN_55; // @[TLB.scala 67:26]
  assign _GEN_69 = _T_66[53] ? _GEN_63 : _GEN_57; // @[TLB.scala 67:26]
  assign _GEN_70 = _T_66[53] ? _GEN_64 : _GEN_58; // @[TLB.scala 67:26]
  assign _T_78 = tlb__T_76_data;
  assign _T_82 = _T_78[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_72 = _T_82 ? 6'h6 : _GEN_66; // @[TLB.scala 68:41]
  assign _GEN_73 = _T_82 | _GEN_67; // @[TLB.scala 68:41]
  assign _T_85 = _T_78[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_75 = _T_85 ? 6'h6 : _GEN_69; // @[TLB.scala 73:41]
  assign _GEN_76 = _T_85 | _GEN_70; // @[TLB.scala 73:41]
  assign _GEN_78 = _T_78[53] ? _GEN_72 : _GEN_66; // @[TLB.scala 67:26]
  assign _GEN_79 = _T_78[53] ? _GEN_73 : _GEN_67; // @[TLB.scala 67:26]
  assign _GEN_81 = _T_78[53] ? _GEN_75 : _GEN_69; // @[TLB.scala 67:26]
  assign _GEN_82 = _T_78[53] ? _GEN_76 : _GEN_70; // @[TLB.scala 67:26]
  assign _T_90 = tlb__T_88_data;
  assign _T_94 = _T_90[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_84 = _T_94 ? 6'h7 : _GEN_78; // @[TLB.scala 68:41]
  assign _GEN_85 = _T_94 | _GEN_79; // @[TLB.scala 68:41]
  assign _T_97 = _T_90[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_87 = _T_97 ? 6'h7 : _GEN_81; // @[TLB.scala 73:41]
  assign _GEN_88 = _T_97 | _GEN_82; // @[TLB.scala 73:41]
  assign _GEN_90 = _T_90[53] ? _GEN_84 : _GEN_78; // @[TLB.scala 67:26]
  assign _GEN_91 = _T_90[53] ? _GEN_85 : _GEN_79; // @[TLB.scala 67:26]
  assign _GEN_93 = _T_90[53] ? _GEN_87 : _GEN_81; // @[TLB.scala 67:26]
  assign _GEN_94 = _T_90[53] ? _GEN_88 : _GEN_82; // @[TLB.scala 67:26]
  assign _T_102 = tlb__T_100_data;
  assign _T_106 = _T_102[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_96 = _T_106 ? 6'h8 : _GEN_90; // @[TLB.scala 68:41]
  assign _GEN_97 = _T_106 | _GEN_91; // @[TLB.scala 68:41]
  assign _T_109 = _T_102[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_99 = _T_109 ? 6'h8 : _GEN_93; // @[TLB.scala 73:41]
  assign _GEN_100 = _T_109 | _GEN_94; // @[TLB.scala 73:41]
  assign _GEN_102 = _T_102[53] ? _GEN_96 : _GEN_90; // @[TLB.scala 67:26]
  assign _GEN_103 = _T_102[53] ? _GEN_97 : _GEN_91; // @[TLB.scala 67:26]
  assign _GEN_105 = _T_102[53] ? _GEN_99 : _GEN_93; // @[TLB.scala 67:26]
  assign _GEN_106 = _T_102[53] ? _GEN_100 : _GEN_94; // @[TLB.scala 67:26]
  assign _T_114 = tlb__T_112_data;
  assign _T_118 = _T_114[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_108 = _T_118 ? 6'h9 : _GEN_102; // @[TLB.scala 68:41]
  assign _GEN_109 = _T_118 | _GEN_103; // @[TLB.scala 68:41]
  assign _T_121 = _T_114[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_111 = _T_121 ? 6'h9 : _GEN_105; // @[TLB.scala 73:41]
  assign _GEN_112 = _T_121 | _GEN_106; // @[TLB.scala 73:41]
  assign _GEN_114 = _T_114[53] ? _GEN_108 : _GEN_102; // @[TLB.scala 67:26]
  assign _GEN_115 = _T_114[53] ? _GEN_109 : _GEN_103; // @[TLB.scala 67:26]
  assign _GEN_117 = _T_114[53] ? _GEN_111 : _GEN_105; // @[TLB.scala 67:26]
  assign _GEN_118 = _T_114[53] ? _GEN_112 : _GEN_106; // @[TLB.scala 67:26]
  assign _T_126 = tlb__T_124_data;
  assign _T_130 = _T_126[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_120 = _T_130 ? 6'ha : _GEN_114; // @[TLB.scala 68:41]
  assign _GEN_121 = _T_130 | _GEN_115; // @[TLB.scala 68:41]
  assign _T_133 = _T_126[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_123 = _T_133 ? 6'ha : _GEN_117; // @[TLB.scala 73:41]
  assign _GEN_124 = _T_133 | _GEN_118; // @[TLB.scala 73:41]
  assign _GEN_126 = _T_126[53] ? _GEN_120 : _GEN_114; // @[TLB.scala 67:26]
  assign _GEN_127 = _T_126[53] ? _GEN_121 : _GEN_115; // @[TLB.scala 67:26]
  assign _GEN_129 = _T_126[53] ? _GEN_123 : _GEN_117; // @[TLB.scala 67:26]
  assign _GEN_130 = _T_126[53] ? _GEN_124 : _GEN_118; // @[TLB.scala 67:26]
  assign _T_138 = tlb__T_136_data;
  assign _T_142 = _T_138[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_132 = _T_142 ? 6'hb : _GEN_126; // @[TLB.scala 68:41]
  assign _GEN_133 = _T_142 | _GEN_127; // @[TLB.scala 68:41]
  assign _T_145 = _T_138[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_135 = _T_145 ? 6'hb : _GEN_129; // @[TLB.scala 73:41]
  assign _GEN_136 = _T_145 | _GEN_130; // @[TLB.scala 73:41]
  assign _GEN_138 = _T_138[53] ? _GEN_132 : _GEN_126; // @[TLB.scala 67:26]
  assign _GEN_139 = _T_138[53] ? _GEN_133 : _GEN_127; // @[TLB.scala 67:26]
  assign _GEN_141 = _T_138[53] ? _GEN_135 : _GEN_129; // @[TLB.scala 67:26]
  assign _GEN_142 = _T_138[53] ? _GEN_136 : _GEN_130; // @[TLB.scala 67:26]
  assign _T_150 = tlb__T_148_data;
  assign _T_154 = _T_150[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_144 = _T_154 ? 6'hc : _GEN_138; // @[TLB.scala 68:41]
  assign _GEN_145 = _T_154 | _GEN_139; // @[TLB.scala 68:41]
  assign _T_157 = _T_150[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_147 = _T_157 ? 6'hc : _GEN_141; // @[TLB.scala 73:41]
  assign _GEN_148 = _T_157 | _GEN_142; // @[TLB.scala 73:41]
  assign _GEN_150 = _T_150[53] ? _GEN_144 : _GEN_138; // @[TLB.scala 67:26]
  assign _GEN_151 = _T_150[53] ? _GEN_145 : _GEN_139; // @[TLB.scala 67:26]
  assign _GEN_153 = _T_150[53] ? _GEN_147 : _GEN_141; // @[TLB.scala 67:26]
  assign _GEN_154 = _T_150[53] ? _GEN_148 : _GEN_142; // @[TLB.scala 67:26]
  assign _T_162 = tlb__T_160_data;
  assign _T_166 = _T_162[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_156 = _T_166 ? 6'hd : _GEN_150; // @[TLB.scala 68:41]
  assign _GEN_157 = _T_166 | _GEN_151; // @[TLB.scala 68:41]
  assign _T_169 = _T_162[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_159 = _T_169 ? 6'hd : _GEN_153; // @[TLB.scala 73:41]
  assign _GEN_160 = _T_169 | _GEN_154; // @[TLB.scala 73:41]
  assign _GEN_162 = _T_162[53] ? _GEN_156 : _GEN_150; // @[TLB.scala 67:26]
  assign _GEN_163 = _T_162[53] ? _GEN_157 : _GEN_151; // @[TLB.scala 67:26]
  assign _GEN_165 = _T_162[53] ? _GEN_159 : _GEN_153; // @[TLB.scala 67:26]
  assign _GEN_166 = _T_162[53] ? _GEN_160 : _GEN_154; // @[TLB.scala 67:26]
  assign _T_174 = tlb__T_172_data;
  assign _T_178 = _T_174[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_168 = _T_178 ? 6'he : _GEN_162; // @[TLB.scala 68:41]
  assign _GEN_169 = _T_178 | _GEN_163; // @[TLB.scala 68:41]
  assign _T_181 = _T_174[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_171 = _T_181 ? 6'he : _GEN_165; // @[TLB.scala 73:41]
  assign _GEN_172 = _T_181 | _GEN_166; // @[TLB.scala 73:41]
  assign _GEN_174 = _T_174[53] ? _GEN_168 : _GEN_162; // @[TLB.scala 67:26]
  assign _GEN_175 = _T_174[53] ? _GEN_169 : _GEN_163; // @[TLB.scala 67:26]
  assign _GEN_177 = _T_174[53] ? _GEN_171 : _GEN_165; // @[TLB.scala 67:26]
  assign _GEN_178 = _T_174[53] ? _GEN_172 : _GEN_166; // @[TLB.scala 67:26]
  assign _T_186 = tlb__T_184_data;
  assign _T_190 = _T_186[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_180 = _T_190 ? 6'hf : _GEN_174; // @[TLB.scala 68:41]
  assign _GEN_181 = _T_190 | _GEN_175; // @[TLB.scala 68:41]
  assign _T_193 = _T_186[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_183 = _T_193 ? 6'hf : _GEN_177; // @[TLB.scala 73:41]
  assign _GEN_184 = _T_193 | _GEN_178; // @[TLB.scala 73:41]
  assign _GEN_186 = _T_186[53] ? _GEN_180 : _GEN_174; // @[TLB.scala 67:26]
  assign _GEN_187 = _T_186[53] ? _GEN_181 : _GEN_175; // @[TLB.scala 67:26]
  assign _GEN_189 = _T_186[53] ? _GEN_183 : _GEN_177; // @[TLB.scala 67:26]
  assign _GEN_190 = _T_186[53] ? _GEN_184 : _GEN_178; // @[TLB.scala 67:26]
  assign _T_198 = tlb__T_196_data;
  assign _T_202 = _T_198[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_192 = _T_202 ? 6'h10 : _GEN_186; // @[TLB.scala 68:41]
  assign _GEN_193 = _T_202 | _GEN_187; // @[TLB.scala 68:41]
  assign _T_205 = _T_198[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_195 = _T_205 ? 6'h10 : _GEN_189; // @[TLB.scala 73:41]
  assign _GEN_196 = _T_205 | _GEN_190; // @[TLB.scala 73:41]
  assign _GEN_198 = _T_198[53] ? _GEN_192 : _GEN_186; // @[TLB.scala 67:26]
  assign _GEN_199 = _T_198[53] ? _GEN_193 : _GEN_187; // @[TLB.scala 67:26]
  assign _GEN_201 = _T_198[53] ? _GEN_195 : _GEN_189; // @[TLB.scala 67:26]
  assign _GEN_202 = _T_198[53] ? _GEN_196 : _GEN_190; // @[TLB.scala 67:26]
  assign _T_210 = tlb__T_208_data;
  assign _T_214 = _T_210[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_204 = _T_214 ? 6'h11 : _GEN_198; // @[TLB.scala 68:41]
  assign _GEN_205 = _T_214 | _GEN_199; // @[TLB.scala 68:41]
  assign _T_217 = _T_210[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_207 = _T_217 ? 6'h11 : _GEN_201; // @[TLB.scala 73:41]
  assign _GEN_208 = _T_217 | _GEN_202; // @[TLB.scala 73:41]
  assign _GEN_210 = _T_210[53] ? _GEN_204 : _GEN_198; // @[TLB.scala 67:26]
  assign _GEN_211 = _T_210[53] ? _GEN_205 : _GEN_199; // @[TLB.scala 67:26]
  assign _GEN_213 = _T_210[53] ? _GEN_207 : _GEN_201; // @[TLB.scala 67:26]
  assign _GEN_214 = _T_210[53] ? _GEN_208 : _GEN_202; // @[TLB.scala 67:26]
  assign _T_222 = tlb__T_220_data;
  assign _T_226 = _T_222[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_216 = _T_226 ? 6'h12 : _GEN_210; // @[TLB.scala 68:41]
  assign _GEN_217 = _T_226 | _GEN_211; // @[TLB.scala 68:41]
  assign _T_229 = _T_222[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_219 = _T_229 ? 6'h12 : _GEN_213; // @[TLB.scala 73:41]
  assign _GEN_220 = _T_229 | _GEN_214; // @[TLB.scala 73:41]
  assign _GEN_222 = _T_222[53] ? _GEN_216 : _GEN_210; // @[TLB.scala 67:26]
  assign _GEN_223 = _T_222[53] ? _GEN_217 : _GEN_211; // @[TLB.scala 67:26]
  assign _GEN_225 = _T_222[53] ? _GEN_219 : _GEN_213; // @[TLB.scala 67:26]
  assign _GEN_226 = _T_222[53] ? _GEN_220 : _GEN_214; // @[TLB.scala 67:26]
  assign _T_234 = tlb__T_232_data;
  assign _T_238 = _T_234[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_228 = _T_238 ? 6'h13 : _GEN_222; // @[TLB.scala 68:41]
  assign _GEN_229 = _T_238 | _GEN_223; // @[TLB.scala 68:41]
  assign _T_241 = _T_234[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_231 = _T_241 ? 6'h13 : _GEN_225; // @[TLB.scala 73:41]
  assign _GEN_232 = _T_241 | _GEN_226; // @[TLB.scala 73:41]
  assign _GEN_234 = _T_234[53] ? _GEN_228 : _GEN_222; // @[TLB.scala 67:26]
  assign _GEN_235 = _T_234[53] ? _GEN_229 : _GEN_223; // @[TLB.scala 67:26]
  assign _GEN_237 = _T_234[53] ? _GEN_231 : _GEN_225; // @[TLB.scala 67:26]
  assign _GEN_238 = _T_234[53] ? _GEN_232 : _GEN_226; // @[TLB.scala 67:26]
  assign _T_246 = tlb__T_244_data;
  assign _T_250 = _T_246[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_240 = _T_250 ? 6'h14 : _GEN_234; // @[TLB.scala 68:41]
  assign _GEN_241 = _T_250 | _GEN_235; // @[TLB.scala 68:41]
  assign _T_253 = _T_246[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_243 = _T_253 ? 6'h14 : _GEN_237; // @[TLB.scala 73:41]
  assign _GEN_244 = _T_253 | _GEN_238; // @[TLB.scala 73:41]
  assign _GEN_246 = _T_246[53] ? _GEN_240 : _GEN_234; // @[TLB.scala 67:26]
  assign _GEN_247 = _T_246[53] ? _GEN_241 : _GEN_235; // @[TLB.scala 67:26]
  assign _GEN_249 = _T_246[53] ? _GEN_243 : _GEN_237; // @[TLB.scala 67:26]
  assign _GEN_250 = _T_246[53] ? _GEN_244 : _GEN_238; // @[TLB.scala 67:26]
  assign _T_258 = tlb__T_256_data;
  assign _T_262 = _T_258[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_252 = _T_262 ? 6'h15 : _GEN_246; // @[TLB.scala 68:41]
  assign _GEN_253 = _T_262 | _GEN_247; // @[TLB.scala 68:41]
  assign _T_265 = _T_258[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_255 = _T_265 ? 6'h15 : _GEN_249; // @[TLB.scala 73:41]
  assign _GEN_256 = _T_265 | _GEN_250; // @[TLB.scala 73:41]
  assign _GEN_258 = _T_258[53] ? _GEN_252 : _GEN_246; // @[TLB.scala 67:26]
  assign _GEN_259 = _T_258[53] ? _GEN_253 : _GEN_247; // @[TLB.scala 67:26]
  assign _GEN_261 = _T_258[53] ? _GEN_255 : _GEN_249; // @[TLB.scala 67:26]
  assign _GEN_262 = _T_258[53] ? _GEN_256 : _GEN_250; // @[TLB.scala 67:26]
  assign _T_270 = tlb__T_268_data;
  assign _T_274 = _T_270[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_264 = _T_274 ? 6'h16 : _GEN_258; // @[TLB.scala 68:41]
  assign _GEN_265 = _T_274 | _GEN_259; // @[TLB.scala 68:41]
  assign _T_277 = _T_270[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_267 = _T_277 ? 6'h16 : _GEN_261; // @[TLB.scala 73:41]
  assign _GEN_268 = _T_277 | _GEN_262; // @[TLB.scala 73:41]
  assign _GEN_270 = _T_270[53] ? _GEN_264 : _GEN_258; // @[TLB.scala 67:26]
  assign _GEN_271 = _T_270[53] ? _GEN_265 : _GEN_259; // @[TLB.scala 67:26]
  assign _GEN_273 = _T_270[53] ? _GEN_267 : _GEN_261; // @[TLB.scala 67:26]
  assign _GEN_274 = _T_270[53] ? _GEN_268 : _GEN_262; // @[TLB.scala 67:26]
  assign _T_282 = tlb__T_280_data;
  assign _T_286 = _T_282[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_276 = _T_286 ? 6'h17 : _GEN_270; // @[TLB.scala 68:41]
  assign _GEN_277 = _T_286 | _GEN_271; // @[TLB.scala 68:41]
  assign _T_289 = _T_282[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_279 = _T_289 ? 6'h17 : _GEN_273; // @[TLB.scala 73:41]
  assign _GEN_280 = _T_289 | _GEN_274; // @[TLB.scala 73:41]
  assign _GEN_282 = _T_282[53] ? _GEN_276 : _GEN_270; // @[TLB.scala 67:26]
  assign _GEN_283 = _T_282[53] ? _GEN_277 : _GEN_271; // @[TLB.scala 67:26]
  assign _GEN_285 = _T_282[53] ? _GEN_279 : _GEN_273; // @[TLB.scala 67:26]
  assign _GEN_286 = _T_282[53] ? _GEN_280 : _GEN_274; // @[TLB.scala 67:26]
  assign _T_294 = tlb__T_292_data;
  assign _T_298 = _T_294[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_288 = _T_298 ? 6'h18 : _GEN_282; // @[TLB.scala 68:41]
  assign _GEN_289 = _T_298 | _GEN_283; // @[TLB.scala 68:41]
  assign _T_301 = _T_294[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_291 = _T_301 ? 6'h18 : _GEN_285; // @[TLB.scala 73:41]
  assign _GEN_292 = _T_301 | _GEN_286; // @[TLB.scala 73:41]
  assign _GEN_294 = _T_294[53] ? _GEN_288 : _GEN_282; // @[TLB.scala 67:26]
  assign _GEN_295 = _T_294[53] ? _GEN_289 : _GEN_283; // @[TLB.scala 67:26]
  assign _GEN_297 = _T_294[53] ? _GEN_291 : _GEN_285; // @[TLB.scala 67:26]
  assign _GEN_298 = _T_294[53] ? _GEN_292 : _GEN_286; // @[TLB.scala 67:26]
  assign _T_306 = tlb__T_304_data;
  assign _T_310 = _T_306[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_300 = _T_310 ? 6'h19 : _GEN_294; // @[TLB.scala 68:41]
  assign _GEN_301 = _T_310 | _GEN_295; // @[TLB.scala 68:41]
  assign _T_313 = _T_306[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_303 = _T_313 ? 6'h19 : _GEN_297; // @[TLB.scala 73:41]
  assign _GEN_304 = _T_313 | _GEN_298; // @[TLB.scala 73:41]
  assign _GEN_306 = _T_306[53] ? _GEN_300 : _GEN_294; // @[TLB.scala 67:26]
  assign _GEN_307 = _T_306[53] ? _GEN_301 : _GEN_295; // @[TLB.scala 67:26]
  assign _GEN_309 = _T_306[53] ? _GEN_303 : _GEN_297; // @[TLB.scala 67:26]
  assign _GEN_310 = _T_306[53] ? _GEN_304 : _GEN_298; // @[TLB.scala 67:26]
  assign _T_318 = tlb__T_316_data;
  assign _T_322 = _T_318[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_312 = _T_322 ? 6'h1a : _GEN_306; // @[TLB.scala 68:41]
  assign _GEN_313 = _T_322 | _GEN_307; // @[TLB.scala 68:41]
  assign _T_325 = _T_318[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_315 = _T_325 ? 6'h1a : _GEN_309; // @[TLB.scala 73:41]
  assign _GEN_316 = _T_325 | _GEN_310; // @[TLB.scala 73:41]
  assign _GEN_318 = _T_318[53] ? _GEN_312 : _GEN_306; // @[TLB.scala 67:26]
  assign _GEN_319 = _T_318[53] ? _GEN_313 : _GEN_307; // @[TLB.scala 67:26]
  assign _GEN_321 = _T_318[53] ? _GEN_315 : _GEN_309; // @[TLB.scala 67:26]
  assign _GEN_322 = _T_318[53] ? _GEN_316 : _GEN_310; // @[TLB.scala 67:26]
  assign _T_330 = tlb__T_328_data;
  assign _T_334 = _T_330[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_324 = _T_334 ? 6'h1b : _GEN_318; // @[TLB.scala 68:41]
  assign _GEN_325 = _T_334 | _GEN_319; // @[TLB.scala 68:41]
  assign _T_337 = _T_330[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_327 = _T_337 ? 6'h1b : _GEN_321; // @[TLB.scala 73:41]
  assign _GEN_328 = _T_337 | _GEN_322; // @[TLB.scala 73:41]
  assign _GEN_330 = _T_330[53] ? _GEN_324 : _GEN_318; // @[TLB.scala 67:26]
  assign _GEN_331 = _T_330[53] ? _GEN_325 : _GEN_319; // @[TLB.scala 67:26]
  assign _GEN_333 = _T_330[53] ? _GEN_327 : _GEN_321; // @[TLB.scala 67:26]
  assign _GEN_334 = _T_330[53] ? _GEN_328 : _GEN_322; // @[TLB.scala 67:26]
  assign _T_342 = tlb__T_340_data;
  assign _T_346 = _T_342[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_336 = _T_346 ? 6'h1c : _GEN_330; // @[TLB.scala 68:41]
  assign _GEN_337 = _T_346 | _GEN_331; // @[TLB.scala 68:41]
  assign _T_349 = _T_342[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_339 = _T_349 ? 6'h1c : _GEN_333; // @[TLB.scala 73:41]
  assign _GEN_340 = _T_349 | _GEN_334; // @[TLB.scala 73:41]
  assign _GEN_342 = _T_342[53] ? _GEN_336 : _GEN_330; // @[TLB.scala 67:26]
  assign _GEN_343 = _T_342[53] ? _GEN_337 : _GEN_331; // @[TLB.scala 67:26]
  assign _GEN_345 = _T_342[53] ? _GEN_339 : _GEN_333; // @[TLB.scala 67:26]
  assign _GEN_346 = _T_342[53] ? _GEN_340 : _GEN_334; // @[TLB.scala 67:26]
  assign _T_354 = tlb__T_352_data;
  assign _T_358 = _T_354[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_348 = _T_358 ? 6'h1d : _GEN_342; // @[TLB.scala 68:41]
  assign _GEN_349 = _T_358 | _GEN_343; // @[TLB.scala 68:41]
  assign _T_361 = _T_354[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_351 = _T_361 ? 6'h1d : _GEN_345; // @[TLB.scala 73:41]
  assign _GEN_352 = _T_361 | _GEN_346; // @[TLB.scala 73:41]
  assign _GEN_354 = _T_354[53] ? _GEN_348 : _GEN_342; // @[TLB.scala 67:26]
  assign _GEN_355 = _T_354[53] ? _GEN_349 : _GEN_343; // @[TLB.scala 67:26]
  assign _GEN_357 = _T_354[53] ? _GEN_351 : _GEN_345; // @[TLB.scala 67:26]
  assign _GEN_358 = _T_354[53] ? _GEN_352 : _GEN_346; // @[TLB.scala 67:26]
  assign _T_366 = tlb__T_364_data;
  assign _T_370 = _T_366[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_360 = _T_370 ? 6'h1e : _GEN_354; // @[TLB.scala 68:41]
  assign _GEN_361 = _T_370 | _GEN_355; // @[TLB.scala 68:41]
  assign _T_373 = _T_366[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_363 = _T_373 ? 6'h1e : _GEN_357; // @[TLB.scala 73:41]
  assign _GEN_364 = _T_373 | _GEN_358; // @[TLB.scala 73:41]
  assign _GEN_366 = _T_366[53] ? _GEN_360 : _GEN_354; // @[TLB.scala 67:26]
  assign _GEN_367 = _T_366[53] ? _GEN_361 : _GEN_355; // @[TLB.scala 67:26]
  assign _GEN_369 = _T_366[53] ? _GEN_363 : _GEN_357; // @[TLB.scala 67:26]
  assign _GEN_370 = _T_366[53] ? _GEN_364 : _GEN_358; // @[TLB.scala 67:26]
  assign _T_378 = tlb__T_376_data;
  assign _T_382 = _T_378[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_372 = _T_382 ? 6'h1f : _GEN_366; // @[TLB.scala 68:41]
  assign _GEN_373 = _T_382 | _GEN_367; // @[TLB.scala 68:41]
  assign _T_385 = _T_378[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_375 = _T_385 ? 6'h1f : _GEN_369; // @[TLB.scala 73:41]
  assign _GEN_376 = _T_385 | _GEN_370; // @[TLB.scala 73:41]
  assign _GEN_378 = _T_378[53] ? _GEN_372 : _GEN_366; // @[TLB.scala 67:26]
  assign _GEN_379 = _T_378[53] ? _GEN_373 : _GEN_367; // @[TLB.scala 67:26]
  assign _GEN_381 = _T_378[53] ? _GEN_375 : _GEN_369; // @[TLB.scala 67:26]
  assign _GEN_382 = _T_378[53] ? _GEN_376 : _GEN_370; // @[TLB.scala 67:26]
  assign _T_390 = tlb__T_388_data;
  assign _T_394 = _T_390[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_384 = _T_394 ? 6'h20 : _GEN_378; // @[TLB.scala 68:41]
  assign _GEN_385 = _T_394 | _GEN_379; // @[TLB.scala 68:41]
  assign _T_397 = _T_390[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_387 = _T_397 ? 6'h20 : _GEN_381; // @[TLB.scala 73:41]
  assign _GEN_388 = _T_397 | _GEN_382; // @[TLB.scala 73:41]
  assign _GEN_390 = _T_390[53] ? _GEN_384 : _GEN_378; // @[TLB.scala 67:26]
  assign _GEN_391 = _T_390[53] ? _GEN_385 : _GEN_379; // @[TLB.scala 67:26]
  assign _GEN_393 = _T_390[53] ? _GEN_387 : _GEN_381; // @[TLB.scala 67:26]
  assign _GEN_394 = _T_390[53] ? _GEN_388 : _GEN_382; // @[TLB.scala 67:26]
  assign _T_402 = tlb__T_400_data;
  assign _T_406 = _T_402[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_396 = _T_406 ? 6'h21 : _GEN_390; // @[TLB.scala 68:41]
  assign _GEN_397 = _T_406 | _GEN_391; // @[TLB.scala 68:41]
  assign _T_409 = _T_402[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_399 = _T_409 ? 6'h21 : _GEN_393; // @[TLB.scala 73:41]
  assign _GEN_400 = _T_409 | _GEN_394; // @[TLB.scala 73:41]
  assign _GEN_402 = _T_402[53] ? _GEN_396 : _GEN_390; // @[TLB.scala 67:26]
  assign _GEN_403 = _T_402[53] ? _GEN_397 : _GEN_391; // @[TLB.scala 67:26]
  assign _GEN_405 = _T_402[53] ? _GEN_399 : _GEN_393; // @[TLB.scala 67:26]
  assign _GEN_406 = _T_402[53] ? _GEN_400 : _GEN_394; // @[TLB.scala 67:26]
  assign _T_414 = tlb__T_412_data;
  assign _T_418 = _T_414[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_408 = _T_418 ? 6'h22 : _GEN_402; // @[TLB.scala 68:41]
  assign _GEN_409 = _T_418 | _GEN_403; // @[TLB.scala 68:41]
  assign _T_421 = _T_414[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_411 = _T_421 ? 6'h22 : _GEN_405; // @[TLB.scala 73:41]
  assign _GEN_412 = _T_421 | _GEN_406; // @[TLB.scala 73:41]
  assign _GEN_414 = _T_414[53] ? _GEN_408 : _GEN_402; // @[TLB.scala 67:26]
  assign _GEN_415 = _T_414[53] ? _GEN_409 : _GEN_403; // @[TLB.scala 67:26]
  assign _GEN_417 = _T_414[53] ? _GEN_411 : _GEN_405; // @[TLB.scala 67:26]
  assign _GEN_418 = _T_414[53] ? _GEN_412 : _GEN_406; // @[TLB.scala 67:26]
  assign _T_426 = tlb__T_424_data;
  assign _T_430 = _T_426[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_420 = _T_430 ? 6'h23 : _GEN_414; // @[TLB.scala 68:41]
  assign _GEN_421 = _T_430 | _GEN_415; // @[TLB.scala 68:41]
  assign _T_433 = _T_426[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_423 = _T_433 ? 6'h23 : _GEN_417; // @[TLB.scala 73:41]
  assign _GEN_424 = _T_433 | _GEN_418; // @[TLB.scala 73:41]
  assign _GEN_426 = _T_426[53] ? _GEN_420 : _GEN_414; // @[TLB.scala 67:26]
  assign _GEN_427 = _T_426[53] ? _GEN_421 : _GEN_415; // @[TLB.scala 67:26]
  assign _GEN_429 = _T_426[53] ? _GEN_423 : _GEN_417; // @[TLB.scala 67:26]
  assign _GEN_430 = _T_426[53] ? _GEN_424 : _GEN_418; // @[TLB.scala 67:26]
  assign _T_438 = tlb__T_436_data;
  assign _T_442 = _T_438[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_432 = _T_442 ? 6'h24 : _GEN_426; // @[TLB.scala 68:41]
  assign _GEN_433 = _T_442 | _GEN_427; // @[TLB.scala 68:41]
  assign _T_445 = _T_438[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_435 = _T_445 ? 6'h24 : _GEN_429; // @[TLB.scala 73:41]
  assign _GEN_436 = _T_445 | _GEN_430; // @[TLB.scala 73:41]
  assign _GEN_438 = _T_438[53] ? _GEN_432 : _GEN_426; // @[TLB.scala 67:26]
  assign _GEN_439 = _T_438[53] ? _GEN_433 : _GEN_427; // @[TLB.scala 67:26]
  assign _GEN_441 = _T_438[53] ? _GEN_435 : _GEN_429; // @[TLB.scala 67:26]
  assign _GEN_442 = _T_438[53] ? _GEN_436 : _GEN_430; // @[TLB.scala 67:26]
  assign _T_450 = tlb__T_448_data;
  assign _T_454 = _T_450[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_444 = _T_454 ? 6'h25 : _GEN_438; // @[TLB.scala 68:41]
  assign _GEN_445 = _T_454 | _GEN_439; // @[TLB.scala 68:41]
  assign _T_457 = _T_450[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_447 = _T_457 ? 6'h25 : _GEN_441; // @[TLB.scala 73:41]
  assign _GEN_448 = _T_457 | _GEN_442; // @[TLB.scala 73:41]
  assign _GEN_450 = _T_450[53] ? _GEN_444 : _GEN_438; // @[TLB.scala 67:26]
  assign _GEN_451 = _T_450[53] ? _GEN_445 : _GEN_439; // @[TLB.scala 67:26]
  assign _GEN_453 = _T_450[53] ? _GEN_447 : _GEN_441; // @[TLB.scala 67:26]
  assign _GEN_454 = _T_450[53] ? _GEN_448 : _GEN_442; // @[TLB.scala 67:26]
  assign _T_462 = tlb__T_460_data;
  assign _T_466 = _T_462[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_456 = _T_466 ? 6'h26 : _GEN_450; // @[TLB.scala 68:41]
  assign _GEN_457 = _T_466 | _GEN_451; // @[TLB.scala 68:41]
  assign _T_469 = _T_462[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_459 = _T_469 ? 6'h26 : _GEN_453; // @[TLB.scala 73:41]
  assign _GEN_460 = _T_469 | _GEN_454; // @[TLB.scala 73:41]
  assign _GEN_462 = _T_462[53] ? _GEN_456 : _GEN_450; // @[TLB.scala 67:26]
  assign _GEN_463 = _T_462[53] ? _GEN_457 : _GEN_451; // @[TLB.scala 67:26]
  assign _GEN_465 = _T_462[53] ? _GEN_459 : _GEN_453; // @[TLB.scala 67:26]
  assign _GEN_466 = _T_462[53] ? _GEN_460 : _GEN_454; // @[TLB.scala 67:26]
  assign _T_474 = tlb__T_472_data;
  assign _T_478 = _T_474[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_468 = _T_478 ? 6'h27 : _GEN_462; // @[TLB.scala 68:41]
  assign _GEN_469 = _T_478 | _GEN_463; // @[TLB.scala 68:41]
  assign _T_481 = _T_474[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_471 = _T_481 ? 6'h27 : _GEN_465; // @[TLB.scala 73:41]
  assign _GEN_472 = _T_481 | _GEN_466; // @[TLB.scala 73:41]
  assign _GEN_474 = _T_474[53] ? _GEN_468 : _GEN_462; // @[TLB.scala 67:26]
  assign _GEN_475 = _T_474[53] ? _GEN_469 : _GEN_463; // @[TLB.scala 67:26]
  assign _GEN_477 = _T_474[53] ? _GEN_471 : _GEN_465; // @[TLB.scala 67:26]
  assign _GEN_478 = _T_474[53] ? _GEN_472 : _GEN_466; // @[TLB.scala 67:26]
  assign _T_486 = tlb__T_484_data;
  assign _T_490 = _T_486[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_480 = _T_490 ? 6'h28 : _GEN_474; // @[TLB.scala 68:41]
  assign _GEN_481 = _T_490 | _GEN_475; // @[TLB.scala 68:41]
  assign _T_493 = _T_486[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_483 = _T_493 ? 6'h28 : _GEN_477; // @[TLB.scala 73:41]
  assign _GEN_484 = _T_493 | _GEN_478; // @[TLB.scala 73:41]
  assign _GEN_486 = _T_486[53] ? _GEN_480 : _GEN_474; // @[TLB.scala 67:26]
  assign _GEN_487 = _T_486[53] ? _GEN_481 : _GEN_475; // @[TLB.scala 67:26]
  assign _GEN_489 = _T_486[53] ? _GEN_483 : _GEN_477; // @[TLB.scala 67:26]
  assign _GEN_490 = _T_486[53] ? _GEN_484 : _GEN_478; // @[TLB.scala 67:26]
  assign _T_498 = tlb__T_496_data;
  assign _T_502 = _T_498[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_492 = _T_502 ? 6'h29 : _GEN_486; // @[TLB.scala 68:41]
  assign _GEN_493 = _T_502 | _GEN_487; // @[TLB.scala 68:41]
  assign _T_505 = _T_498[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_495 = _T_505 ? 6'h29 : _GEN_489; // @[TLB.scala 73:41]
  assign _GEN_496 = _T_505 | _GEN_490; // @[TLB.scala 73:41]
  assign _GEN_498 = _T_498[53] ? _GEN_492 : _GEN_486; // @[TLB.scala 67:26]
  assign _GEN_499 = _T_498[53] ? _GEN_493 : _GEN_487; // @[TLB.scala 67:26]
  assign _GEN_501 = _T_498[53] ? _GEN_495 : _GEN_489; // @[TLB.scala 67:26]
  assign _GEN_502 = _T_498[53] ? _GEN_496 : _GEN_490; // @[TLB.scala 67:26]
  assign _T_510 = tlb__T_508_data;
  assign _T_514 = _T_510[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_504 = _T_514 ? 6'h2a : _GEN_498; // @[TLB.scala 68:41]
  assign _GEN_505 = _T_514 | _GEN_499; // @[TLB.scala 68:41]
  assign _T_517 = _T_510[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_507 = _T_517 ? 6'h2a : _GEN_501; // @[TLB.scala 73:41]
  assign _GEN_508 = _T_517 | _GEN_502; // @[TLB.scala 73:41]
  assign _GEN_510 = _T_510[53] ? _GEN_504 : _GEN_498; // @[TLB.scala 67:26]
  assign _GEN_511 = _T_510[53] ? _GEN_505 : _GEN_499; // @[TLB.scala 67:26]
  assign _GEN_513 = _T_510[53] ? _GEN_507 : _GEN_501; // @[TLB.scala 67:26]
  assign _GEN_514 = _T_510[53] ? _GEN_508 : _GEN_502; // @[TLB.scala 67:26]
  assign _T_522 = tlb__T_520_data;
  assign _T_526 = _T_522[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_516 = _T_526 ? 6'h2b : _GEN_510; // @[TLB.scala 68:41]
  assign _GEN_517 = _T_526 | _GEN_511; // @[TLB.scala 68:41]
  assign _T_529 = _T_522[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_519 = _T_529 ? 6'h2b : _GEN_513; // @[TLB.scala 73:41]
  assign _GEN_520 = _T_529 | _GEN_514; // @[TLB.scala 73:41]
  assign _GEN_522 = _T_522[53] ? _GEN_516 : _GEN_510; // @[TLB.scala 67:26]
  assign _GEN_523 = _T_522[53] ? _GEN_517 : _GEN_511; // @[TLB.scala 67:26]
  assign _GEN_525 = _T_522[53] ? _GEN_519 : _GEN_513; // @[TLB.scala 67:26]
  assign _GEN_526 = _T_522[53] ? _GEN_520 : _GEN_514; // @[TLB.scala 67:26]
  assign _T_534 = tlb__T_532_data;
  assign _T_538 = _T_534[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_528 = _T_538 ? 6'h2c : _GEN_522; // @[TLB.scala 68:41]
  assign _GEN_529 = _T_538 | _GEN_523; // @[TLB.scala 68:41]
  assign _T_541 = _T_534[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_531 = _T_541 ? 6'h2c : _GEN_525; // @[TLB.scala 73:41]
  assign _GEN_532 = _T_541 | _GEN_526; // @[TLB.scala 73:41]
  assign _GEN_534 = _T_534[53] ? _GEN_528 : _GEN_522; // @[TLB.scala 67:26]
  assign _GEN_535 = _T_534[53] ? _GEN_529 : _GEN_523; // @[TLB.scala 67:26]
  assign _GEN_537 = _T_534[53] ? _GEN_531 : _GEN_525; // @[TLB.scala 67:26]
  assign _GEN_538 = _T_534[53] ? _GEN_532 : _GEN_526; // @[TLB.scala 67:26]
  assign _T_546 = tlb__T_544_data;
  assign _T_550 = _T_546[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_540 = _T_550 ? 6'h2d : _GEN_534; // @[TLB.scala 68:41]
  assign _GEN_541 = _T_550 | _GEN_535; // @[TLB.scala 68:41]
  assign _T_553 = _T_546[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_543 = _T_553 ? 6'h2d : _GEN_537; // @[TLB.scala 73:41]
  assign _GEN_544 = _T_553 | _GEN_538; // @[TLB.scala 73:41]
  assign _GEN_546 = _T_546[53] ? _GEN_540 : _GEN_534; // @[TLB.scala 67:26]
  assign _GEN_547 = _T_546[53] ? _GEN_541 : _GEN_535; // @[TLB.scala 67:26]
  assign _GEN_549 = _T_546[53] ? _GEN_543 : _GEN_537; // @[TLB.scala 67:26]
  assign _GEN_550 = _T_546[53] ? _GEN_544 : _GEN_538; // @[TLB.scala 67:26]
  assign _T_558 = tlb__T_556_data;
  assign _T_562 = _T_558[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_552 = _T_562 ? 6'h2e : _GEN_546; // @[TLB.scala 68:41]
  assign _GEN_553 = _T_562 | _GEN_547; // @[TLB.scala 68:41]
  assign _T_565 = _T_558[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_555 = _T_565 ? 6'h2e : _GEN_549; // @[TLB.scala 73:41]
  assign _GEN_556 = _T_565 | _GEN_550; // @[TLB.scala 73:41]
  assign _GEN_558 = _T_558[53] ? _GEN_552 : _GEN_546; // @[TLB.scala 67:26]
  assign _GEN_559 = _T_558[53] ? _GEN_553 : _GEN_547; // @[TLB.scala 67:26]
  assign _GEN_561 = _T_558[53] ? _GEN_555 : _GEN_549; // @[TLB.scala 67:26]
  assign _GEN_562 = _T_558[53] ? _GEN_556 : _GEN_550; // @[TLB.scala 67:26]
  assign _T_570 = tlb__T_568_data;
  assign _T_574 = _T_570[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_564 = _T_574 ? 6'h2f : _GEN_558; // @[TLB.scala 68:41]
  assign _GEN_565 = _T_574 | _GEN_559; // @[TLB.scala 68:41]
  assign _T_577 = _T_570[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_567 = _T_577 ? 6'h2f : _GEN_561; // @[TLB.scala 73:41]
  assign _GEN_568 = _T_577 | _GEN_562; // @[TLB.scala 73:41]
  assign _GEN_570 = _T_570[53] ? _GEN_564 : _GEN_558; // @[TLB.scala 67:26]
  assign _GEN_571 = _T_570[53] ? _GEN_565 : _GEN_559; // @[TLB.scala 67:26]
  assign _GEN_573 = _T_570[53] ? _GEN_567 : _GEN_561; // @[TLB.scala 67:26]
  assign _GEN_574 = _T_570[53] ? _GEN_568 : _GEN_562; // @[TLB.scala 67:26]
  assign _T_582 = tlb__T_580_data;
  assign _T_586 = _T_582[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_576 = _T_586 ? 6'h30 : _GEN_570; // @[TLB.scala 68:41]
  assign _GEN_577 = _T_586 | _GEN_571; // @[TLB.scala 68:41]
  assign _T_589 = _T_582[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_579 = _T_589 ? 6'h30 : _GEN_573; // @[TLB.scala 73:41]
  assign _GEN_580 = _T_589 | _GEN_574; // @[TLB.scala 73:41]
  assign _GEN_582 = _T_582[53] ? _GEN_576 : _GEN_570; // @[TLB.scala 67:26]
  assign _GEN_583 = _T_582[53] ? _GEN_577 : _GEN_571; // @[TLB.scala 67:26]
  assign _GEN_585 = _T_582[53] ? _GEN_579 : _GEN_573; // @[TLB.scala 67:26]
  assign _GEN_586 = _T_582[53] ? _GEN_580 : _GEN_574; // @[TLB.scala 67:26]
  assign _T_594 = tlb__T_592_data;
  assign _T_598 = _T_594[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_588 = _T_598 ? 6'h31 : _GEN_582; // @[TLB.scala 68:41]
  assign _GEN_589 = _T_598 | _GEN_583; // @[TLB.scala 68:41]
  assign _T_601 = _T_594[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_591 = _T_601 ? 6'h31 : _GEN_585; // @[TLB.scala 73:41]
  assign _GEN_592 = _T_601 | _GEN_586; // @[TLB.scala 73:41]
  assign _GEN_594 = _T_594[53] ? _GEN_588 : _GEN_582; // @[TLB.scala 67:26]
  assign _GEN_595 = _T_594[53] ? _GEN_589 : _GEN_583; // @[TLB.scala 67:26]
  assign _GEN_597 = _T_594[53] ? _GEN_591 : _GEN_585; // @[TLB.scala 67:26]
  assign _GEN_598 = _T_594[53] ? _GEN_592 : _GEN_586; // @[TLB.scala 67:26]
  assign _T_606 = tlb__T_604_data;
  assign _T_610 = _T_606[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_600 = _T_610 ? 6'h32 : _GEN_594; // @[TLB.scala 68:41]
  assign _GEN_601 = _T_610 | _GEN_595; // @[TLB.scala 68:41]
  assign _T_613 = _T_606[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_603 = _T_613 ? 6'h32 : _GEN_597; // @[TLB.scala 73:41]
  assign _GEN_604 = _T_613 | _GEN_598; // @[TLB.scala 73:41]
  assign _GEN_606 = _T_606[53] ? _GEN_600 : _GEN_594; // @[TLB.scala 67:26]
  assign _GEN_607 = _T_606[53] ? _GEN_601 : _GEN_595; // @[TLB.scala 67:26]
  assign _GEN_609 = _T_606[53] ? _GEN_603 : _GEN_597; // @[TLB.scala 67:26]
  assign _GEN_610 = _T_606[53] ? _GEN_604 : _GEN_598; // @[TLB.scala 67:26]
  assign _T_618 = tlb__T_616_data;
  assign _T_622 = _T_618[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_612 = _T_622 ? 6'h33 : _GEN_606; // @[TLB.scala 68:41]
  assign _GEN_613 = _T_622 | _GEN_607; // @[TLB.scala 68:41]
  assign _T_625 = _T_618[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_615 = _T_625 ? 6'h33 : _GEN_609; // @[TLB.scala 73:41]
  assign _GEN_616 = _T_625 | _GEN_610; // @[TLB.scala 73:41]
  assign _GEN_618 = _T_618[53] ? _GEN_612 : _GEN_606; // @[TLB.scala 67:26]
  assign _GEN_619 = _T_618[53] ? _GEN_613 : _GEN_607; // @[TLB.scala 67:26]
  assign _GEN_621 = _T_618[53] ? _GEN_615 : _GEN_609; // @[TLB.scala 67:26]
  assign _GEN_622 = _T_618[53] ? _GEN_616 : _GEN_610; // @[TLB.scala 67:26]
  assign _T_630 = tlb__T_628_data;
  assign _T_634 = _T_630[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_624 = _T_634 ? 6'h34 : _GEN_618; // @[TLB.scala 68:41]
  assign _GEN_625 = _T_634 | _GEN_619; // @[TLB.scala 68:41]
  assign _T_637 = _T_630[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_627 = _T_637 ? 6'h34 : _GEN_621; // @[TLB.scala 73:41]
  assign _GEN_628 = _T_637 | _GEN_622; // @[TLB.scala 73:41]
  assign _GEN_630 = _T_630[53] ? _GEN_624 : _GEN_618; // @[TLB.scala 67:26]
  assign _GEN_631 = _T_630[53] ? _GEN_625 : _GEN_619; // @[TLB.scala 67:26]
  assign _GEN_633 = _T_630[53] ? _GEN_627 : _GEN_621; // @[TLB.scala 67:26]
  assign _GEN_634 = _T_630[53] ? _GEN_628 : _GEN_622; // @[TLB.scala 67:26]
  assign _T_642 = tlb__T_640_data;
  assign _T_646 = _T_642[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_636 = _T_646 ? 6'h35 : _GEN_630; // @[TLB.scala 68:41]
  assign _GEN_637 = _T_646 | _GEN_631; // @[TLB.scala 68:41]
  assign _T_649 = _T_642[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_639 = _T_649 ? 6'h35 : _GEN_633; // @[TLB.scala 73:41]
  assign _GEN_640 = _T_649 | _GEN_634; // @[TLB.scala 73:41]
  assign _GEN_642 = _T_642[53] ? _GEN_636 : _GEN_630; // @[TLB.scala 67:26]
  assign _GEN_643 = _T_642[53] ? _GEN_637 : _GEN_631; // @[TLB.scala 67:26]
  assign _GEN_645 = _T_642[53] ? _GEN_639 : _GEN_633; // @[TLB.scala 67:26]
  assign _GEN_646 = _T_642[53] ? _GEN_640 : _GEN_634; // @[TLB.scala 67:26]
  assign _T_654 = tlb__T_652_data;
  assign _T_658 = _T_654[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_648 = _T_658 ? 6'h36 : _GEN_642; // @[TLB.scala 68:41]
  assign _GEN_649 = _T_658 | _GEN_643; // @[TLB.scala 68:41]
  assign _T_661 = _T_654[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_651 = _T_661 ? 6'h36 : _GEN_645; // @[TLB.scala 73:41]
  assign _GEN_652 = _T_661 | _GEN_646; // @[TLB.scala 73:41]
  assign _GEN_654 = _T_654[53] ? _GEN_648 : _GEN_642; // @[TLB.scala 67:26]
  assign _GEN_655 = _T_654[53] ? _GEN_649 : _GEN_643; // @[TLB.scala 67:26]
  assign _GEN_657 = _T_654[53] ? _GEN_651 : _GEN_645; // @[TLB.scala 67:26]
  assign _GEN_658 = _T_654[53] ? _GEN_652 : _GEN_646; // @[TLB.scala 67:26]
  assign _T_666 = tlb__T_664_data;
  assign _T_670 = _T_666[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_660 = _T_670 ? 6'h37 : _GEN_654; // @[TLB.scala 68:41]
  assign _GEN_661 = _T_670 | _GEN_655; // @[TLB.scala 68:41]
  assign _T_673 = _T_666[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_663 = _T_673 ? 6'h37 : _GEN_657; // @[TLB.scala 73:41]
  assign _GEN_664 = _T_673 | _GEN_658; // @[TLB.scala 73:41]
  assign _GEN_666 = _T_666[53] ? _GEN_660 : _GEN_654; // @[TLB.scala 67:26]
  assign _GEN_667 = _T_666[53] ? _GEN_661 : _GEN_655; // @[TLB.scala 67:26]
  assign _GEN_669 = _T_666[53] ? _GEN_663 : _GEN_657; // @[TLB.scala 67:26]
  assign _GEN_670 = _T_666[53] ? _GEN_664 : _GEN_658; // @[TLB.scala 67:26]
  assign _T_678 = tlb__T_676_data;
  assign _T_682 = _T_678[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_672 = _T_682 ? 6'h38 : _GEN_666; // @[TLB.scala 68:41]
  assign _GEN_673 = _T_682 | _GEN_667; // @[TLB.scala 68:41]
  assign _T_685 = _T_678[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_675 = _T_685 ? 6'h38 : _GEN_669; // @[TLB.scala 73:41]
  assign _GEN_676 = _T_685 | _GEN_670; // @[TLB.scala 73:41]
  assign _GEN_678 = _T_678[53] ? _GEN_672 : _GEN_666; // @[TLB.scala 67:26]
  assign _GEN_679 = _T_678[53] ? _GEN_673 : _GEN_667; // @[TLB.scala 67:26]
  assign _GEN_681 = _T_678[53] ? _GEN_675 : _GEN_669; // @[TLB.scala 67:26]
  assign _GEN_682 = _T_678[53] ? _GEN_676 : _GEN_670; // @[TLB.scala 67:26]
  assign _T_690 = tlb__T_688_data;
  assign _T_694 = _T_690[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_684 = _T_694 ? 6'h39 : _GEN_678; // @[TLB.scala 68:41]
  assign _GEN_685 = _T_694 | _GEN_679; // @[TLB.scala 68:41]
  assign _T_697 = _T_690[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_687 = _T_697 ? 6'h39 : _GEN_681; // @[TLB.scala 73:41]
  assign _GEN_688 = _T_697 | _GEN_682; // @[TLB.scala 73:41]
  assign _GEN_690 = _T_690[53] ? _GEN_684 : _GEN_678; // @[TLB.scala 67:26]
  assign _GEN_691 = _T_690[53] ? _GEN_685 : _GEN_679; // @[TLB.scala 67:26]
  assign _GEN_693 = _T_690[53] ? _GEN_687 : _GEN_681; // @[TLB.scala 67:26]
  assign _GEN_694 = _T_690[53] ? _GEN_688 : _GEN_682; // @[TLB.scala 67:26]
  assign _T_702 = tlb__T_700_data;
  assign _T_706 = _T_702[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_696 = _T_706 ? 6'h3a : _GEN_690; // @[TLB.scala 68:41]
  assign _GEN_697 = _T_706 | _GEN_691; // @[TLB.scala 68:41]
  assign _T_709 = _T_702[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_699 = _T_709 ? 6'h3a : _GEN_693; // @[TLB.scala 73:41]
  assign _GEN_700 = _T_709 | _GEN_694; // @[TLB.scala 73:41]
  assign _GEN_702 = _T_702[53] ? _GEN_696 : _GEN_690; // @[TLB.scala 67:26]
  assign _GEN_703 = _T_702[53] ? _GEN_697 : _GEN_691; // @[TLB.scala 67:26]
  assign _GEN_705 = _T_702[53] ? _GEN_699 : _GEN_693; // @[TLB.scala 67:26]
  assign _GEN_706 = _T_702[53] ? _GEN_700 : _GEN_694; // @[TLB.scala 67:26]
  assign _T_714 = tlb__T_712_data;
  assign _T_718 = _T_714[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_708 = _T_718 ? 6'h3b : _GEN_702; // @[TLB.scala 68:41]
  assign _GEN_709 = _T_718 | _GEN_703; // @[TLB.scala 68:41]
  assign _T_721 = _T_714[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_711 = _T_721 ? 6'h3b : _GEN_705; // @[TLB.scala 73:41]
  assign _GEN_712 = _T_721 | _GEN_706; // @[TLB.scala 73:41]
  assign _GEN_714 = _T_714[53] ? _GEN_708 : _GEN_702; // @[TLB.scala 67:26]
  assign _GEN_715 = _T_714[53] ? _GEN_709 : _GEN_703; // @[TLB.scala 67:26]
  assign _GEN_717 = _T_714[53] ? _GEN_711 : _GEN_705; // @[TLB.scala 67:26]
  assign _GEN_718 = _T_714[53] ? _GEN_712 : _GEN_706; // @[TLB.scala 67:26]
  assign _T_726 = tlb__T_724_data;
  assign _T_730 = _T_726[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_720 = _T_730 ? 6'h3c : _GEN_714; // @[TLB.scala 68:41]
  assign _GEN_721 = _T_730 | _GEN_715; // @[TLB.scala 68:41]
  assign _T_733 = _T_726[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_723 = _T_733 ? 6'h3c : _GEN_717; // @[TLB.scala 73:41]
  assign _GEN_724 = _T_733 | _GEN_718; // @[TLB.scala 73:41]
  assign _GEN_726 = _T_726[53] ? _GEN_720 : _GEN_714; // @[TLB.scala 67:26]
  assign _GEN_727 = _T_726[53] ? _GEN_721 : _GEN_715; // @[TLB.scala 67:26]
  assign _GEN_729 = _T_726[53] ? _GEN_723 : _GEN_717; // @[TLB.scala 67:26]
  assign _GEN_730 = _T_726[53] ? _GEN_724 : _GEN_718; // @[TLB.scala 67:26]
  assign _T_738 = tlb__T_736_data;
  assign _T_742 = _T_738[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_732 = _T_742 ? 6'h3d : _GEN_726; // @[TLB.scala 68:41]
  assign _GEN_733 = _T_742 | _GEN_727; // @[TLB.scala 68:41]
  assign _T_745 = _T_738[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_735 = _T_745 ? 6'h3d : _GEN_729; // @[TLB.scala 73:41]
  assign _GEN_736 = _T_745 | _GEN_730; // @[TLB.scala 73:41]
  assign _GEN_738 = _T_738[53] ? _GEN_732 : _GEN_726; // @[TLB.scala 67:26]
  assign _GEN_739 = _T_738[53] ? _GEN_733 : _GEN_727; // @[TLB.scala 67:26]
  assign _GEN_741 = _T_738[53] ? _GEN_735 : _GEN_729; // @[TLB.scala 67:26]
  assign _GEN_742 = _T_738[53] ? _GEN_736 : _GEN_730; // @[TLB.scala 67:26]
  assign _T_750 = tlb__T_748_data;
  assign _T_754 = _T_750[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_744 = _T_754 ? 6'h3e : _GEN_738; // @[TLB.scala 68:41]
  assign _GEN_745 = _T_754 | _GEN_739; // @[TLB.scala 68:41]
  assign _T_757 = _T_750[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_747 = _T_757 ? 6'h3e : _GEN_741; // @[TLB.scala 73:41]
  assign _GEN_748 = _T_757 | _GEN_742; // @[TLB.scala 73:41]
  assign _GEN_750 = _T_750[53] ? _GEN_744 : _GEN_738; // @[TLB.scala 67:26]
  assign _GEN_751 = _T_750[53] ? _GEN_745 : _GEN_739; // @[TLB.scala 67:26]
  assign _GEN_753 = _T_750[53] ? _GEN_747 : _GEN_741; // @[TLB.scala 67:26]
  assign _GEN_754 = _T_750[53] ? _GEN_748 : _GEN_742; // @[TLB.scala 67:26]
  assign _T_762 = tlb__T_760_data;
  assign _T_766 = _T_762[51:0] == iPortTagIn; // @[TLB.scala 68:25]
  assign _GEN_756 = _T_766 ? 6'h3f : _GEN_750; // @[TLB.scala 68:41]
  assign _GEN_757 = _T_766 | _GEN_751; // @[TLB.scala 68:41]
  assign _T_769 = _T_762[51:0] == dPortTagIn; // @[TLB.scala 73:25]
  assign _GEN_759 = _T_769 ? 6'h3f : _GEN_753; // @[TLB.scala 73:41]
  assign _GEN_760 = _T_769 | _GEN_754; // @[TLB.scala 73:41]
  assign iPortIdx = _T_762[53] ? _GEN_756 : _GEN_750; // @[TLB.scala 67:26]
  assign iPortHit = _T_762[53] ? _GEN_757 : _GEN_751; // @[TLB.scala 67:26]
  assign dPortIdx = _T_762[53] ? _GEN_759 : _GEN_753; // @[TLB.scala 67:26]
  assign dPortHit = _T_762[53] ? _GEN_760 : _GEN_754; // @[TLB.scala 67:26]
  assign _T_774 = {{3'd0}, io_iPort_vaddr_bits[63:3]}; // @[TLB.scala 87:56]
  assign _T_776 = {iPortIdx,_T_774[8:0]}; // @[Cat.scala 29:58]
  assign _T_777 = {{3'd0}, io_dPort_vaddr_bits[63:3]}; // @[TLB.scala 88:56]
  assign _T_779 = {dPortIdx,_T_777[8:0]}; // @[Cat.scala 29:58]
  assign _T_781 = ~lru_io_lru_idx[5]; // @[TLB.scala 90:28]
  assign pseudoLRU_idx2 = {_T_781,lru_io_lru_idx[4:0]}; // @[Cat.scala 29:58]
  assign _T_784 = ~iPortHit; // @[TLB.scala 95:26]
  assign _T_786 = ~dPortHit; // @[TLB.scala 96:26]
  assign io_iPort_paddr = {{49'd0}, _T_776}; // @[TLB.scala 87:18]
  assign io_iPort_miss_valid = _T_784 & io_iPort_vaddr_valid; // @[TLB.scala 95:23]
  assign io_iPort_miss_bits_vaddr = io_iPort_vaddr_bits; // @[TLB.scala 93:28]
  assign io_iPort_miss_bits_tlbIdx = io_dPort_miss_valid ? pseudoLRU_idx2 : lru_io_lru_idx; // @[TLB.scala 91:29]
  assign io_dPort_paddr = {{49'd0}, _T_779}; // @[TLB.scala 88:18]
  assign io_dPort_miss_valid = _T_786 & io_dPort_vaddr_valid; // @[TLB.scala 96:23]
  assign io_dPort_miss_bits_vaddr = io_dPort_vaddr_bits; // @[TLB.scala 94:28]
  assign io_dPort_miss_bits_tlbIdx = lru_io_lru_idx; // @[TLB.scala 92:29]
  assign lru_clock = clock;
  assign lru_reset = reset;
  assign lru_io_idx_1_valid = iPortHit & io_iPort_vaddr_valid; // @[TLB.scala 84:22]
  assign lru_io_idx_1_bits = _T_762[53] ? _GEN_756 : _GEN_750; // @[TLB.scala 82:21]
  assign lru_io_idx_2_valid = dPortHit & io_dPort_vaddr_valid; // @[TLB.scala 85:22]
  assign lru_io_idx_2_bits = _T_762[53] ? _GEN_759 : _GEN_753; // @[TLB.scala 83:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tlb[initvar] = _RAND_0[53:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tlb__T_788_en & tlb__T_788_mask) begin
      tlb[tlb__T_788_addr] <= tlb__T_788_data; // @[TLB.scala 53:16]
    end
  end
endmodule
