module DecodeUnit(
  input  [31:0] io_finst_inst,
  input         io_finst_tag,
  input  [63:0] io_finst_pc,
  output        io_dinst_rd_valid,
  output [4:0]  io_dinst_rd_bits,
  output [4:0]  io_dinst_rs1,
  output [4:0]  io_dinst_rs2,
  output [25:0] io_dinst_imm,
  output        io_dinst_shift_val_valid,
  output [5:0]  io_dinst_shift_val_bits,
  output [1:0]  io_dinst_shift_type,
  output        io_dinst_cond_valid,
  output [3:0]  io_dinst_cond_bits,
  output        io_dinst_is32bit,
  output [4:0]  io_dinst_itype,
  output [3:0]  io_dinst_op,
  output        io_dinst_nzcv_valid,
  output [3:0]  io_dinst_nzcv_bits,
  output        io_dinst_tag,
  output        io_dinst_inst32_valid,
  output [31:0] io_dinst_inst32_bits,
  output [63:0] io_dinst_pc
);
  wire [31:0] _T_1; // @[Lookup.scala 31:38]
  wire  _T_2; // @[Lookup.scala 31:38]
  wire  _T_4; // @[Lookup.scala 31:38]
  wire [31:0] _T_5; // @[Lookup.scala 31:38]
  wire  _T_6; // @[Lookup.scala 31:38]
  wire [31:0] _T_7; // @[Lookup.scala 31:38]
  wire  _T_8; // @[Lookup.scala 31:38]
  wire  _T_10; // @[Lookup.scala 31:38]
  wire  _T_12; // @[Lookup.scala 31:38]
  wire  _T_14; // @[Lookup.scala 31:38]
  wire  _T_16; // @[Lookup.scala 31:38]
  wire  _T_18; // @[Lookup.scala 31:38]
  wire  _T_20; // @[Lookup.scala 31:38]
  wire  _T_22; // @[Lookup.scala 31:38]
  wire  _T_24; // @[Lookup.scala 31:38]
  wire  _T_26; // @[Lookup.scala 31:38]
  wire  _T_28; // @[Lookup.scala 31:38]
  wire  _T_30; // @[Lookup.scala 31:38]
  wire  _T_32; // @[Lookup.scala 31:38]
  wire  _T_34; // @[Lookup.scala 31:38]
  wire  _T_36; // @[Lookup.scala 31:38]
  wire  _T_38; // @[Lookup.scala 31:38]
  wire  _T_40; // @[Lookup.scala 31:38]
  wire [31:0] _T_41; // @[Lookup.scala 31:38]
  wire  _T_42; // @[Lookup.scala 31:38]
  wire [31:0] _T_43; // @[Lookup.scala 31:38]
  wire  _T_44; // @[Lookup.scala 31:38]
  wire  _T_46; // @[Lookup.scala 31:38]
  wire  _T_48; // @[Lookup.scala 31:38]
  wire  _T_50; // @[Lookup.scala 31:38]
  wire [31:0] _T_51; // @[Lookup.scala 31:38]
  wire  _T_52; // @[Lookup.scala 31:38]
  wire [31:0] _T_53; // @[Lookup.scala 31:38]
  wire  _T_54; // @[Lookup.scala 31:38]
  wire  _T_56; // @[Lookup.scala 31:38]
  wire  _T_58; // @[Lookup.scala 31:38]
  wire  _T_60; // @[Lookup.scala 31:38]
  wire  _T_62; // @[Lookup.scala 31:38]
  wire  _T_64; // @[Lookup.scala 31:38]
  wire  _T_66; // @[Lookup.scala 31:38]
  wire  _T_68; // @[Lookup.scala 31:38]
  wire  _T_70; // @[Lookup.scala 31:38]
  wire  _T_72; // @[Lookup.scala 31:38]
  wire  _T_74; // @[Lookup.scala 31:38]
  wire  _T_76; // @[Lookup.scala 31:38]
  wire  _T_78; // @[Lookup.scala 31:38]
  wire  _T_80; // @[Lookup.scala 31:38]
  wire  _T_82; // @[Lookup.scala 31:38]
  wire  _T_84; // @[Lookup.scala 31:38]
  wire [31:0] _T_85; // @[Lookup.scala 31:38]
  wire  _T_86; // @[Lookup.scala 31:38]
  wire  _T_88; // @[Lookup.scala 31:38]
  wire  _T_90; // @[Lookup.scala 31:38]
  wire  _T_92; // @[Lookup.scala 31:38]
  wire  _T_94; // @[Lookup.scala 31:38]
  wire  _T_96; // @[Lookup.scala 31:38]
  wire  _T_98; // @[Lookup.scala 31:38]
  wire  _T_100; // @[Lookup.scala 31:38]
  wire [31:0] _T_101; // @[Lookup.scala 31:38]
  wire  _T_102; // @[Lookup.scala 31:38]
  wire  _T_104; // @[Lookup.scala 31:38]
  wire  _T_106; // @[Lookup.scala 31:38]
  wire  _T_108; // @[Lookup.scala 31:38]
  wire  _T_110; // @[Lookup.scala 31:38]
  wire  _T_112; // @[Lookup.scala 31:38]
  wire  _T_114; // @[Lookup.scala 31:38]
  wire  _T_116; // @[Lookup.scala 31:38]
  wire  _T_118; // @[Lookup.scala 31:38]
  wire  _T_120; // @[Lookup.scala 31:38]
  wire  _T_122; // @[Lookup.scala 31:38]
  wire  _T_124; // @[Lookup.scala 31:38]
  wire  _T_126; // @[Lookup.scala 31:38]
  wire  _T_128; // @[Lookup.scala 31:38]
  wire  _T_130; // @[Lookup.scala 31:38]
  wire  _T_132; // @[Lookup.scala 31:38]
  wire  _T_134; // @[Lookup.scala 31:38]
  wire  _T_136; // @[Lookup.scala 31:38]
  wire  _T_138; // @[Lookup.scala 31:38]
  wire  _T_140; // @[Lookup.scala 31:38]
  wire  _T_142; // @[Lookup.scala 31:38]
  wire  _T_144; // @[Lookup.scala 31:38]
  wire  _T_146; // @[Lookup.scala 31:38]
  wire  _T_148; // @[Lookup.scala 31:38]
  wire  _T_150; // @[Lookup.scala 31:38]
  wire  _T_152; // @[Lookup.scala 31:38]
  wire  _T_154; // @[Lookup.scala 31:38]
  wire  _T_156; // @[Lookup.scala 31:38]
  wire  _T_158; // @[Lookup.scala 31:38]
  wire  _T_160; // @[Lookup.scala 31:38]
  wire [31:0] _T_161; // @[Lookup.scala 31:38]
  wire  _T_162; // @[Lookup.scala 31:38]
  wire  _T_164; // @[Lookup.scala 31:38]
  wire  _T_166; // @[Lookup.scala 31:38]
  wire  _T_168; // @[Lookup.scala 31:38]
  wire  _T_170; // @[Lookup.scala 31:38]
  wire  _T_172; // @[Lookup.scala 31:38]
  wire  _T_174; // @[Lookup.scala 31:38]
  wire  _T_176; // @[Lookup.scala 31:38]
  wire  _T_178; // @[Lookup.scala 31:38]
  wire  _T_180; // @[Lookup.scala 31:38]
  wire  _T_182; // @[Lookup.scala 31:38]
  wire [31:0] _T_183; // @[Lookup.scala 31:38]
  wire  _T_184; // @[Lookup.scala 31:38]
  wire  _T_186; // @[Lookup.scala 31:38]
  wire  _T_188; // @[Lookup.scala 31:38]
  wire  _T_190; // @[Lookup.scala 31:38]
  wire  _T_192; // @[Lookup.scala 31:38]
  wire  _T_194; // @[Lookup.scala 31:38]
  wire  _T_196; // @[Lookup.scala 31:38]
  wire  _T_198; // @[Lookup.scala 31:38]
  wire [31:0] _T_199; // @[Lookup.scala 31:38]
  wire  _T_200; // @[Lookup.scala 31:38]
  wire [31:0] _T_201; // @[Lookup.scala 31:38]
  wire  _T_202; // @[Lookup.scala 31:38]
  wire  _T_204; // @[Lookup.scala 31:38]
  wire [31:0] _T_205; // @[Lookup.scala 31:38]
  wire  _T_206; // @[Lookup.scala 31:38]
  wire  _T_208; // @[Lookup.scala 31:38]
  wire  _T_210; // @[Lookup.scala 31:38]
  wire [31:0] _T_211; // @[Lookup.scala 31:38]
  wire  _T_212; // @[Lookup.scala 31:38]
  wire  _T_214; // @[Lookup.scala 31:38]
  wire  _T_216; // @[Lookup.scala 31:38]
  wire  _T_218; // @[Lookup.scala 31:38]
  wire [31:0] _T_219; // @[Lookup.scala 31:38]
  wire  _T_220; // @[Lookup.scala 31:38]
  wire  _T_222; // @[Lookup.scala 31:38]
  wire  _T_224; // @[Lookup.scala 31:38]
  wire  _T_226; // @[Lookup.scala 31:38]
  wire  _T_228; // @[Lookup.scala 31:38]
  wire  _T_230; // @[Lookup.scala 31:38]
  wire  _T_232; // @[Lookup.scala 31:38]
  wire  _T_234; // @[Lookup.scala 31:38]
  wire  _T_236; // @[Lookup.scala 31:38]
  wire  _T_238; // @[Lookup.scala 31:38]
  wire  _T_240; // @[Lookup.scala 31:38]
  wire  _T_242; // @[Lookup.scala 31:38]
  wire  _T_244; // @[Lookup.scala 31:38]
  wire  _T_246; // @[Lookup.scala 31:38]
  wire  _T_248; // @[Lookup.scala 31:38]
  wire  _T_250; // @[Lookup.scala 31:38]
  wire  _T_252; // @[Lookup.scala 31:38]
  wire  _T_254; // @[Lookup.scala 31:38]
  wire  _T_256; // @[Lookup.scala 31:38]
  wire  _T_258; // @[Lookup.scala 31:38]
  wire [31:0] _T_259; // @[Lookup.scala 31:38]
  wire  _T_260; // @[Lookup.scala 31:38]
  wire  _T_262; // @[Lookup.scala 31:38]
  wire  _T_264; // @[Lookup.scala 31:38]
  wire  _T_266; // @[Lookup.scala 31:38]
  wire  _T_268; // @[Lookup.scala 31:38]
  wire  _T_270; // @[Lookup.scala 31:38]
  wire  _T_272; // @[Lookup.scala 31:38]
  wire  _T_274; // @[Lookup.scala 31:38]
  wire  _T_276; // @[Lookup.scala 31:38]
  wire  _T_278; // @[Lookup.scala 31:38]
  wire  _T_280; // @[Lookup.scala 31:38]
  wire  _T_282; // @[Lookup.scala 31:38]
  wire  _T_284; // @[Lookup.scala 31:38]
  wire  _T_286; // @[Lookup.scala 31:38]
  wire  _T_288; // @[Lookup.scala 31:38]
  wire  _T_290; // @[Lookup.scala 31:38]
  wire  _T_292; // @[Lookup.scala 31:38]
  wire  _T_294; // @[Lookup.scala 31:38]
  wire  _T_296; // @[Lookup.scala 31:38]
  wire  _T_298; // @[Lookup.scala 31:38]
  wire  _T_300; // @[Lookup.scala 31:38]
  wire  _T_302; // @[Lookup.scala 31:38]
  wire  _T_304; // @[Lookup.scala 31:38]
  wire  _T_306; // @[Lookup.scala 31:38]
  wire  _T_308; // @[Lookup.scala 31:38]
  wire  _T_310; // @[Lookup.scala 31:38]
  wire  _T_312; // @[Lookup.scala 31:38]
  wire  _T_314; // @[Lookup.scala 31:38]
  wire  _T_316; // @[Lookup.scala 31:38]
  wire  _T_318; // @[Lookup.scala 31:38]
  wire  _T_320; // @[Lookup.scala 31:38]
  wire  _T_322; // @[Lookup.scala 31:38]
  wire  _T_324; // @[Lookup.scala 31:38]
  wire  _T_326; // @[Lookup.scala 31:38]
  wire  _T_328; // @[Lookup.scala 31:38]
  wire  _T_330; // @[Lookup.scala 31:38]
  wire  _T_332; // @[Lookup.scala 31:38]
  wire  _T_334; // @[Lookup.scala 31:38]
  wire  _T_336; // @[Lookup.scala 31:38]
  wire  _T_338; // @[Lookup.scala 31:38]
  wire  _T_340; // @[Lookup.scala 31:38]
  wire  _T_342; // @[Lookup.scala 31:38]
  wire  _T_344; // @[Lookup.scala 31:38]
  wire  _T_346; // @[Lookup.scala 31:38]
  wire  _T_348; // @[Lookup.scala 31:38]
  wire  _T_350; // @[Lookup.scala 31:38]
  wire  _T_352; // @[Lookup.scala 31:38]
  wire  _T_354; // @[Lookup.scala 31:38]
  wire  _T_356; // @[Lookup.scala 31:38]
  wire  _T_358; // @[Lookup.scala 31:38]
  wire  _T_360; // @[Lookup.scala 31:38]
  wire  _T_362; // @[Lookup.scala 31:38]
  wire  _T_364; // @[Lookup.scala 31:38]
  wire  _T_366; // @[Lookup.scala 31:38]
  wire  _T_368; // @[Lookup.scala 31:38]
  wire  _T_370; // @[Lookup.scala 31:38]
  wire  _T_372; // @[Lookup.scala 31:38]
  wire  _T_374; // @[Lookup.scala 31:38]
  wire  _T_376; // @[Lookup.scala 31:38]
  wire  _T_378; // @[Lookup.scala 31:38]
  wire [4:0] _T_379; // @[Lookup.scala 33:37]
  wire [4:0] _T_380; // @[Lookup.scala 33:37]
  wire [4:0] _T_381; // @[Lookup.scala 33:37]
  wire [4:0] _T_382; // @[Lookup.scala 33:37]
  wire [4:0] _T_383; // @[Lookup.scala 33:37]
  wire [4:0] _T_384; // @[Lookup.scala 33:37]
  wire [4:0] _T_385; // @[Lookup.scala 33:37]
  wire [4:0] _T_386; // @[Lookup.scala 33:37]
  wire [4:0] _T_387; // @[Lookup.scala 33:37]
  wire [4:0] _T_388; // @[Lookup.scala 33:37]
  wire [4:0] _T_389; // @[Lookup.scala 33:37]
  wire [4:0] _T_390; // @[Lookup.scala 33:37]
  wire [4:0] _T_391; // @[Lookup.scala 33:37]
  wire [4:0] _T_392; // @[Lookup.scala 33:37]
  wire [4:0] _T_393; // @[Lookup.scala 33:37]
  wire [4:0] _T_394; // @[Lookup.scala 33:37]
  wire [4:0] _T_395; // @[Lookup.scala 33:37]
  wire [4:0] _T_396; // @[Lookup.scala 33:37]
  wire [4:0] _T_397; // @[Lookup.scala 33:37]
  wire [4:0] _T_398; // @[Lookup.scala 33:37]
  wire [4:0] _T_399; // @[Lookup.scala 33:37]
  wire [4:0] _T_400; // @[Lookup.scala 33:37]
  wire [4:0] _T_401; // @[Lookup.scala 33:37]
  wire [4:0] _T_402; // @[Lookup.scala 33:37]
  wire [4:0] _T_403; // @[Lookup.scala 33:37]
  wire [4:0] _T_404; // @[Lookup.scala 33:37]
  wire [4:0] _T_405; // @[Lookup.scala 33:37]
  wire [4:0] _T_406; // @[Lookup.scala 33:37]
  wire [4:0] _T_407; // @[Lookup.scala 33:37]
  wire [4:0] _T_408; // @[Lookup.scala 33:37]
  wire [4:0] _T_409; // @[Lookup.scala 33:37]
  wire [4:0] _T_410; // @[Lookup.scala 33:37]
  wire [4:0] _T_411; // @[Lookup.scala 33:37]
  wire [4:0] _T_412; // @[Lookup.scala 33:37]
  wire [4:0] _T_413; // @[Lookup.scala 33:37]
  wire [4:0] _T_414; // @[Lookup.scala 33:37]
  wire [4:0] _T_415; // @[Lookup.scala 33:37]
  wire [4:0] _T_416; // @[Lookup.scala 33:37]
  wire [4:0] _T_417; // @[Lookup.scala 33:37]
  wire [4:0] _T_418; // @[Lookup.scala 33:37]
  wire [4:0] _T_419; // @[Lookup.scala 33:37]
  wire [4:0] _T_420; // @[Lookup.scala 33:37]
  wire [4:0] _T_421; // @[Lookup.scala 33:37]
  wire [4:0] _T_422; // @[Lookup.scala 33:37]
  wire [4:0] _T_423; // @[Lookup.scala 33:37]
  wire [4:0] _T_424; // @[Lookup.scala 33:37]
  wire [4:0] _T_425; // @[Lookup.scala 33:37]
  wire [4:0] _T_426; // @[Lookup.scala 33:37]
  wire [4:0] _T_427; // @[Lookup.scala 33:37]
  wire [4:0] _T_428; // @[Lookup.scala 33:37]
  wire [4:0] _T_429; // @[Lookup.scala 33:37]
  wire [4:0] _T_430; // @[Lookup.scala 33:37]
  wire [4:0] _T_431; // @[Lookup.scala 33:37]
  wire [4:0] _T_432; // @[Lookup.scala 33:37]
  wire [4:0] _T_433; // @[Lookup.scala 33:37]
  wire [4:0] _T_434; // @[Lookup.scala 33:37]
  wire [4:0] _T_435; // @[Lookup.scala 33:37]
  wire [4:0] _T_436; // @[Lookup.scala 33:37]
  wire [4:0] _T_437; // @[Lookup.scala 33:37]
  wire [4:0] _T_438; // @[Lookup.scala 33:37]
  wire [4:0] _T_439; // @[Lookup.scala 33:37]
  wire [4:0] _T_440; // @[Lookup.scala 33:37]
  wire [4:0] _T_441; // @[Lookup.scala 33:37]
  wire [4:0] _T_442; // @[Lookup.scala 33:37]
  wire [4:0] _T_443; // @[Lookup.scala 33:37]
  wire [4:0] _T_444; // @[Lookup.scala 33:37]
  wire [4:0] _T_445; // @[Lookup.scala 33:37]
  wire [4:0] _T_446; // @[Lookup.scala 33:37]
  wire [4:0] _T_447; // @[Lookup.scala 33:37]
  wire [4:0] _T_448; // @[Lookup.scala 33:37]
  wire [4:0] _T_449; // @[Lookup.scala 33:37]
  wire [4:0] _T_450; // @[Lookup.scala 33:37]
  wire [4:0] _T_451; // @[Lookup.scala 33:37]
  wire [4:0] _T_452; // @[Lookup.scala 33:37]
  wire [4:0] _T_453; // @[Lookup.scala 33:37]
  wire [4:0] _T_454; // @[Lookup.scala 33:37]
  wire [4:0] _T_455; // @[Lookup.scala 33:37]
  wire [4:0] _T_456; // @[Lookup.scala 33:37]
  wire [4:0] _T_457; // @[Lookup.scala 33:37]
  wire [4:0] _T_458; // @[Lookup.scala 33:37]
  wire [4:0] _T_459; // @[Lookup.scala 33:37]
  wire [4:0] _T_460; // @[Lookup.scala 33:37]
  wire [4:0] _T_461; // @[Lookup.scala 33:37]
  wire [4:0] _T_462; // @[Lookup.scala 33:37]
  wire [4:0] _T_463; // @[Lookup.scala 33:37]
  wire [4:0] _T_464; // @[Lookup.scala 33:37]
  wire [4:0] _T_465; // @[Lookup.scala 33:37]
  wire [4:0] _T_466; // @[Lookup.scala 33:37]
  wire [4:0] _T_467; // @[Lookup.scala 33:37]
  wire [4:0] _T_468; // @[Lookup.scala 33:37]
  wire [4:0] _T_469; // @[Lookup.scala 33:37]
  wire [4:0] _T_470; // @[Lookup.scala 33:37]
  wire [4:0] _T_471; // @[Lookup.scala 33:37]
  wire [4:0] _T_472; // @[Lookup.scala 33:37]
  wire [4:0] _T_473; // @[Lookup.scala 33:37]
  wire [4:0] _T_474; // @[Lookup.scala 33:37]
  wire [4:0] _T_475; // @[Lookup.scala 33:37]
  wire [4:0] _T_476; // @[Lookup.scala 33:37]
  wire [4:0] _T_477; // @[Lookup.scala 33:37]
  wire [4:0] _T_478; // @[Lookup.scala 33:37]
  wire [4:0] _T_479; // @[Lookup.scala 33:37]
  wire [4:0] _T_480; // @[Lookup.scala 33:37]
  wire [4:0] _T_481; // @[Lookup.scala 33:37]
  wire [4:0] _T_482; // @[Lookup.scala 33:37]
  wire [4:0] _T_483; // @[Lookup.scala 33:37]
  wire [4:0] _T_484; // @[Lookup.scala 33:37]
  wire [4:0] _T_485; // @[Lookup.scala 33:37]
  wire [4:0] _T_486; // @[Lookup.scala 33:37]
  wire [4:0] _T_487; // @[Lookup.scala 33:37]
  wire [4:0] _T_488; // @[Lookup.scala 33:37]
  wire [4:0] _T_489; // @[Lookup.scala 33:37]
  wire [4:0] _T_490; // @[Lookup.scala 33:37]
  wire [4:0] _T_491; // @[Lookup.scala 33:37]
  wire [4:0] _T_492; // @[Lookup.scala 33:37]
  wire [4:0] _T_493; // @[Lookup.scala 33:37]
  wire [4:0] _T_494; // @[Lookup.scala 33:37]
  wire [4:0] _T_495; // @[Lookup.scala 33:37]
  wire [4:0] _T_496; // @[Lookup.scala 33:37]
  wire [4:0] _T_497; // @[Lookup.scala 33:37]
  wire [4:0] _T_498; // @[Lookup.scala 33:37]
  wire [4:0] _T_499; // @[Lookup.scala 33:37]
  wire [4:0] _T_500; // @[Lookup.scala 33:37]
  wire [4:0] _T_501; // @[Lookup.scala 33:37]
  wire [4:0] _T_502; // @[Lookup.scala 33:37]
  wire [4:0] _T_503; // @[Lookup.scala 33:37]
  wire [4:0] _T_504; // @[Lookup.scala 33:37]
  wire [4:0] _T_505; // @[Lookup.scala 33:37]
  wire [4:0] _T_506; // @[Lookup.scala 33:37]
  wire [4:0] _T_507; // @[Lookup.scala 33:37]
  wire [4:0] _T_508; // @[Lookup.scala 33:37]
  wire [4:0] _T_509; // @[Lookup.scala 33:37]
  wire [4:0] _T_510; // @[Lookup.scala 33:37]
  wire [4:0] _T_511; // @[Lookup.scala 33:37]
  wire [4:0] _T_512; // @[Lookup.scala 33:37]
  wire [4:0] _T_513; // @[Lookup.scala 33:37]
  wire [4:0] _T_514; // @[Lookup.scala 33:37]
  wire [4:0] _T_515; // @[Lookup.scala 33:37]
  wire [4:0] _T_516; // @[Lookup.scala 33:37]
  wire [4:0] _T_517; // @[Lookup.scala 33:37]
  wire [4:0] _T_518; // @[Lookup.scala 33:37]
  wire [4:0] _T_519; // @[Lookup.scala 33:37]
  wire [4:0] _T_520; // @[Lookup.scala 33:37]
  wire [4:0] _T_521; // @[Lookup.scala 33:37]
  wire [4:0] _T_522; // @[Lookup.scala 33:37]
  wire [4:0] _T_523; // @[Lookup.scala 33:37]
  wire [4:0] _T_524; // @[Lookup.scala 33:37]
  wire [4:0] _T_525; // @[Lookup.scala 33:37]
  wire [4:0] _T_526; // @[Lookup.scala 33:37]
  wire [4:0] _T_527; // @[Lookup.scala 33:37]
  wire [4:0] _T_528; // @[Lookup.scala 33:37]
  wire [4:0] _T_529; // @[Lookup.scala 33:37]
  wire [4:0] _T_530; // @[Lookup.scala 33:37]
  wire [4:0] _T_531; // @[Lookup.scala 33:37]
  wire [4:0] _T_532; // @[Lookup.scala 33:37]
  wire [4:0] _T_533; // @[Lookup.scala 33:37]
  wire [4:0] _T_534; // @[Lookup.scala 33:37]
  wire [4:0] _T_535; // @[Lookup.scala 33:37]
  wire [4:0] _T_536; // @[Lookup.scala 33:37]
  wire [4:0] _T_537; // @[Lookup.scala 33:37]
  wire [4:0] _T_538; // @[Lookup.scala 33:37]
  wire [4:0] _T_539; // @[Lookup.scala 33:37]
  wire [4:0] _T_540; // @[Lookup.scala 33:37]
  wire [4:0] _T_541; // @[Lookup.scala 33:37]
  wire [4:0] _T_542; // @[Lookup.scala 33:37]
  wire [4:0] _T_543; // @[Lookup.scala 33:37]
  wire [4:0] _T_544; // @[Lookup.scala 33:37]
  wire [4:0] _T_545; // @[Lookup.scala 33:37]
  wire [4:0] _T_546; // @[Lookup.scala 33:37]
  wire [4:0] _T_547; // @[Lookup.scala 33:37]
  wire [4:0] _T_548; // @[Lookup.scala 33:37]
  wire [4:0] _T_549; // @[Lookup.scala 33:37]
  wire [4:0] _T_550; // @[Lookup.scala 33:37]
  wire [4:0] _T_551; // @[Lookup.scala 33:37]
  wire [4:0] _T_552; // @[Lookup.scala 33:37]
  wire [4:0] _T_553; // @[Lookup.scala 33:37]
  wire [4:0] _T_554; // @[Lookup.scala 33:37]
  wire [4:0] _T_555; // @[Lookup.scala 33:37]
  wire [4:0] _T_556; // @[Lookup.scala 33:37]
  wire [4:0] _T_557; // @[Lookup.scala 33:37]
  wire [4:0] _T_558; // @[Lookup.scala 33:37]
  wire [4:0] _T_559; // @[Lookup.scala 33:37]
  wire [4:0] _T_560; // @[Lookup.scala 33:37]
  wire [4:0] _T_561; // @[Lookup.scala 33:37]
  wire [4:0] _T_562; // @[Lookup.scala 33:37]
  wire [4:0] _T_563; // @[Lookup.scala 33:37]
  wire [4:0] _T_564; // @[Lookup.scala 33:37]
  wire [4:0] _T_565; // @[Lookup.scala 33:37]
  wire [4:0] _T_566; // @[Lookup.scala 33:37]
  wire [4:0] dinst_itype; // @[Lookup.scala 33:37]
  wire [3:0] _T_568; // @[Lookup.scala 33:37]
  wire [3:0] _T_569; // @[Lookup.scala 33:37]
  wire [3:0] _T_570; // @[Lookup.scala 33:37]
  wire [3:0] _T_571; // @[Lookup.scala 33:37]
  wire [3:0] _T_572; // @[Lookup.scala 33:37]
  wire [3:0] _T_573; // @[Lookup.scala 33:37]
  wire [3:0] _T_574; // @[Lookup.scala 33:37]
  wire [3:0] _T_575; // @[Lookup.scala 33:37]
  wire [3:0] _T_576; // @[Lookup.scala 33:37]
  wire [3:0] _T_577; // @[Lookup.scala 33:37]
  wire [3:0] _T_578; // @[Lookup.scala 33:37]
  wire [3:0] _T_579; // @[Lookup.scala 33:37]
  wire [3:0] _T_580; // @[Lookup.scala 33:37]
  wire [3:0] _T_581; // @[Lookup.scala 33:37]
  wire [3:0] _T_582; // @[Lookup.scala 33:37]
  wire [3:0] _T_583; // @[Lookup.scala 33:37]
  wire [3:0] _T_584; // @[Lookup.scala 33:37]
  wire [3:0] _T_585; // @[Lookup.scala 33:37]
  wire [3:0] _T_586; // @[Lookup.scala 33:37]
  wire [3:0] _T_587; // @[Lookup.scala 33:37]
  wire [3:0] _T_588; // @[Lookup.scala 33:37]
  wire [3:0] _T_589; // @[Lookup.scala 33:37]
  wire [3:0] _T_590; // @[Lookup.scala 33:37]
  wire [3:0] _T_591; // @[Lookup.scala 33:37]
  wire [3:0] _T_592; // @[Lookup.scala 33:37]
  wire [3:0] _T_593; // @[Lookup.scala 33:37]
  wire [3:0] _T_594; // @[Lookup.scala 33:37]
  wire [3:0] _T_595; // @[Lookup.scala 33:37]
  wire [3:0] _T_596; // @[Lookup.scala 33:37]
  wire [3:0] _T_597; // @[Lookup.scala 33:37]
  wire [3:0] _T_598; // @[Lookup.scala 33:37]
  wire [3:0] _T_599; // @[Lookup.scala 33:37]
  wire [3:0] _T_600; // @[Lookup.scala 33:37]
  wire [3:0] _T_601; // @[Lookup.scala 33:37]
  wire [3:0] _T_602; // @[Lookup.scala 33:37]
  wire [3:0] _T_603; // @[Lookup.scala 33:37]
  wire [3:0] _T_604; // @[Lookup.scala 33:37]
  wire [3:0] _T_605; // @[Lookup.scala 33:37]
  wire [3:0] _T_606; // @[Lookup.scala 33:37]
  wire [3:0] _T_607; // @[Lookup.scala 33:37]
  wire [3:0] _T_608; // @[Lookup.scala 33:37]
  wire [3:0] _T_609; // @[Lookup.scala 33:37]
  wire [3:0] _T_610; // @[Lookup.scala 33:37]
  wire [3:0] _T_611; // @[Lookup.scala 33:37]
  wire [3:0] _T_612; // @[Lookup.scala 33:37]
  wire [3:0] _T_613; // @[Lookup.scala 33:37]
  wire [3:0] _T_614; // @[Lookup.scala 33:37]
  wire [3:0] _T_615; // @[Lookup.scala 33:37]
  wire [3:0] _T_616; // @[Lookup.scala 33:37]
  wire [3:0] _T_617; // @[Lookup.scala 33:37]
  wire [3:0] _T_618; // @[Lookup.scala 33:37]
  wire [3:0] _T_619; // @[Lookup.scala 33:37]
  wire [3:0] _T_620; // @[Lookup.scala 33:37]
  wire [3:0] _T_621; // @[Lookup.scala 33:37]
  wire [3:0] _T_622; // @[Lookup.scala 33:37]
  wire [3:0] _T_623; // @[Lookup.scala 33:37]
  wire [3:0] _T_624; // @[Lookup.scala 33:37]
  wire [3:0] _T_625; // @[Lookup.scala 33:37]
  wire [3:0] _T_626; // @[Lookup.scala 33:37]
  wire [3:0] _T_627; // @[Lookup.scala 33:37]
  wire [3:0] _T_628; // @[Lookup.scala 33:37]
  wire [3:0] _T_629; // @[Lookup.scala 33:37]
  wire [3:0] _T_630; // @[Lookup.scala 33:37]
  wire [3:0] _T_631; // @[Lookup.scala 33:37]
  wire [3:0] _T_632; // @[Lookup.scala 33:37]
  wire [3:0] _T_633; // @[Lookup.scala 33:37]
  wire [3:0] _T_634; // @[Lookup.scala 33:37]
  wire [3:0] _T_635; // @[Lookup.scala 33:37]
  wire [3:0] _T_636; // @[Lookup.scala 33:37]
  wire [3:0] _T_637; // @[Lookup.scala 33:37]
  wire [3:0] _T_638; // @[Lookup.scala 33:37]
  wire [3:0] _T_639; // @[Lookup.scala 33:37]
  wire [3:0] _T_640; // @[Lookup.scala 33:37]
  wire [3:0] _T_641; // @[Lookup.scala 33:37]
  wire [3:0] _T_642; // @[Lookup.scala 33:37]
  wire [3:0] _T_643; // @[Lookup.scala 33:37]
  wire [3:0] _T_644; // @[Lookup.scala 33:37]
  wire [3:0] _T_645; // @[Lookup.scala 33:37]
  wire [3:0] _T_646; // @[Lookup.scala 33:37]
  wire [3:0] _T_647; // @[Lookup.scala 33:37]
  wire [3:0] _T_648; // @[Lookup.scala 33:37]
  wire [3:0] _T_649; // @[Lookup.scala 33:37]
  wire [3:0] _T_650; // @[Lookup.scala 33:37]
  wire [3:0] _T_651; // @[Lookup.scala 33:37]
  wire [3:0] _T_652; // @[Lookup.scala 33:37]
  wire [3:0] _T_653; // @[Lookup.scala 33:37]
  wire [3:0] _T_654; // @[Lookup.scala 33:37]
  wire [3:0] _T_655; // @[Lookup.scala 33:37]
  wire [3:0] _T_656; // @[Lookup.scala 33:37]
  wire [3:0] _T_657; // @[Lookup.scala 33:37]
  wire [3:0] _T_658; // @[Lookup.scala 33:37]
  wire [3:0] _T_659; // @[Lookup.scala 33:37]
  wire [3:0] _T_660; // @[Lookup.scala 33:37]
  wire [3:0] _T_661; // @[Lookup.scala 33:37]
  wire [3:0] _T_662; // @[Lookup.scala 33:37]
  wire [3:0] _T_663; // @[Lookup.scala 33:37]
  wire [3:0] _T_664; // @[Lookup.scala 33:37]
  wire [3:0] _T_665; // @[Lookup.scala 33:37]
  wire [3:0] _T_666; // @[Lookup.scala 33:37]
  wire [3:0] _T_667; // @[Lookup.scala 33:37]
  wire [3:0] _T_668; // @[Lookup.scala 33:37]
  wire [3:0] _T_669; // @[Lookup.scala 33:37]
  wire [3:0] _T_670; // @[Lookup.scala 33:37]
  wire [3:0] _T_671; // @[Lookup.scala 33:37]
  wire [3:0] _T_672; // @[Lookup.scala 33:37]
  wire [3:0] _T_673; // @[Lookup.scala 33:37]
  wire [3:0] _T_674; // @[Lookup.scala 33:37]
  wire [3:0] _T_675; // @[Lookup.scala 33:37]
  wire [3:0] _T_676; // @[Lookup.scala 33:37]
  wire [3:0] _T_677; // @[Lookup.scala 33:37]
  wire [3:0] _T_678; // @[Lookup.scala 33:37]
  wire [3:0] _T_679; // @[Lookup.scala 33:37]
  wire [3:0] _T_680; // @[Lookup.scala 33:37]
  wire [3:0] _T_681; // @[Lookup.scala 33:37]
  wire [3:0] _T_682; // @[Lookup.scala 33:37]
  wire [3:0] _T_683; // @[Lookup.scala 33:37]
  wire [3:0] _T_684; // @[Lookup.scala 33:37]
  wire [3:0] _T_685; // @[Lookup.scala 33:37]
  wire [3:0] _T_686; // @[Lookup.scala 33:37]
  wire [3:0] _T_687; // @[Lookup.scala 33:37]
  wire [3:0] _T_688; // @[Lookup.scala 33:37]
  wire [3:0] _T_689; // @[Lookup.scala 33:37]
  wire [3:0] _T_690; // @[Lookup.scala 33:37]
  wire [3:0] _T_691; // @[Lookup.scala 33:37]
  wire [3:0] _T_692; // @[Lookup.scala 33:37]
  wire [3:0] _T_693; // @[Lookup.scala 33:37]
  wire [3:0] _T_694; // @[Lookup.scala 33:37]
  wire [3:0] _T_695; // @[Lookup.scala 33:37]
  wire [3:0] _T_696; // @[Lookup.scala 33:37]
  wire [3:0] _T_697; // @[Lookup.scala 33:37]
  wire [3:0] _T_698; // @[Lookup.scala 33:37]
  wire [3:0] _T_699; // @[Lookup.scala 33:37]
  wire [3:0] _T_700; // @[Lookup.scala 33:37]
  wire [3:0] _T_701; // @[Lookup.scala 33:37]
  wire [3:0] _T_702; // @[Lookup.scala 33:37]
  wire [3:0] _T_703; // @[Lookup.scala 33:37]
  wire [3:0] _T_704; // @[Lookup.scala 33:37]
  wire [3:0] _T_705; // @[Lookup.scala 33:37]
  wire [3:0] _T_706; // @[Lookup.scala 33:37]
  wire [3:0] _T_707; // @[Lookup.scala 33:37]
  wire [3:0] _T_708; // @[Lookup.scala 33:37]
  wire [3:0] _T_709; // @[Lookup.scala 33:37]
  wire [3:0] _T_710; // @[Lookup.scala 33:37]
  wire [3:0] _T_711; // @[Lookup.scala 33:37]
  wire [3:0] _T_712; // @[Lookup.scala 33:37]
  wire [3:0] _T_713; // @[Lookup.scala 33:37]
  wire [3:0] _T_714; // @[Lookup.scala 33:37]
  wire [3:0] _T_715; // @[Lookup.scala 33:37]
  wire [3:0] _T_716; // @[Lookup.scala 33:37]
  wire [3:0] _T_717; // @[Lookup.scala 33:37]
  wire [3:0] _T_718; // @[Lookup.scala 33:37]
  wire [3:0] _T_719; // @[Lookup.scala 33:37]
  wire [3:0] _T_720; // @[Lookup.scala 33:37]
  wire [3:0] _T_721; // @[Lookup.scala 33:37]
  wire [3:0] _T_722; // @[Lookup.scala 33:37]
  wire [3:0] _T_723; // @[Lookup.scala 33:37]
  wire [3:0] _T_724; // @[Lookup.scala 33:37]
  wire [3:0] _T_725; // @[Lookup.scala 33:37]
  wire [3:0] _T_726; // @[Lookup.scala 33:37]
  wire [3:0] _T_727; // @[Lookup.scala 33:37]
  wire [3:0] _T_728; // @[Lookup.scala 33:37]
  wire [3:0] _T_729; // @[Lookup.scala 33:37]
  wire [3:0] _T_730; // @[Lookup.scala 33:37]
  wire [3:0] _T_731; // @[Lookup.scala 33:37]
  wire [3:0] _T_732; // @[Lookup.scala 33:37]
  wire [3:0] _T_733; // @[Lookup.scala 33:37]
  wire [3:0] _T_734; // @[Lookup.scala 33:37]
  wire [3:0] _T_735; // @[Lookup.scala 33:37]
  wire [3:0] _T_736; // @[Lookup.scala 33:37]
  wire [3:0] _T_737; // @[Lookup.scala 33:37]
  wire [3:0] _T_738; // @[Lookup.scala 33:37]
  wire [3:0] _T_739; // @[Lookup.scala 33:37]
  wire [3:0] _T_740; // @[Lookup.scala 33:37]
  wire [3:0] _T_741; // @[Lookup.scala 33:37]
  wire [3:0] _T_742; // @[Lookup.scala 33:37]
  wire [3:0] _T_743; // @[Lookup.scala 33:37]
  wire [3:0] _T_744; // @[Lookup.scala 33:37]
  wire [3:0] _T_745; // @[Lookup.scala 33:37]
  wire [3:0] _T_746; // @[Lookup.scala 33:37]
  wire [3:0] _T_747; // @[Lookup.scala 33:37]
  wire [3:0] _T_748; // @[Lookup.scala 33:37]
  wire [3:0] _T_749; // @[Lookup.scala 33:37]
  wire [3:0] _T_750; // @[Lookup.scala 33:37]
  wire [3:0] _T_751; // @[Lookup.scala 33:37]
  wire [3:0] _T_752; // @[Lookup.scala 33:37]
  wire [3:0] _T_753; // @[Lookup.scala 33:37]
  wire [3:0] _T_754; // @[Lookup.scala 33:37]
  wire [3:0] _T_755; // @[Lookup.scala 33:37]
  wire  _T_758; // @[Lookup.scala 33:37]
  wire  _T_759; // @[Lookup.scala 33:37]
  wire  _T_760; // @[Lookup.scala 33:37]
  wire  _T_761; // @[Lookup.scala 33:37]
  wire  _T_762; // @[Lookup.scala 33:37]
  wire  _T_763; // @[Lookup.scala 33:37]
  wire  _T_764; // @[Lookup.scala 33:37]
  wire  _T_765; // @[Lookup.scala 33:37]
  wire  _T_766; // @[Lookup.scala 33:37]
  wire  _T_767; // @[Lookup.scala 33:37]
  wire  _T_768; // @[Lookup.scala 33:37]
  wire  _T_769; // @[Lookup.scala 33:37]
  wire  _T_770; // @[Lookup.scala 33:37]
  wire  _T_771; // @[Lookup.scala 33:37]
  wire  _T_772; // @[Lookup.scala 33:37]
  wire  _T_773; // @[Lookup.scala 33:37]
  wire  _T_774; // @[Lookup.scala 33:37]
  wire  _T_775; // @[Lookup.scala 33:37]
  wire  _T_776; // @[Lookup.scala 33:37]
  wire  _T_777; // @[Lookup.scala 33:37]
  wire  _T_778; // @[Lookup.scala 33:37]
  wire  _T_779; // @[Lookup.scala 33:37]
  wire  _T_780; // @[Lookup.scala 33:37]
  wire  _T_781; // @[Lookup.scala 33:37]
  wire  _T_782; // @[Lookup.scala 33:37]
  wire  _T_783; // @[Lookup.scala 33:37]
  wire  _T_784; // @[Lookup.scala 33:37]
  wire  _T_785; // @[Lookup.scala 33:37]
  wire  _T_786; // @[Lookup.scala 33:37]
  wire  _T_787; // @[Lookup.scala 33:37]
  wire  _T_788; // @[Lookup.scala 33:37]
  wire  _T_789; // @[Lookup.scala 33:37]
  wire  _T_790; // @[Lookup.scala 33:37]
  wire  _T_791; // @[Lookup.scala 33:37]
  wire  _T_792; // @[Lookup.scala 33:37]
  wire  _T_793; // @[Lookup.scala 33:37]
  wire  _T_794; // @[Lookup.scala 33:37]
  wire  _T_795; // @[Lookup.scala 33:37]
  wire  _T_796; // @[Lookup.scala 33:37]
  wire  _T_797; // @[Lookup.scala 33:37]
  wire  _T_798; // @[Lookup.scala 33:37]
  wire  _T_799; // @[Lookup.scala 33:37]
  wire  _T_800; // @[Lookup.scala 33:37]
  wire  _T_801; // @[Lookup.scala 33:37]
  wire  _T_802; // @[Lookup.scala 33:37]
  wire  _T_803; // @[Lookup.scala 33:37]
  wire  _T_804; // @[Lookup.scala 33:37]
  wire  _T_805; // @[Lookup.scala 33:37]
  wire  _T_806; // @[Lookup.scala 33:37]
  wire  _T_807; // @[Lookup.scala 33:37]
  wire  _T_808; // @[Lookup.scala 33:37]
  wire  _T_809; // @[Lookup.scala 33:37]
  wire  _T_810; // @[Lookup.scala 33:37]
  wire  _T_811; // @[Lookup.scala 33:37]
  wire  _T_812; // @[Lookup.scala 33:37]
  wire  _T_813; // @[Lookup.scala 33:37]
  wire  _T_814; // @[Lookup.scala 33:37]
  wire  _T_815; // @[Lookup.scala 33:37]
  wire  _T_816; // @[Lookup.scala 33:37]
  wire  _T_817; // @[Lookup.scala 33:37]
  wire  _T_818; // @[Lookup.scala 33:37]
  wire  _T_819; // @[Lookup.scala 33:37]
  wire  _T_820; // @[Lookup.scala 33:37]
  wire  _T_821; // @[Lookup.scala 33:37]
  wire  _T_822; // @[Lookup.scala 33:37]
  wire  _T_823; // @[Lookup.scala 33:37]
  wire  _T_824; // @[Lookup.scala 33:37]
  wire  _T_825; // @[Lookup.scala 33:37]
  wire  _T_826; // @[Lookup.scala 33:37]
  wire  _T_827; // @[Lookup.scala 33:37]
  wire  _T_828; // @[Lookup.scala 33:37]
  wire  _T_829; // @[Lookup.scala 33:37]
  wire  _T_830; // @[Lookup.scala 33:37]
  wire  _T_831; // @[Lookup.scala 33:37]
  wire  _T_832; // @[Lookup.scala 33:37]
  wire  _T_833; // @[Lookup.scala 33:37]
  wire  _T_834; // @[Lookup.scala 33:37]
  wire  _T_835; // @[Lookup.scala 33:37]
  wire  _T_836; // @[Lookup.scala 33:37]
  wire  _T_837; // @[Lookup.scala 33:37]
  wire  _T_838; // @[Lookup.scala 33:37]
  wire  _T_839; // @[Lookup.scala 33:37]
  wire  _T_840; // @[Lookup.scala 33:37]
  wire  _T_841; // @[Lookup.scala 33:37]
  wire  _T_842; // @[Lookup.scala 33:37]
  wire  _T_843; // @[Lookup.scala 33:37]
  wire  _T_844; // @[Lookup.scala 33:37]
  wire  _T_845; // @[Lookup.scala 33:37]
  wire  _T_846; // @[Lookup.scala 33:37]
  wire  _T_847; // @[Lookup.scala 33:37]
  wire  _T_848; // @[Lookup.scala 33:37]
  wire  _T_849; // @[Lookup.scala 33:37]
  wire  _T_850; // @[Lookup.scala 33:37]
  wire  _T_851; // @[Lookup.scala 33:37]
  wire  _T_852; // @[Lookup.scala 33:37]
  wire  _T_853; // @[Lookup.scala 33:37]
  wire  _T_854; // @[Lookup.scala 33:37]
  wire  _T_855; // @[Lookup.scala 33:37]
  wire  _T_856; // @[Lookup.scala 33:37]
  wire  _T_857; // @[Lookup.scala 33:37]
  wire  _T_858; // @[Lookup.scala 33:37]
  wire  _T_859; // @[Lookup.scala 33:37]
  wire  _T_860; // @[Lookup.scala 33:37]
  wire  _T_861; // @[Lookup.scala 33:37]
  wire  _T_862; // @[Lookup.scala 33:37]
  wire  _T_863; // @[Lookup.scala 33:37]
  wire  _T_864; // @[Lookup.scala 33:37]
  wire  _T_865; // @[Lookup.scala 33:37]
  wire  _T_866; // @[Lookup.scala 33:37]
  wire  _T_867; // @[Lookup.scala 33:37]
  wire  _T_868; // @[Lookup.scala 33:37]
  wire  _T_869; // @[Lookup.scala 33:37]
  wire  _T_870; // @[Lookup.scala 33:37]
  wire  _T_871; // @[Lookup.scala 33:37]
  wire  _T_872; // @[Lookup.scala 33:37]
  wire  _T_873; // @[Lookup.scala 33:37]
  wire  _T_874; // @[Lookup.scala 33:37]
  wire  _T_875; // @[Lookup.scala 33:37]
  wire  _T_876; // @[Lookup.scala 33:37]
  wire  _T_877; // @[Lookup.scala 33:37]
  wire  _T_878; // @[Lookup.scala 33:37]
  wire  _T_879; // @[Lookup.scala 33:37]
  wire  _T_880; // @[Lookup.scala 33:37]
  wire  _T_881; // @[Lookup.scala 33:37]
  wire  _T_882; // @[Lookup.scala 33:37]
  wire  _T_883; // @[Lookup.scala 33:37]
  wire  _T_884; // @[Lookup.scala 33:37]
  wire  _T_885; // @[Lookup.scala 33:37]
  wire  _T_886; // @[Lookup.scala 33:37]
  wire  _T_887; // @[Lookup.scala 33:37]
  wire  _T_888; // @[Lookup.scala 33:37]
  wire  _T_889; // @[Lookup.scala 33:37]
  wire  _T_890; // @[Lookup.scala 33:37]
  wire  _T_891; // @[Lookup.scala 33:37]
  wire  _T_892; // @[Lookup.scala 33:37]
  wire  _T_893; // @[Lookup.scala 33:37]
  wire  _T_894; // @[Lookup.scala 33:37]
  wire  _T_895; // @[Lookup.scala 33:37]
  wire  _T_896; // @[Lookup.scala 33:37]
  wire  _T_897; // @[Lookup.scala 33:37]
  wire  _T_898; // @[Lookup.scala 33:37]
  wire  _T_899; // @[Lookup.scala 33:37]
  wire  _T_900; // @[Lookup.scala 33:37]
  wire  _T_901; // @[Lookup.scala 33:37]
  wire  _T_902; // @[Lookup.scala 33:37]
  wire  _T_903; // @[Lookup.scala 33:37]
  wire  _T_904; // @[Lookup.scala 33:37]
  wire  _T_905; // @[Lookup.scala 33:37]
  wire  _T_906; // @[Lookup.scala 33:37]
  wire  _T_907; // @[Lookup.scala 33:37]
  wire  _T_908; // @[Lookup.scala 33:37]
  wire  _T_909; // @[Lookup.scala 33:37]
  wire  _T_910; // @[Lookup.scala 33:37]
  wire  _T_911; // @[Lookup.scala 33:37]
  wire  _T_912; // @[Lookup.scala 33:37]
  wire  _T_913; // @[Lookup.scala 33:37]
  wire  _T_914; // @[Lookup.scala 33:37]
  wire  _T_915; // @[Lookup.scala 33:37]
  wire  _T_916; // @[Lookup.scala 33:37]
  wire  _T_917; // @[Lookup.scala 33:37]
  wire  _T_918; // @[Lookup.scala 33:37]
  wire  _T_919; // @[Lookup.scala 33:37]
  wire  _T_920; // @[Lookup.scala 33:37]
  wire  _T_921; // @[Lookup.scala 33:37]
  wire  _T_922; // @[Lookup.scala 33:37]
  wire  _T_923; // @[Lookup.scala 33:37]
  wire  _T_924; // @[Lookup.scala 33:37]
  wire  _T_925; // @[Lookup.scala 33:37]
  wire  _T_926; // @[Lookup.scala 33:37]
  wire  _T_927; // @[Lookup.scala 33:37]
  wire  _T_928; // @[Lookup.scala 33:37]
  wire  _T_929; // @[Lookup.scala 33:37]
  wire  _T_930; // @[Lookup.scala 33:37]
  wire  _T_931; // @[Lookup.scala 33:37]
  wire  _T_932; // @[Lookup.scala 33:37]
  wire  _T_933; // @[Lookup.scala 33:37]
  wire  _T_934; // @[Lookup.scala 33:37]
  wire  _T_935; // @[Lookup.scala 33:37]
  wire  _T_936; // @[Lookup.scala 33:37]
  wire  _T_937; // @[Lookup.scala 33:37]
  wire  _T_938; // @[Lookup.scala 33:37]
  wire  _T_939; // @[Lookup.scala 33:37]
  wire  _T_940; // @[Lookup.scala 33:37]
  wire  _T_941; // @[Lookup.scala 33:37]
  wire  _T_942; // @[Lookup.scala 33:37]
  wire  _T_943; // @[Lookup.scala 33:37]
  wire  _T_944; // @[Lookup.scala 33:37]
  wire  _T_1037; // @[Lookup.scala 33:37]
  wire  _T_1038; // @[Lookup.scala 33:37]
  wire  _T_1039; // @[Lookup.scala 33:37]
  wire  _T_1040; // @[Lookup.scala 33:37]
  wire  _T_1041; // @[Lookup.scala 33:37]
  wire  _T_1042; // @[Lookup.scala 33:37]
  wire  _T_1043; // @[Lookup.scala 33:37]
  wire  _T_1044; // @[Lookup.scala 33:37]
  wire  _T_1045; // @[Lookup.scala 33:37]
  wire  _T_1046; // @[Lookup.scala 33:37]
  wire  _T_1047; // @[Lookup.scala 33:37]
  wire  _T_1048; // @[Lookup.scala 33:37]
  wire  _T_1049; // @[Lookup.scala 33:37]
  wire  _T_1050; // @[Lookup.scala 33:37]
  wire  _T_1051; // @[Lookup.scala 33:37]
  wire  _T_1052; // @[Lookup.scala 33:37]
  wire  _T_1053; // @[Lookup.scala 33:37]
  wire  _T_1054; // @[Lookup.scala 33:37]
  wire  _T_1055; // @[Lookup.scala 33:37]
  wire  _T_1056; // @[Lookup.scala 33:37]
  wire  _T_1057; // @[Lookup.scala 33:37]
  wire  _T_1058; // @[Lookup.scala 33:37]
  wire  _T_1059; // @[Lookup.scala 33:37]
  wire  _T_1060; // @[Lookup.scala 33:37]
  wire  _T_1061; // @[Lookup.scala 33:37]
  wire  _T_1062; // @[Lookup.scala 33:37]
  wire  _T_1063; // @[Lookup.scala 33:37]
  wire  _T_1064; // @[Lookup.scala 33:37]
  wire  _T_1065; // @[Lookup.scala 33:37]
  wire  _T_1066; // @[Lookup.scala 33:37]
  wire  _T_1067; // @[Lookup.scala 33:37]
  wire  _T_1068; // @[Lookup.scala 33:37]
  wire  _T_1069; // @[Lookup.scala 33:37]
  wire  _T_1070; // @[Lookup.scala 33:37]
  wire  _T_1071; // @[Lookup.scala 33:37]
  wire  _T_1072; // @[Lookup.scala 33:37]
  wire  _T_1073; // @[Lookup.scala 33:37]
  wire  _T_1074; // @[Lookup.scala 33:37]
  wire  _T_1075; // @[Lookup.scala 33:37]
  wire  _T_1076; // @[Lookup.scala 33:37]
  wire  _T_1077; // @[Lookup.scala 33:37]
  wire  _T_1078; // @[Lookup.scala 33:37]
  wire  _T_1079; // @[Lookup.scala 33:37]
  wire  _T_1080; // @[Lookup.scala 33:37]
  wire  _T_1081; // @[Lookup.scala 33:37]
  wire  _T_1082; // @[Lookup.scala 33:37]
  wire  _T_1083; // @[Lookup.scala 33:37]
  wire  _T_1084; // @[Lookup.scala 33:37]
  wire  _T_1085; // @[Lookup.scala 33:37]
  wire  _T_1086; // @[Lookup.scala 33:37]
  wire  _T_1087; // @[Lookup.scala 33:37]
  wire  _T_1088; // @[Lookup.scala 33:37]
  wire  _T_1089; // @[Lookup.scala 33:37]
  wire  _T_1090; // @[Lookup.scala 33:37]
  wire  _T_1091; // @[Lookup.scala 33:37]
  wire  _T_1092; // @[Lookup.scala 33:37]
  wire  _T_1093; // @[Lookup.scala 33:37]
  wire  _T_1094; // @[Lookup.scala 33:37]
  wire  _T_1095; // @[Lookup.scala 33:37]
  wire  _T_1096; // @[Lookup.scala 33:37]
  wire  _T_1097; // @[Lookup.scala 33:37]
  wire  _T_1098; // @[Lookup.scala 33:37]
  wire  _T_1099; // @[Lookup.scala 33:37]
  wire  _T_1100; // @[Lookup.scala 33:37]
  wire  _T_1101; // @[Lookup.scala 33:37]
  wire  _T_1102; // @[Lookup.scala 33:37]
  wire  _T_1103; // @[Lookup.scala 33:37]
  wire  _T_1104; // @[Lookup.scala 33:37]
  wire  _T_1105; // @[Lookup.scala 33:37]
  wire  _T_1106; // @[Lookup.scala 33:37]
  wire  _T_1107; // @[Lookup.scala 33:37]
  wire  _T_1108; // @[Lookup.scala 33:37]
  wire  _T_1109; // @[Lookup.scala 33:37]
  wire  _T_1110; // @[Lookup.scala 33:37]
  wire  _T_1111; // @[Lookup.scala 33:37]
  wire  _T_1112; // @[Lookup.scala 33:37]
  wire  _T_1113; // @[Lookup.scala 33:37]
  wire  _T_1114; // @[Lookup.scala 33:37]
  wire  _T_1115; // @[Lookup.scala 33:37]
  wire  _T_1116; // @[Lookup.scala 33:37]
  wire  _T_1117; // @[Lookup.scala 33:37]
  wire  _T_1118; // @[Lookup.scala 33:37]
  wire  _T_1119; // @[Lookup.scala 33:37]
  wire  _T_1120; // @[Lookup.scala 33:37]
  wire  _T_1121; // @[Lookup.scala 33:37]
  wire  _T_1122; // @[Lookup.scala 33:37]
  wire  _T_1123; // @[Lookup.scala 33:37]
  wire  _T_1124; // @[Lookup.scala 33:37]
  wire  _T_1125; // @[Lookup.scala 33:37]
  wire  _T_1126; // @[Lookup.scala 33:37]
  wire  _T_1127; // @[Lookup.scala 33:37]
  wire  _T_1128; // @[Lookup.scala 33:37]
  wire  _T_1129; // @[Lookup.scala 33:37]
  wire  _T_1130; // @[Lookup.scala 33:37]
  wire  _T_1131; // @[Lookup.scala 33:37]
  wire  _T_1132; // @[Lookup.scala 33:37]
  wire  _T_1133; // @[Lookup.scala 33:37]
  wire  _T_1134; // @[Lookup.scala 33:37]
  wire  _T_1215; // @[Lookup.scala 33:37]
  wire  _T_1216; // @[Lookup.scala 33:37]
  wire  _T_1217; // @[Lookup.scala 33:37]
  wire  _T_1218; // @[Lookup.scala 33:37]
  wire  _T_1219; // @[Lookup.scala 33:37]
  wire  _T_1220; // @[Lookup.scala 33:37]
  wire  _T_1221; // @[Lookup.scala 33:37]
  wire  _T_1222; // @[Lookup.scala 33:37]
  wire  _T_1223; // @[Lookup.scala 33:37]
  wire  _T_1224; // @[Lookup.scala 33:37]
  wire  _T_1225; // @[Lookup.scala 33:37]
  wire  _T_1226; // @[Lookup.scala 33:37]
  wire  _T_1227; // @[Lookup.scala 33:37]
  wire  _T_1228; // @[Lookup.scala 33:37]
  wire  _T_1229; // @[Lookup.scala 33:37]
  wire  _T_1230; // @[Lookup.scala 33:37]
  wire  _T_1231; // @[Lookup.scala 33:37]
  wire  _T_1232; // @[Lookup.scala 33:37]
  wire  _T_1233; // @[Lookup.scala 33:37]
  wire  _T_1234; // @[Lookup.scala 33:37]
  wire  _T_1235; // @[Lookup.scala 33:37]
  wire  _T_1236; // @[Lookup.scala 33:37]
  wire  _T_1237; // @[Lookup.scala 33:37]
  wire  _T_1238; // @[Lookup.scala 33:37]
  wire  _T_1239; // @[Lookup.scala 33:37]
  wire  _T_1240; // @[Lookup.scala 33:37]
  wire  _T_1241; // @[Lookup.scala 33:37]
  wire  _T_1242; // @[Lookup.scala 33:37]
  wire  _T_1243; // @[Lookup.scala 33:37]
  wire  _T_1244; // @[Lookup.scala 33:37]
  wire  _T_1245; // @[Lookup.scala 33:37]
  wire  _T_1246; // @[Lookup.scala 33:37]
  wire  _T_1247; // @[Lookup.scala 33:37]
  wire  _T_1248; // @[Lookup.scala 33:37]
  wire  _T_1249; // @[Lookup.scala 33:37]
  wire  _T_1250; // @[Lookup.scala 33:37]
  wire  _T_1251; // @[Lookup.scala 33:37]
  wire  _T_1252; // @[Lookup.scala 33:37]
  wire  _T_1253; // @[Lookup.scala 33:37]
  wire  _T_1254; // @[Lookup.scala 33:37]
  wire  _T_1255; // @[Lookup.scala 33:37]
  wire  _T_1256; // @[Lookup.scala 33:37]
  wire  _T_1257; // @[Lookup.scala 33:37]
  wire  _T_1258; // @[Lookup.scala 33:37]
  wire  _T_1259; // @[Lookup.scala 33:37]
  wire  _T_1260; // @[Lookup.scala 33:37]
  wire  _T_1261; // @[Lookup.scala 33:37]
  wire  _T_1262; // @[Lookup.scala 33:37]
  wire  _T_1263; // @[Lookup.scala 33:37]
  wire  _T_1264; // @[Lookup.scala 33:37]
  wire  _T_1265; // @[Lookup.scala 33:37]
  wire  _T_1266; // @[Lookup.scala 33:37]
  wire  _T_1267; // @[Lookup.scala 33:37]
  wire  _T_1268; // @[Lookup.scala 33:37]
  wire  _T_1269; // @[Lookup.scala 33:37]
  wire  _T_1270; // @[Lookup.scala 33:37]
  wire  _T_1271; // @[Lookup.scala 33:37]
  wire  _T_1272; // @[Lookup.scala 33:37]
  wire  _T_1273; // @[Lookup.scala 33:37]
  wire  _T_1274; // @[Lookup.scala 33:37]
  wire  _T_1275; // @[Lookup.scala 33:37]
  wire  _T_1276; // @[Lookup.scala 33:37]
  wire  _T_1277; // @[Lookup.scala 33:37]
  wire  _T_1278; // @[Lookup.scala 33:37]
  wire  _T_1279; // @[Lookup.scala 33:37]
  wire  _T_1280; // @[Lookup.scala 33:37]
  wire  _T_1281; // @[Lookup.scala 33:37]
  wire  _T_1282; // @[Lookup.scala 33:37]
  wire  _T_1283; // @[Lookup.scala 33:37]
  wire  _T_1284; // @[Lookup.scala 33:37]
  wire  _T_1285; // @[Lookup.scala 33:37]
  wire  _T_1286; // @[Lookup.scala 33:37]
  wire  _T_1287; // @[Lookup.scala 33:37]
  wire  _T_1288; // @[Lookup.scala 33:37]
  wire  _T_1289; // @[Lookup.scala 33:37]
  wire  _T_1290; // @[Lookup.scala 33:37]
  wire  _T_1291; // @[Lookup.scala 33:37]
  wire  _T_1292; // @[Lookup.scala 33:37]
  wire  _T_1293; // @[Lookup.scala 33:37]
  wire  _T_1294; // @[Lookup.scala 33:37]
  wire  _T_1295; // @[Lookup.scala 33:37]
  wire  _T_1296; // @[Lookup.scala 33:37]
  wire  _T_1297; // @[Lookup.scala 33:37]
  wire  _T_1298; // @[Lookup.scala 33:37]
  wire  _T_1299; // @[Lookup.scala 33:37]
  wire  _T_1300; // @[Lookup.scala 33:37]
  wire  _T_1301; // @[Lookup.scala 33:37]
  wire  _T_1302; // @[Lookup.scala 33:37]
  wire  _T_1303; // @[Lookup.scala 33:37]
  wire  _T_1304; // @[Lookup.scala 33:37]
  wire  _T_1305; // @[Lookup.scala 33:37]
  wire  _T_1306; // @[Lookup.scala 33:37]
  wire  _T_1307; // @[Lookup.scala 33:37]
  wire  _T_1308; // @[Lookup.scala 33:37]
  wire  _T_1309; // @[Lookup.scala 33:37]
  wire  _T_1310; // @[Lookup.scala 33:37]
  wire  _T_1311; // @[Lookup.scala 33:37]
  wire  _T_1312; // @[Lookup.scala 33:37]
  wire  _T_1313; // @[Lookup.scala 33:37]
  wire  _T_1314; // @[Lookup.scala 33:37]
  wire  _T_1315; // @[Lookup.scala 33:37]
  wire  _T_1316; // @[Lookup.scala 33:37]
  wire  _T_1317; // @[Lookup.scala 33:37]
  wire  _T_1318; // @[Lookup.scala 33:37]
  wire  _T_1319; // @[Lookup.scala 33:37]
  wire  _T_1320; // @[Lookup.scala 33:37]
  wire  _T_1321; // @[Lookup.scala 33:37]
  wire  _T_1322; // @[Lookup.scala 33:37]
  wire  _T_1434; // @[Lookup.scala 33:37]
  wire  _T_1435; // @[Lookup.scala 33:37]
  wire  _T_1436; // @[Lookup.scala 33:37]
  wire  _T_1437; // @[Lookup.scala 33:37]
  wire  _T_1438; // @[Lookup.scala 33:37]
  wire  _T_1439; // @[Lookup.scala 33:37]
  wire  _T_1440; // @[Lookup.scala 33:37]
  wire  _T_1441; // @[Lookup.scala 33:37]
  wire  _T_1442; // @[Lookup.scala 33:37]
  wire  _T_1443; // @[Lookup.scala 33:37]
  wire  _T_1444; // @[Lookup.scala 33:37]
  wire  _T_1445; // @[Lookup.scala 33:37]
  wire  _T_1446; // @[Lookup.scala 33:37]
  wire  _T_1447; // @[Lookup.scala 33:37]
  wire  _T_1448; // @[Lookup.scala 33:37]
  wire  _T_1449; // @[Lookup.scala 33:37]
  wire  _T_1450; // @[Lookup.scala 33:37]
  wire  _T_1451; // @[Lookup.scala 33:37]
  wire  _T_1452; // @[Lookup.scala 33:37]
  wire  _T_1453; // @[Lookup.scala 33:37]
  wire  _T_1454; // @[Lookup.scala 33:37]
  wire  _T_1455; // @[Lookup.scala 33:37]
  wire  _T_1456; // @[Lookup.scala 33:37]
  wire  _T_1457; // @[Lookup.scala 33:37]
  wire  _T_1458; // @[Lookup.scala 33:37]
  wire  _T_1459; // @[Lookup.scala 33:37]
  wire  _T_1460; // @[Lookup.scala 33:37]
  wire  _T_1461; // @[Lookup.scala 33:37]
  wire  _T_1462; // @[Lookup.scala 33:37]
  wire  _T_1463; // @[Lookup.scala 33:37]
  wire  _T_1464; // @[Lookup.scala 33:37]
  wire  _T_1465; // @[Lookup.scala 33:37]
  wire  _T_1466; // @[Lookup.scala 33:37]
  wire  _T_1467; // @[Lookup.scala 33:37]
  wire  _T_1468; // @[Lookup.scala 33:37]
  wire  _T_1469; // @[Lookup.scala 33:37]
  wire  _T_1470; // @[Lookup.scala 33:37]
  wire  _T_1471; // @[Lookup.scala 33:37]
  wire  _T_1472; // @[Lookup.scala 33:37]
  wire  _T_1473; // @[Lookup.scala 33:37]
  wire  _T_1474; // @[Lookup.scala 33:37]
  wire  _T_1475; // @[Lookup.scala 33:37]
  wire  _T_1476; // @[Lookup.scala 33:37]
  wire  _T_1477; // @[Lookup.scala 33:37]
  wire  _T_1478; // @[Lookup.scala 33:37]
  wire  _T_1479; // @[Lookup.scala 33:37]
  wire  _T_1480; // @[Lookup.scala 33:37]
  wire  _T_1481; // @[Lookup.scala 33:37]
  wire  _T_1482; // @[Lookup.scala 33:37]
  wire  _T_1483; // @[Lookup.scala 33:37]
  wire  _T_1484; // @[Lookup.scala 33:37]
  wire  _T_1485; // @[Lookup.scala 33:37]
  wire  _T_1486; // @[Lookup.scala 33:37]
  wire  _T_1487; // @[Lookup.scala 33:37]
  wire  _T_1488; // @[Lookup.scala 33:37]
  wire  _T_1489; // @[Lookup.scala 33:37]
  wire  _T_1490; // @[Lookup.scala 33:37]
  wire  _T_1491; // @[Lookup.scala 33:37]
  wire  _T_1492; // @[Lookup.scala 33:37]
  wire  _T_1493; // @[Lookup.scala 33:37]
  wire  _T_1494; // @[Lookup.scala 33:37]
  wire  _T_1495; // @[Lookup.scala 33:37]
  wire  _T_1496; // @[Lookup.scala 33:37]
  wire  _T_1497; // @[Lookup.scala 33:37]
  wire  _T_1498; // @[Lookup.scala 33:37]
  wire  _T_1499; // @[Lookup.scala 33:37]
  wire  _T_1500; // @[Lookup.scala 33:37]
  wire  _T_1501; // @[Lookup.scala 33:37]
  wire  _T_1502; // @[Lookup.scala 33:37]
  wire  _T_1503; // @[Lookup.scala 33:37]
  wire  _T_1504; // @[Lookup.scala 33:37]
  wire  _T_1505; // @[Lookup.scala 33:37]
  wire  _T_1506; // @[Lookup.scala 33:37]
  wire  _T_1507; // @[Lookup.scala 33:37]
  wire  _T_1508; // @[Lookup.scala 33:37]
  wire  _T_1509; // @[Lookup.scala 33:37]
  wire  _T_1510; // @[Lookup.scala 33:37]
  wire  _T_1511; // @[Lookup.scala 33:37]
  wire  _T_1517; // @[Lookup.scala 33:37]
  wire  _T_1518; // @[Lookup.scala 33:37]
  wire  _T_1519; // @[Lookup.scala 33:37]
  wire  _T_1520; // @[Lookup.scala 33:37]
  wire  _T_1521; // @[Lookup.scala 33:37]
  wire  _T_1522; // @[Lookup.scala 33:37]
  wire  _T_1523; // @[Lookup.scala 33:37]
  wire  _T_1524; // @[Lookup.scala 33:37]
  wire  _T_1525; // @[Lookup.scala 33:37]
  wire  _T_1526; // @[Lookup.scala 33:37]
  wire  _T_1527; // @[Lookup.scala 33:37]
  wire  _T_1528; // @[Lookup.scala 33:37]
  wire  _T_1529; // @[Lookup.scala 33:37]
  wire  _T_1530; // @[Lookup.scala 33:37]
  wire  _T_1531; // @[Lookup.scala 33:37]
  wire  _T_1532; // @[Lookup.scala 33:37]
  wire  _T_1533; // @[Lookup.scala 33:37]
  wire  _T_1534; // @[Lookup.scala 33:37]
  wire  _T_1535; // @[Lookup.scala 33:37]
  wire  _T_1536; // @[Lookup.scala 33:37]
  wire  _T_1537; // @[Lookup.scala 33:37]
  wire  _T_1538; // @[Lookup.scala 33:37]
  wire  _T_1539; // @[Lookup.scala 33:37]
  wire  _T_1540; // @[Lookup.scala 33:37]
  wire  _T_1541; // @[Lookup.scala 33:37]
  wire  _T_1542; // @[Lookup.scala 33:37]
  wire  _T_1543; // @[Lookup.scala 33:37]
  wire  _T_1544; // @[Lookup.scala 33:37]
  wire  _T_1545; // @[Lookup.scala 33:37]
  wire  _T_1546; // @[Lookup.scala 33:37]
  wire  _T_1547; // @[Lookup.scala 33:37]
  wire  _T_1548; // @[Lookup.scala 33:37]
  wire  _T_1549; // @[Lookup.scala 33:37]
  wire  _T_1550; // @[Lookup.scala 33:37]
  wire  _T_1551; // @[Lookup.scala 33:37]
  wire  _T_1552; // @[Lookup.scala 33:37]
  wire  _T_1553; // @[Lookup.scala 33:37]
  wire  _T_1554; // @[Lookup.scala 33:37]
  wire  _T_1555; // @[Lookup.scala 33:37]
  wire  _T_1556; // @[Lookup.scala 33:37]
  wire  _T_1557; // @[Lookup.scala 33:37]
  wire  _T_1558; // @[Lookup.scala 33:37]
  wire  _T_1559; // @[Lookup.scala 33:37]
  wire  _T_1560; // @[Lookup.scala 33:37]
  wire  _T_1561; // @[Lookup.scala 33:37]
  wire  _T_1562; // @[Lookup.scala 33:37]
  wire  _T_1563; // @[Lookup.scala 33:37]
  wire  _T_1564; // @[Lookup.scala 33:37]
  wire  _T_1565; // @[Lookup.scala 33:37]
  wire  _T_1566; // @[Lookup.scala 33:37]
  wire  _T_1567; // @[Lookup.scala 33:37]
  wire  _T_1568; // @[Lookup.scala 33:37]
  wire  _T_1569; // @[Lookup.scala 33:37]
  wire  _T_1570; // @[Lookup.scala 33:37]
  wire  _T_1571; // @[Lookup.scala 33:37]
  wire  _T_1572; // @[Lookup.scala 33:37]
  wire  _T_1573; // @[Lookup.scala 33:37]
  wire  _T_1574; // @[Lookup.scala 33:37]
  wire  _T_1575; // @[Lookup.scala 33:37]
  wire  _T_1576; // @[Lookup.scala 33:37]
  wire  _T_1577; // @[Lookup.scala 33:37]
  wire  _T_1578; // @[Lookup.scala 33:37]
  wire  _T_1579; // @[Lookup.scala 33:37]
  wire  _T_1580; // @[Lookup.scala 33:37]
  wire  _T_1581; // @[Lookup.scala 33:37]
  wire  _T_1582; // @[Lookup.scala 33:37]
  wire  _T_1583; // @[Lookup.scala 33:37]
  wire  _T_1584; // @[Lookup.scala 33:37]
  wire  _T_1585; // @[Lookup.scala 33:37]
  wire  _T_1586; // @[Lookup.scala 33:37]
  wire  _T_1587; // @[Lookup.scala 33:37]
  wire  _T_1588; // @[Lookup.scala 33:37]
  wire  _T_1589; // @[Lookup.scala 33:37]
  wire  _T_1590; // @[Lookup.scala 33:37]
  wire  _T_1591; // @[Lookup.scala 33:37]
  wire  _T_1592; // @[Lookup.scala 33:37]
  wire  _T_1593; // @[Lookup.scala 33:37]
  wire  _T_1594; // @[Lookup.scala 33:37]
  wire  _T_1595; // @[Lookup.scala 33:37]
  wire  _T_1596; // @[Lookup.scala 33:37]
  wire  _T_1597; // @[Lookup.scala 33:37]
  wire  _T_1598; // @[Lookup.scala 33:37]
  wire  _T_1599; // @[Lookup.scala 33:37]
  wire  _T_1600; // @[Lookup.scala 33:37]
  wire  _T_1601; // @[Lookup.scala 33:37]
  wire  _T_1602; // @[Lookup.scala 33:37]
  wire  _T_1603; // @[Lookup.scala 33:37]
  wire  _T_1604; // @[Lookup.scala 33:37]
  wire  _T_1605; // @[Lookup.scala 33:37]
  wire  _T_1606; // @[Lookup.scala 33:37]
  wire  _T_1607; // @[Lookup.scala 33:37]
  wire  _T_1608; // @[Lookup.scala 33:37]
  wire  _T_1609; // @[Lookup.scala 33:37]
  wire  _T_1610; // @[Lookup.scala 33:37]
  wire  _T_1611; // @[Lookup.scala 33:37]
  wire  _T_1612; // @[Lookup.scala 33:37]
  wire  _T_1613; // @[Lookup.scala 33:37]
  wire  _T_1614; // @[Lookup.scala 33:37]
  wire  _T_1615; // @[Lookup.scala 33:37]
  wire  _T_1616; // @[Lookup.scala 33:37]
  wire  _T_1617; // @[Lookup.scala 33:37]
  wire  _T_1618; // @[Lookup.scala 33:37]
  wire  _T_1619; // @[Lookup.scala 33:37]
  wire  _T_1620; // @[Lookup.scala 33:37]
  wire  _T_1621; // @[Lookup.scala 33:37]
  wire  _T_1622; // @[Lookup.scala 33:37]
  wire  _T_1623; // @[Lookup.scala 33:37]
  wire  _T_1624; // @[Lookup.scala 33:37]
  wire  _T_1625; // @[Lookup.scala 33:37]
  wire  _T_1626; // @[Lookup.scala 33:37]
  wire  _T_1627; // @[Lookup.scala 33:37]
  wire  _T_1628; // @[Lookup.scala 33:37]
  wire  _T_1629; // @[Lookup.scala 33:37]
  wire  _T_1630; // @[Lookup.scala 33:37]
  wire  _T_1631; // @[Lookup.scala 33:37]
  wire  _T_1632; // @[Lookup.scala 33:37]
  wire  _T_1633; // @[Lookup.scala 33:37]
  wire  _T_1634; // @[Lookup.scala 33:37]
  wire  _T_1635; // @[Lookup.scala 33:37]
  wire  _T_1636; // @[Lookup.scala 33:37]
  wire  _T_1637; // @[Lookup.scala 33:37]
  wire  _T_1638; // @[Lookup.scala 33:37]
  wire  _T_1639; // @[Lookup.scala 33:37]
  wire  _T_1640; // @[Lookup.scala 33:37]
  wire  _T_1641; // @[Lookup.scala 33:37]
  wire  _T_1642; // @[Lookup.scala 33:37]
  wire  _T_1643; // @[Lookup.scala 33:37]
  wire  _T_1644; // @[Lookup.scala 33:37]
  wire  _T_1645; // @[Lookup.scala 33:37]
  wire  _T_1646; // @[Lookup.scala 33:37]
  wire  _T_1647; // @[Lookup.scala 33:37]
  wire  _T_1648; // @[Lookup.scala 33:37]
  wire  _T_1649; // @[Lookup.scala 33:37]
  wire  _T_1650; // @[Lookup.scala 33:37]
  wire  _T_1651; // @[Lookup.scala 33:37]
  wire  _T_1652; // @[Lookup.scala 33:37]
  wire  _T_1653; // @[Lookup.scala 33:37]
  wire  _T_1654; // @[Lookup.scala 33:37]
  wire  _T_1655; // @[Lookup.scala 33:37]
  wire  _T_1656; // @[Lookup.scala 33:37]
  wire  _T_1657; // @[Lookup.scala 33:37]
  wire  _T_1658; // @[Lookup.scala 33:37]
  wire  _T_1659; // @[Lookup.scala 33:37]
  wire  _T_1660; // @[Lookup.scala 33:37]
  wire  _T_1661; // @[Lookup.scala 33:37]
  wire  _T_1662; // @[Lookup.scala 33:37]
  wire  _T_1663; // @[Lookup.scala 33:37]
  wire  _T_1664; // @[Lookup.scala 33:37]
  wire  _T_1665; // @[Lookup.scala 33:37]
  wire  _T_1666; // @[Lookup.scala 33:37]
  wire  _T_1667; // @[Lookup.scala 33:37]
  wire  _T_1668; // @[Lookup.scala 33:37]
  wire  _T_1669; // @[Lookup.scala 33:37]
  wire  _T_1670; // @[Lookup.scala 33:37]
  wire  _T_1671; // @[Lookup.scala 33:37]
  wire  _T_1672; // @[Lookup.scala 33:37]
  wire  _T_1673; // @[Lookup.scala 33:37]
  wire  _T_1674; // @[Lookup.scala 33:37]
  wire  _T_1675; // @[Lookup.scala 33:37]
  wire  _T_1676; // @[Lookup.scala 33:37]
  wire  _T_1677; // @[Lookup.scala 33:37]
  wire  _T_1678; // @[Lookup.scala 33:37]
  wire  _T_1679; // @[Lookup.scala 33:37]
  wire  _T_1680; // @[Lookup.scala 33:37]
  wire  _T_1681; // @[Lookup.scala 33:37]
  wire  _T_1682; // @[Lookup.scala 33:37]
  wire  _T_1683; // @[Lookup.scala 33:37]
  wire  _T_1684; // @[Lookup.scala 33:37]
  wire  _T_1685; // @[Lookup.scala 33:37]
  wire  _T_1686; // @[Lookup.scala 33:37]
  wire  _T_1687; // @[Lookup.scala 33:37]
  wire  _T_1688; // @[Lookup.scala 33:37]
  wire  _T_1689; // @[Lookup.scala 33:37]
  wire  _T_1690; // @[Lookup.scala 33:37]
  wire  _T_1691; // @[Lookup.scala 33:37]
  wire  _T_1692; // @[Lookup.scala 33:37]
  wire  _T_1693; // @[Lookup.scala 33:37]
  wire  _T_1694; // @[Lookup.scala 33:37]
  wire  _T_1695; // @[Lookup.scala 33:37]
  wire  _T_1696; // @[Lookup.scala 33:37]
  wire  _T_1697; // @[Lookup.scala 33:37]
  wire  _T_1698; // @[Lookup.scala 33:37]
  wire  _T_1699; // @[Lookup.scala 33:37]
  wire  _T_1700; // @[Lookup.scala 33:37]
  wire  _T_1722; // @[Mux.scala 80:60]
  wire [4:0] _T_1723; // @[Mux.scala 80:57]
  wire  _T_1725; // @[Mux.scala 80:60]
  wire [4:0] _T_1726; // @[Mux.scala 80:57]
  wire  _T_1727; // @[Mux.scala 80:60]
  wire [4:0] _T_1728; // @[Mux.scala 80:57]
  wire  _T_1729; // @[Mux.scala 80:60]
  wire [4:0] _T_1730; // @[Mux.scala 80:57]
  wire  _T_1731; // @[Mux.scala 80:60]
  wire [4:0] _T_1732; // @[Mux.scala 80:57]
  wire  _T_1733; // @[Mux.scala 80:60]
  wire [4:0] _T_1734; // @[Mux.scala 80:57]
  wire  _T_1735; // @[Mux.scala 80:60]
  wire [4:0] _T_1736; // @[Mux.scala 80:57]
  wire  _T_1737; // @[Mux.scala 80:60]
  wire [4:0] _T_1738; // @[Mux.scala 80:57]
  wire  _T_1739; // @[Mux.scala 80:60]
  wire [4:0] _T_1740; // @[Mux.scala 80:57]
  wire  _T_1741; // @[Mux.scala 80:60]
  wire [4:0] _T_1742; // @[Mux.scala 80:57]
  wire [4:0] _T_1744; // @[Mux.scala 80:57]
  wire  _T_1745; // @[Mux.scala 80:60]
  wire [4:0] _T_1746; // @[Mux.scala 80:57]
  wire  _T_1747; // @[Mux.scala 80:60]
  wire [4:0] _T_1748; // @[Mux.scala 80:57]
  wire  _T_1749; // @[Mux.scala 80:60]
  wire [4:0] _T_1750; // @[Mux.scala 80:57]
  wire  _T_1751; // @[Mux.scala 80:60]
  wire [4:0] _T_1752; // @[Mux.scala 80:57]
  wire  _T_1753; // @[Mux.scala 80:60]
  wire [4:0] _T_1754; // @[Mux.scala 80:57]
  wire  _T_1755; // @[Mux.scala 80:60]
  wire [4:0] _T_1756; // @[Mux.scala 80:57]
  wire  _T_1757; // @[Mux.scala 80:60]
  wire [4:0] _T_1758; // @[Mux.scala 80:57]
  wire  _T_1759; // @[Mux.scala 80:60]
  wire [4:0] _T_1760; // @[Mux.scala 80:57]
  wire  _T_1761; // @[Mux.scala 80:60]
  wire  _T_1783; // @[Mux.scala 80:60]
  wire [4:0] _T_1784; // @[Mux.scala 80:57]
  wire [4:0] _T_1787; // @[Mux.scala 80:57]
  wire [4:0] _T_1789; // @[Mux.scala 80:57]
  wire [4:0] _T_1791; // @[Mux.scala 80:57]
  wire [4:0] _T_1793; // @[Mux.scala 80:57]
  wire [4:0] _T_1795; // @[Mux.scala 80:57]
  wire [4:0] _T_1797; // @[Mux.scala 80:57]
  wire [4:0] _T_1799; // @[Mux.scala 80:57]
  wire [4:0] _T_1801; // @[Mux.scala 80:57]
  wire  _T_1802; // @[Mux.scala 80:60]
  wire [4:0] _T_1803; // @[Mux.scala 80:57]
  wire  _T_1804; // @[Mux.scala 80:60]
  wire [4:0] _T_1805; // @[Mux.scala 80:57]
  wire [4:0] _T_1807; // @[Mux.scala 80:57]
  wire [4:0] _T_1809; // @[Mux.scala 80:57]
  wire [4:0] _T_1811; // @[Mux.scala 80:57]
  wire [4:0] _T_1813; // @[Mux.scala 80:57]
  wire [4:0] _T_1815; // @[Mux.scala 80:57]
  wire [4:0] _T_1817; // @[Mux.scala 80:57]
  wire [4:0] _T_1819; // @[Mux.scala 80:57]
  wire [4:0] _T_1821; // @[Mux.scala 80:57]
  wire [4:0] _T_1840; // @[Mux.scala 80:57]
  wire [4:0] _T_1843; // @[Mux.scala 80:57]
  wire [4:0] _T_1845; // @[Mux.scala 80:57]
  wire [4:0] _T_1847; // @[Mux.scala 80:57]
  wire  _T_1848; // @[Mux.scala 80:60]
  wire [4:0] _T_1849; // @[Mux.scala 80:57]
  wire [4:0] _T_1851; // @[Mux.scala 80:57]
  wire [4:0] _T_1853; // @[Mux.scala 80:57]
  wire [4:0] _T_1855; // @[Mux.scala 80:57]
  wire [4:0] _T_1857; // @[Mux.scala 80:57]
  wire  _T_1858; // @[Mux.scala 80:60]
  wire [4:0] _T_1859; // @[Mux.scala 80:57]
  wire [4:0] _T_1861; // @[Mux.scala 80:57]
  wire [4:0] _T_1863; // @[Mux.scala 80:57]
  wire [4:0] _T_1865; // @[Mux.scala 80:57]
  wire [4:0] _T_1867; // @[Mux.scala 80:57]
  wire [20:0] _T_1879; // @[Cat.scala 29:58]
  wire [12:0] _T_1891; // @[Mux.scala 80:57]
  wire [12:0] _T_1894; // @[Mux.scala 80:57]
  wire [17:0] _T_1896; // @[Mux.scala 80:57]
  wire [18:0] _T_1898; // @[Mux.scala 80:57]
  wire [18:0] _T_1900; // @[Mux.scala 80:57]
  wire [18:0] _T_1902; // @[Mux.scala 80:57]
  wire  _T_1903; // @[Mux.scala 80:60]
  wire [25:0] _T_1904; // @[Mux.scala 80:57]
  wire [25:0] _T_1906; // @[Mux.scala 80:57]
  wire  _T_1907; // @[Mux.scala 80:60]
  wire [25:0] _T_1908; // @[Mux.scala 80:57]
  wire [25:0] _T_1910; // @[Mux.scala 80:57]
  wire [25:0] _T_1912; // @[Mux.scala 80:57]
  wire [25:0] _T_1914; // @[Mux.scala 80:57]
  wire [25:0] _T_1916; // @[Mux.scala 80:57]
  wire [25:0] _T_1918; // @[Mux.scala 80:57]
  wire [25:0] _T_1920; // @[Mux.scala 80:57]
  wire [25:0] _T_1922; // @[Mux.scala 80:57]
  wire [25:0] _T_1924; // @[Mux.scala 80:57]
  wire [3:0] _T_1930; // @[Decode.scala 131:21]
  wire [5:0] _T_1933; // @[Mux.scala 80:57]
  wire [5:0] _T_1936; // @[Mux.scala 80:57]
  wire [5:0] _T_1938; // @[Mux.scala 80:57]
  wire [5:0] _T_1940; // @[Mux.scala 80:57]
  wire [1:0] _T_1945; // @[Mux.scala 80:57]
  wire [1:0] _T_1948; // @[Mux.scala 80:57]
  wire [1:0] _T_1950; // @[Mux.scala 80:57]
  wire [1:0] _T_1952; // @[Mux.scala 80:57]
  wire [3:0] _T_1960; // @[Mux.scala 80:57]
  wire [3:0] _T_1963; // @[Mux.scala 80:57]
  wire [3:0] _T_1965; // @[Mux.scala 80:57]
  wire [3:0] _T_1971; // @[Mux.scala 80:57]
  wire  _T_1976; // @[Decode.scala 164:16]
  assign _T_1 = io_finst_inst & 32'h9f000000; // @[Lookup.scala 31:38]
  assign _T_2 = 32'h10000000 == _T_1; // @[Lookup.scala 31:38]
  assign _T_4 = 32'h90000000 == _T_1; // @[Lookup.scala 31:38]
  assign _T_5 = io_finst_inst & 32'hff20001f; // @[Lookup.scala 31:38]
  assign _T_6 = 32'h6a00001f == _T_5; // @[Lookup.scala 31:38]
  assign _T_7 = io_finst_inst & 32'hff200000; // @[Lookup.scala 31:38]
  assign _T_8 = 32'ha000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_10 = 32'ha200000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_12 = 32'h2a000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_14 = 32'h2a200000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_16 = 32'h4a000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_18 = 32'h4a200000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_20 = 32'h6a000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_22 = 32'h6a200000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_24 = 32'hea00001f == _T_5; // @[Lookup.scala 31:38]
  assign _T_26 = 32'h8a000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_28 = 32'h8a200000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_30 = 32'haa000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_32 = 32'haa200000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_34 = 32'hca000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_36 = 32'hca200000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_38 = 32'hea000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_40 = 32'hea200000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_41 = io_finst_inst & 32'hffc0001f; // @[Lookup.scala 31:38]
  assign _T_42 = 32'h7200001f == _T_41; // @[Lookup.scala 31:38]
  assign _T_43 = io_finst_inst & 32'hffc00000; // @[Lookup.scala 31:38]
  assign _T_44 = 32'h12000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_46 = 32'h32000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_48 = 32'h52000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_50 = 32'h72000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_51 = io_finst_inst & 32'hff80001f; // @[Lookup.scala 31:38]
  assign _T_52 = 32'hf200001f == _T_51; // @[Lookup.scala 31:38]
  assign _T_53 = io_finst_inst & 32'hff800000; // @[Lookup.scala 31:38]
  assign _T_54 = 32'h92000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_56 = 32'hb2000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_58 = 32'hd2000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_60 = 32'hf2000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_62 = 32'h12800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_64 = 32'h52800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_66 = 32'h72800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_68 = 32'h92800000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_70 = 32'hd2800000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_72 = 32'hf2800000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_74 = 32'h13000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_76 = 32'h33000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_78 = 32'h53000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_80 = 32'h93400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_82 = 32'hb3400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_84 = 32'hd3400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_85 = io_finst_inst & 32'hffe00c00; // @[Lookup.scala 31:38]
  assign _T_86 = 32'h1a800000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_88 = 32'h1a800400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_90 = 32'h5a800000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_92 = 32'h5a800400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_94 = 32'h9a800000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_96 = 32'h9a800400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_98 = 32'hda800000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_100 = 32'hda800400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_101 = io_finst_inst & 32'hffe00c10; // @[Lookup.scala 31:38]
  assign _T_102 = 32'hba400800 == _T_101; // @[Lookup.scala 31:38]
  assign _T_104 = 32'hfa400800 == _T_101; // @[Lookup.scala 31:38]
  assign _T_106 = 32'h7a400800 == _T_101; // @[Lookup.scala 31:38]
  assign _T_108 = 32'hba400000 == _T_101; // @[Lookup.scala 31:38]
  assign _T_110 = 32'hfa400000 == _T_101; // @[Lookup.scala 31:38]
  assign _T_112 = 32'h7a400000 == _T_101; // @[Lookup.scala 31:38]
  assign _T_114 = 32'h6b00001f == _T_5; // @[Lookup.scala 31:38]
  assign _T_116 = 32'h2b00001f == _T_5; // @[Lookup.scala 31:38]
  assign _T_118 = 32'hb000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_120 = 32'h2b000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_122 = 32'h4b000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_124 = 32'h6b000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_126 = 32'heb00001f == _T_5; // @[Lookup.scala 31:38]
  assign _T_128 = 32'hab00001f == _T_5; // @[Lookup.scala 31:38]
  assign _T_130 = 32'h8b000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_132 = 32'hab000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_134 = 32'hcb000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_136 = 32'heb000000 == _T_7; // @[Lookup.scala 31:38]
  assign _T_138 = 32'h7100001f == _T_51; // @[Lookup.scala 31:38]
  assign _T_140 = 32'h3100001f == _T_51; // @[Lookup.scala 31:38]
  assign _T_142 = 32'h11000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_144 = 32'h31000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_146 = 32'h51000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_148 = 32'h71000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_150 = 32'hf100001f == _T_51; // @[Lookup.scala 31:38]
  assign _T_152 = 32'hb100001f == _T_51; // @[Lookup.scala 31:38]
  assign _T_154 = 32'h91000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_156 = 32'hb1000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_158 = 32'hd1000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_160 = 32'hf1000000 == _T_53; // @[Lookup.scala 31:38]
  assign _T_161 = io_finst_inst & 32'hfffffc00; // @[Lookup.scala 31:38]
  assign _T_162 = 32'h5ac00000 == _T_161; // @[Lookup.scala 31:38]
  assign _T_164 = 32'h5ac00400 == _T_161; // @[Lookup.scala 31:38]
  assign _T_166 = 32'h5ac00800 == _T_161; // @[Lookup.scala 31:38]
  assign _T_168 = 32'h5ac01000 == _T_161; // @[Lookup.scala 31:38]
  assign _T_170 = 32'h5ac01400 == _T_161; // @[Lookup.scala 31:38]
  assign _T_172 = 32'hdac00000 == _T_161; // @[Lookup.scala 31:38]
  assign _T_174 = 32'hdac00400 == _T_161; // @[Lookup.scala 31:38]
  assign _T_176 = 32'hdac00800 == _T_161; // @[Lookup.scala 31:38]
  assign _T_178 = 32'hdac00c00 == _T_161; // @[Lookup.scala 31:38]
  assign _T_180 = 32'hdac01000 == _T_161; // @[Lookup.scala 31:38]
  assign _T_182 = 32'hdac01400 == _T_161; // @[Lookup.scala 31:38]
  assign _T_183 = io_finst_inst & 32'hffe0fc00; // @[Lookup.scala 31:38]
  assign _T_184 = 32'h1ac02000 == _T_183; // @[Lookup.scala 31:38]
  assign _T_186 = 32'h1ac02400 == _T_183; // @[Lookup.scala 31:38]
  assign _T_188 = 32'h1ac02800 == _T_183; // @[Lookup.scala 31:38]
  assign _T_190 = 32'h1ac02c00 == _T_183; // @[Lookup.scala 31:38]
  assign _T_192 = 32'h9ac02000 == _T_183; // @[Lookup.scala 31:38]
  assign _T_194 = 32'h9ac02400 == _T_183; // @[Lookup.scala 31:38]
  assign _T_196 = 32'h9ac02800 == _T_183; // @[Lookup.scala 31:38]
  assign _T_198 = 32'h9ac02c00 == _T_183; // @[Lookup.scala 31:38]
  assign _T_199 = io_finst_inst & 32'hffe08000; // @[Lookup.scala 31:38]
  assign _T_200 = 32'h1b000000 == _T_199; // @[Lookup.scala 31:38]
  assign _T_201 = io_finst_inst & 32'hfc000000; // @[Lookup.scala 31:38]
  assign _T_202 = 32'h14000000 == _T_201; // @[Lookup.scala 31:38]
  assign _T_204 = 32'h94000000 == _T_201; // @[Lookup.scala 31:38]
  assign _T_205 = io_finst_inst & 32'hfffffc1f; // @[Lookup.scala 31:38]
  assign _T_206 = 32'hd61f0000 == _T_205; // @[Lookup.scala 31:38]
  assign _T_208 = 32'hd63f0000 == _T_205; // @[Lookup.scala 31:38]
  assign _T_210 = 32'hd65f0000 == _T_205; // @[Lookup.scala 31:38]
  assign _T_211 = io_finst_inst & 32'hff000000; // @[Lookup.scala 31:38]
  assign _T_212 = 32'h36000000 == _T_211; // @[Lookup.scala 31:38]
  assign _T_214 = 32'h37000000 == _T_211; // @[Lookup.scala 31:38]
  assign _T_216 = 32'hb6000000 == _T_211; // @[Lookup.scala 31:38]
  assign _T_218 = 32'hb7000000 == _T_211; // @[Lookup.scala 31:38]
  assign _T_219 = io_finst_inst & 32'hff000010; // @[Lookup.scala 31:38]
  assign _T_220 = 32'h54000000 == _T_219; // @[Lookup.scala 31:38]
  assign _T_222 = 32'h34000000 == _T_211; // @[Lookup.scala 31:38]
  assign _T_224 = 32'h35000000 == _T_211; // @[Lookup.scala 31:38]
  assign _T_226 = 32'hb4000000 == _T_211; // @[Lookup.scala 31:38]
  assign _T_228 = 32'hb5000000 == _T_211; // @[Lookup.scala 31:38]
  assign _T_230 = 32'h28800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_232 = 32'ha8800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_234 = 32'h28c00000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_236 = 32'ha8c00000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_238 = 32'h68c00000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_240 = 32'h29000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_242 = 32'ha9000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_244 = 32'h29400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_246 = 32'ha9400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_248 = 32'h69400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_250 = 32'h29800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_252 = 32'ha9800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_254 = 32'h29c00000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_256 = 32'ha9c00000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_258 = 32'h69c00000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_259 = io_finst_inst & 32'hffe04c00; // @[Lookup.scala 31:38]
  assign _T_260 = 32'h38204800 == _T_259; // @[Lookup.scala 31:38]
  assign _T_262 = 32'h78204800 == _T_259; // @[Lookup.scala 31:38]
  assign _T_264 = 32'hb8204800 == _T_259; // @[Lookup.scala 31:38]
  assign _T_266 = 32'hf8204800 == _T_259; // @[Lookup.scala 31:38]
  assign _T_268 = 32'h38604800 == _T_259; // @[Lookup.scala 31:38]
  assign _T_270 = 32'h78604800 == _T_259; // @[Lookup.scala 31:38]
  assign _T_272 = 32'hb8604800 == _T_259; // @[Lookup.scala 31:38]
  assign _T_274 = 32'hf8604800 == _T_259; // @[Lookup.scala 31:38]
  assign _T_276 = 32'h39000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_278 = 32'h79000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_280 = 32'hb9000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_282 = 32'hf9000000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_284 = 32'h39400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_286 = 32'h79400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_288 = 32'hb9400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_290 = 32'hf9400000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_292 = 32'hb9800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_294 = 32'h39800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_296 = 32'h39c00000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_298 = 32'h79800000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_300 = 32'h79c00000 == _T_43; // @[Lookup.scala 31:38]
  assign _T_302 = 32'h38000000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_304 = 32'h38400000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_306 = 32'h38800000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_308 = 32'h38c00000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_310 = 32'h78000000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_312 = 32'h78400000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_314 = 32'h78800000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_316 = 32'h78c00000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_318 = 32'hb8000000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_320 = 32'hb8400000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_322 = 32'hb8800000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_324 = 32'hf8000000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_326 = 32'hf8400000 == _T_85; // @[Lookup.scala 31:38]
  assign _T_328 = 32'h38000400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_330 = 32'h38400400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_332 = 32'h38800400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_334 = 32'h38c00400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_336 = 32'h78000400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_338 = 32'h78400400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_340 = 32'h78800400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_342 = 32'h78c00400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_344 = 32'hb8000400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_346 = 32'hb8400400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_348 = 32'hb8800400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_350 = 32'hf8000400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_352 = 32'hf8400400 == _T_85; // @[Lookup.scala 31:38]
  assign _T_354 = 32'h38000c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_356 = 32'h38400c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_358 = 32'h38800c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_360 = 32'h38c00c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_362 = 32'h78000c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_364 = 32'h78400c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_366 = 32'h78800c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_368 = 32'h78c00c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_370 = 32'hb8000c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_372 = 32'hb8400c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_374 = 32'hb8800c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_376 = 32'hf8000c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_378 = 32'hf8400c00 == _T_85; // @[Lookup.scala 31:38]
  assign _T_379 = _T_378 ? 5'h13 : 5'h0; // @[Lookup.scala 33:37]
  assign _T_380 = _T_376 ? 5'h13 : _T_379; // @[Lookup.scala 33:37]
  assign _T_381 = _T_374 ? 5'h13 : _T_380; // @[Lookup.scala 33:37]
  assign _T_382 = _T_372 ? 5'h13 : _T_381; // @[Lookup.scala 33:37]
  assign _T_383 = _T_370 ? 5'h13 : _T_382; // @[Lookup.scala 33:37]
  assign _T_384 = _T_368 ? 5'h13 : _T_383; // @[Lookup.scala 33:37]
  assign _T_385 = _T_366 ? 5'h13 : _T_384; // @[Lookup.scala 33:37]
  assign _T_386 = _T_364 ? 5'h13 : _T_385; // @[Lookup.scala 33:37]
  assign _T_387 = _T_362 ? 5'h13 : _T_386; // @[Lookup.scala 33:37]
  assign _T_388 = _T_360 ? 5'h13 : _T_387; // @[Lookup.scala 33:37]
  assign _T_389 = _T_358 ? 5'h13 : _T_388; // @[Lookup.scala 33:37]
  assign _T_390 = _T_356 ? 5'h13 : _T_389; // @[Lookup.scala 33:37]
  assign _T_391 = _T_354 ? 5'h13 : _T_390; // @[Lookup.scala 33:37]
  assign _T_392 = _T_352 ? 5'h11 : _T_391; // @[Lookup.scala 33:37]
  assign _T_393 = _T_350 ? 5'h11 : _T_392; // @[Lookup.scala 33:37]
  assign _T_394 = _T_348 ? 5'h11 : _T_393; // @[Lookup.scala 33:37]
  assign _T_395 = _T_346 ? 5'h11 : _T_394; // @[Lookup.scala 33:37]
  assign _T_396 = _T_344 ? 5'h11 : _T_395; // @[Lookup.scala 33:37]
  assign _T_397 = _T_342 ? 5'h11 : _T_396; // @[Lookup.scala 33:37]
  assign _T_398 = _T_340 ? 5'h11 : _T_397; // @[Lookup.scala 33:37]
  assign _T_399 = _T_338 ? 5'h11 : _T_398; // @[Lookup.scala 33:37]
  assign _T_400 = _T_336 ? 5'h11 : _T_399; // @[Lookup.scala 33:37]
  assign _T_401 = _T_334 ? 5'h11 : _T_400; // @[Lookup.scala 33:37]
  assign _T_402 = _T_332 ? 5'h11 : _T_401; // @[Lookup.scala 33:37]
  assign _T_403 = _T_330 ? 5'h11 : _T_402; // @[Lookup.scala 33:37]
  assign _T_404 = _T_328 ? 5'h11 : _T_403; // @[Lookup.scala 33:37]
  assign _T_405 = _T_326 ? 5'h10 : _T_404; // @[Lookup.scala 33:37]
  assign _T_406 = _T_324 ? 5'h10 : _T_405; // @[Lookup.scala 33:37]
  assign _T_407 = _T_322 ? 5'h10 : _T_406; // @[Lookup.scala 33:37]
  assign _T_408 = _T_320 ? 5'h10 : _T_407; // @[Lookup.scala 33:37]
  assign _T_409 = _T_318 ? 5'h10 : _T_408; // @[Lookup.scala 33:37]
  assign _T_410 = _T_316 ? 5'h10 : _T_409; // @[Lookup.scala 33:37]
  assign _T_411 = _T_314 ? 5'h10 : _T_410; // @[Lookup.scala 33:37]
  assign _T_412 = _T_312 ? 5'h10 : _T_411; // @[Lookup.scala 33:37]
  assign _T_413 = _T_310 ? 5'h10 : _T_412; // @[Lookup.scala 33:37]
  assign _T_414 = _T_308 ? 5'h10 : _T_413; // @[Lookup.scala 33:37]
  assign _T_415 = _T_306 ? 5'h10 : _T_414; // @[Lookup.scala 33:37]
  assign _T_416 = _T_304 ? 5'h10 : _T_415; // @[Lookup.scala 33:37]
  assign _T_417 = _T_302 ? 5'h10 : _T_416; // @[Lookup.scala 33:37]
  assign _T_418 = _T_300 ? 5'h14 : _T_417; // @[Lookup.scala 33:37]
  assign _T_419 = _T_298 ? 5'h14 : _T_418; // @[Lookup.scala 33:37]
  assign _T_420 = _T_296 ? 5'h14 : _T_419; // @[Lookup.scala 33:37]
  assign _T_421 = _T_294 ? 5'h14 : _T_420; // @[Lookup.scala 33:37]
  assign _T_422 = _T_292 ? 5'h14 : _T_421; // @[Lookup.scala 33:37]
  assign _T_423 = _T_290 ? 5'h14 : _T_422; // @[Lookup.scala 33:37]
  assign _T_424 = _T_288 ? 5'h14 : _T_423; // @[Lookup.scala 33:37]
  assign _T_425 = _T_286 ? 5'h14 : _T_424; // @[Lookup.scala 33:37]
  assign _T_426 = _T_284 ? 5'h14 : _T_425; // @[Lookup.scala 33:37]
  assign _T_427 = _T_282 ? 5'h14 : _T_426; // @[Lookup.scala 33:37]
  assign _T_428 = _T_280 ? 5'h14 : _T_427; // @[Lookup.scala 33:37]
  assign _T_429 = _T_278 ? 5'h14 : _T_428; // @[Lookup.scala 33:37]
  assign _T_430 = _T_276 ? 5'h14 : _T_429; // @[Lookup.scala 33:37]
  assign _T_431 = _T_274 ? 5'h12 : _T_430; // @[Lookup.scala 33:37]
  assign _T_432 = _T_272 ? 5'h12 : _T_431; // @[Lookup.scala 33:37]
  assign _T_433 = _T_270 ? 5'h12 : _T_432; // @[Lookup.scala 33:37]
  assign _T_434 = _T_268 ? 5'h12 : _T_433; // @[Lookup.scala 33:37]
  assign _T_435 = _T_266 ? 5'h12 : _T_434; // @[Lookup.scala 33:37]
  assign _T_436 = _T_264 ? 5'h12 : _T_435; // @[Lookup.scala 33:37]
  assign _T_437 = _T_262 ? 5'h12 : _T_436; // @[Lookup.scala 33:37]
  assign _T_438 = _T_260 ? 5'h12 : _T_437; // @[Lookup.scala 33:37]
  assign _T_439 = _T_258 ? 5'h17 : _T_438; // @[Lookup.scala 33:37]
  assign _T_440 = _T_256 ? 5'h17 : _T_439; // @[Lookup.scala 33:37]
  assign _T_441 = _T_254 ? 5'h17 : _T_440; // @[Lookup.scala 33:37]
  assign _T_442 = _T_252 ? 5'h17 : _T_441; // @[Lookup.scala 33:37]
  assign _T_443 = _T_250 ? 5'h17 : _T_442; // @[Lookup.scala 33:37]
  assign _T_444 = _T_248 ? 5'h16 : _T_443; // @[Lookup.scala 33:37]
  assign _T_445 = _T_246 ? 5'h16 : _T_444; // @[Lookup.scala 33:37]
  assign _T_446 = _T_244 ? 5'h16 : _T_445; // @[Lookup.scala 33:37]
  assign _T_447 = _T_242 ? 5'h16 : _T_446; // @[Lookup.scala 33:37]
  assign _T_448 = _T_240 ? 5'h16 : _T_447; // @[Lookup.scala 33:37]
  assign _T_449 = _T_238 ? 5'h15 : _T_448; // @[Lookup.scala 33:37]
  assign _T_450 = _T_236 ? 5'h15 : _T_449; // @[Lookup.scala 33:37]
  assign _T_451 = _T_234 ? 5'h15 : _T_450; // @[Lookup.scala 33:37]
  assign _T_452 = _T_232 ? 5'h15 : _T_451; // @[Lookup.scala 33:37]
  assign _T_453 = _T_230 ? 5'h15 : _T_452; // @[Lookup.scala 33:37]
  assign _T_454 = _T_228 ? 5'h1b : _T_453; // @[Lookup.scala 33:37]
  assign _T_455 = _T_226 ? 5'h1b : _T_454; // @[Lookup.scala 33:37]
  assign _T_456 = _T_224 ? 5'h1b : _T_455; // @[Lookup.scala 33:37]
  assign _T_457 = _T_222 ? 5'h1b : _T_456; // @[Lookup.scala 33:37]
  assign _T_458 = _T_220 ? 5'h19 : _T_457; // @[Lookup.scala 33:37]
  assign _T_459 = _T_218 ? 5'h1a : _T_458; // @[Lookup.scala 33:37]
  assign _T_460 = _T_216 ? 5'h1a : _T_459; // @[Lookup.scala 33:37]
  assign _T_461 = _T_214 ? 5'h1a : _T_460; // @[Lookup.scala 33:37]
  assign _T_462 = _T_212 ? 5'h1a : _T_461; // @[Lookup.scala 33:37]
  assign _T_463 = _T_210 ? 5'h1c : _T_462; // @[Lookup.scala 33:37]
  assign _T_464 = _T_208 ? 5'h1c : _T_463; // @[Lookup.scala 33:37]
  assign _T_465 = _T_206 ? 5'h1c : _T_464; // @[Lookup.scala 33:37]
  assign _T_466 = _T_204 ? 5'h18 : _T_465; // @[Lookup.scala 33:37]
  assign _T_467 = _T_202 ? 5'h18 : _T_466; // @[Lookup.scala 33:37]
  assign _T_468 = _T_200 ? 5'he : _T_467; // @[Lookup.scala 33:37]
  assign _T_469 = _T_198 ? 5'hd : _T_468; // @[Lookup.scala 33:37]
  assign _T_470 = _T_196 ? 5'hd : _T_469; // @[Lookup.scala 33:37]
  assign _T_471 = _T_194 ? 5'hd : _T_470; // @[Lookup.scala 33:37]
  assign _T_472 = _T_192 ? 5'hd : _T_471; // @[Lookup.scala 33:37]
  assign _T_473 = _T_190 ? 5'hd : _T_472; // @[Lookup.scala 33:37]
  assign _T_474 = _T_188 ? 5'hd : _T_473; // @[Lookup.scala 33:37]
  assign _T_475 = _T_186 ? 5'hd : _T_474; // @[Lookup.scala 33:37]
  assign _T_476 = _T_184 ? 5'hd : _T_475; // @[Lookup.scala 33:37]
  assign _T_477 = _T_182 ? 5'hc : _T_476; // @[Lookup.scala 33:37]
  assign _T_478 = _T_180 ? 5'hc : _T_477; // @[Lookup.scala 33:37]
  assign _T_479 = _T_178 ? 5'hc : _T_478; // @[Lookup.scala 33:37]
  assign _T_480 = _T_176 ? 5'hc : _T_479; // @[Lookup.scala 33:37]
  assign _T_481 = _T_174 ? 5'hc : _T_480; // @[Lookup.scala 33:37]
  assign _T_482 = _T_172 ? 5'hc : _T_481; // @[Lookup.scala 33:37]
  assign _T_483 = _T_170 ? 5'hc : _T_482; // @[Lookup.scala 33:37]
  assign _T_484 = _T_168 ? 5'hc : _T_483; // @[Lookup.scala 33:37]
  assign _T_485 = _T_166 ? 5'hc : _T_484; // @[Lookup.scala 33:37]
  assign _T_486 = _T_164 ? 5'hc : _T_485; // @[Lookup.scala 33:37]
  assign _T_487 = _T_162 ? 5'hc : _T_486; // @[Lookup.scala 33:37]
  assign _T_488 = _T_160 ? 5'h8 : _T_487; // @[Lookup.scala 33:37]
  assign _T_489 = _T_158 ? 5'h8 : _T_488; // @[Lookup.scala 33:37]
  assign _T_490 = _T_156 ? 5'h8 : _T_489; // @[Lookup.scala 33:37]
  assign _T_491 = _T_154 ? 5'h8 : _T_490; // @[Lookup.scala 33:37]
  assign _T_492 = _T_152 ? 5'h8 : _T_491; // @[Lookup.scala 33:37]
  assign _T_493 = _T_150 ? 5'h8 : _T_492; // @[Lookup.scala 33:37]
  assign _T_494 = _T_148 ? 5'h8 : _T_493; // @[Lookup.scala 33:37]
  assign _T_495 = _T_146 ? 5'h8 : _T_494; // @[Lookup.scala 33:37]
  assign _T_496 = _T_144 ? 5'h8 : _T_495; // @[Lookup.scala 33:37]
  assign _T_497 = _T_142 ? 5'h8 : _T_496; // @[Lookup.scala 33:37]
  assign _T_498 = _T_140 ? 5'h8 : _T_497; // @[Lookup.scala 33:37]
  assign _T_499 = _T_138 ? 5'h8 : _T_498; // @[Lookup.scala 33:37]
  assign _T_500 = _T_136 ? 5'h9 : _T_499; // @[Lookup.scala 33:37]
  assign _T_501 = _T_134 ? 5'h9 : _T_500; // @[Lookup.scala 33:37]
  assign _T_502 = _T_132 ? 5'h9 : _T_501; // @[Lookup.scala 33:37]
  assign _T_503 = _T_130 ? 5'h9 : _T_502; // @[Lookup.scala 33:37]
  assign _T_504 = _T_128 ? 5'h9 : _T_503; // @[Lookup.scala 33:37]
  assign _T_505 = _T_126 ? 5'h9 : _T_504; // @[Lookup.scala 33:37]
  assign _T_506 = _T_124 ? 5'h9 : _T_505; // @[Lookup.scala 33:37]
  assign _T_507 = _T_122 ? 5'h9 : _T_506; // @[Lookup.scala 33:37]
  assign _T_508 = _T_120 ? 5'h9 : _T_507; // @[Lookup.scala 33:37]
  assign _T_509 = _T_118 ? 5'h9 : _T_508; // @[Lookup.scala 33:37]
  assign _T_510 = _T_116 ? 5'h9 : _T_509; // @[Lookup.scala 33:37]
  assign _T_511 = _T_114 ? 5'h9 : _T_510; // @[Lookup.scala 33:37]
  assign _T_512 = _T_112 ? 5'h5 : _T_511; // @[Lookup.scala 33:37]
  assign _T_513 = _T_110 ? 5'h5 : _T_512; // @[Lookup.scala 33:37]
  assign _T_514 = _T_108 ? 5'h5 : _T_513; // @[Lookup.scala 33:37]
  assign _T_515 = _T_106 ? 5'h4 : _T_514; // @[Lookup.scala 33:37]
  assign _T_516 = _T_104 ? 5'h4 : _T_515; // @[Lookup.scala 33:37]
  assign _T_517 = _T_102 ? 5'h4 : _T_516; // @[Lookup.scala 33:37]
  assign _T_518 = _T_100 ? 5'h6 : _T_517; // @[Lookup.scala 33:37]
  assign _T_519 = _T_98 ? 5'h6 : _T_518; // @[Lookup.scala 33:37]
  assign _T_520 = _T_96 ? 5'h6 : _T_519; // @[Lookup.scala 33:37]
  assign _T_521 = _T_94 ? 5'h6 : _T_520; // @[Lookup.scala 33:37]
  assign _T_522 = _T_92 ? 5'h6 : _T_521; // @[Lookup.scala 33:37]
  assign _T_523 = _T_90 ? 5'h6 : _T_522; // @[Lookup.scala 33:37]
  assign _T_524 = _T_88 ? 5'h6 : _T_523; // @[Lookup.scala 33:37]
  assign _T_525 = _T_86 ? 5'h6 : _T_524; // @[Lookup.scala 33:37]
  assign _T_526 = _T_84 ? 5'hb : _T_525; // @[Lookup.scala 33:37]
  assign _T_527 = _T_82 ? 5'hb : _T_526; // @[Lookup.scala 33:37]
  assign _T_528 = _T_80 ? 5'hb : _T_527; // @[Lookup.scala 33:37]
  assign _T_529 = _T_78 ? 5'hb : _T_528; // @[Lookup.scala 33:37]
  assign _T_530 = _T_76 ? 5'hb : _T_529; // @[Lookup.scala 33:37]
  assign _T_531 = _T_74 ? 5'hb : _T_530; // @[Lookup.scala 33:37]
  assign _T_532 = _T_72 ? 5'ha : _T_531; // @[Lookup.scala 33:37]
  assign _T_533 = _T_70 ? 5'ha : _T_532; // @[Lookup.scala 33:37]
  assign _T_534 = _T_68 ? 5'ha : _T_533; // @[Lookup.scala 33:37]
  assign _T_535 = _T_66 ? 5'ha : _T_534; // @[Lookup.scala 33:37]
  assign _T_536 = _T_64 ? 5'ha : _T_535; // @[Lookup.scala 33:37]
  assign _T_537 = _T_62 ? 5'ha : _T_536; // @[Lookup.scala 33:37]
  assign _T_538 = _T_60 ? 5'h2 : _T_537; // @[Lookup.scala 33:37]
  assign _T_539 = _T_58 ? 5'h2 : _T_538; // @[Lookup.scala 33:37]
  assign _T_540 = _T_56 ? 5'h2 : _T_539; // @[Lookup.scala 33:37]
  assign _T_541 = _T_54 ? 5'h2 : _T_540; // @[Lookup.scala 33:37]
  assign _T_542 = _T_52 ? 5'h2 : _T_541; // @[Lookup.scala 33:37]
  assign _T_543 = _T_50 ? 5'h2 : _T_542; // @[Lookup.scala 33:37]
  assign _T_544 = _T_48 ? 5'h2 : _T_543; // @[Lookup.scala 33:37]
  assign _T_545 = _T_46 ? 5'h2 : _T_544; // @[Lookup.scala 33:37]
  assign _T_546 = _T_44 ? 5'h2 : _T_545; // @[Lookup.scala 33:37]
  assign _T_547 = _T_42 ? 5'h2 : _T_546; // @[Lookup.scala 33:37]
  assign _T_548 = _T_40 ? 5'h1 : _T_547; // @[Lookup.scala 33:37]
  assign _T_549 = _T_38 ? 5'h1 : _T_548; // @[Lookup.scala 33:37]
  assign _T_550 = _T_36 ? 5'h1 : _T_549; // @[Lookup.scala 33:37]
  assign _T_551 = _T_34 ? 5'h1 : _T_550; // @[Lookup.scala 33:37]
  assign _T_552 = _T_32 ? 5'h1 : _T_551; // @[Lookup.scala 33:37]
  assign _T_553 = _T_30 ? 5'h1 : _T_552; // @[Lookup.scala 33:37]
  assign _T_554 = _T_28 ? 5'h1 : _T_553; // @[Lookup.scala 33:37]
  assign _T_555 = _T_26 ? 5'h1 : _T_554; // @[Lookup.scala 33:37]
  assign _T_556 = _T_24 ? 5'h1 : _T_555; // @[Lookup.scala 33:37]
  assign _T_557 = _T_22 ? 5'h1 : _T_556; // @[Lookup.scala 33:37]
  assign _T_558 = _T_20 ? 5'h1 : _T_557; // @[Lookup.scala 33:37]
  assign _T_559 = _T_18 ? 5'h1 : _T_558; // @[Lookup.scala 33:37]
  assign _T_560 = _T_16 ? 5'h1 : _T_559; // @[Lookup.scala 33:37]
  assign _T_561 = _T_14 ? 5'h1 : _T_560; // @[Lookup.scala 33:37]
  assign _T_562 = _T_12 ? 5'h1 : _T_561; // @[Lookup.scala 33:37]
  assign _T_563 = _T_10 ? 5'h1 : _T_562; // @[Lookup.scala 33:37]
  assign _T_564 = _T_8 ? 5'h1 : _T_563; // @[Lookup.scala 33:37]
  assign _T_565 = _T_6 ? 5'h1 : _T_564; // @[Lookup.scala 33:37]
  assign _T_566 = _T_4 ? 5'h3 : _T_565; // @[Lookup.scala 33:37]
  assign dinst_itype = _T_2 ? 5'h3 : _T_566; // @[Lookup.scala 33:37]
  assign _T_568 = _T_378 ? 4'h7 : 4'h0; // @[Lookup.scala 33:37]
  assign _T_569 = _T_376 ? 4'h3 : _T_568; // @[Lookup.scala 33:37]
  assign _T_570 = _T_374 ? 4'he : _T_569; // @[Lookup.scala 33:37]
  assign _T_571 = _T_372 ? 4'h6 : _T_570; // @[Lookup.scala 33:37]
  assign _T_572 = _T_370 ? 4'h2 : _T_571; // @[Lookup.scala 33:37]
  assign _T_573 = _T_368 ? 4'hd : _T_572; // @[Lookup.scala 33:37]
  assign _T_574 = _T_366 ? 4'hd : _T_573; // @[Lookup.scala 33:37]
  assign _T_575 = _T_364 ? 4'h5 : _T_574; // @[Lookup.scala 33:37]
  assign _T_576 = _T_362 ? 4'h1 : _T_575; // @[Lookup.scala 33:37]
  assign _T_577 = _T_360 ? 4'hc : _T_576; // @[Lookup.scala 33:37]
  assign _T_578 = _T_358 ? 4'hc : _T_577; // @[Lookup.scala 33:37]
  assign _T_579 = _T_356 ? 4'h4 : _T_578; // @[Lookup.scala 33:37]
  assign _T_580 = _T_354 ? 4'h0 : _T_579; // @[Lookup.scala 33:37]
  assign _T_581 = _T_352 ? 4'h7 : _T_580; // @[Lookup.scala 33:37]
  assign _T_582 = _T_350 ? 4'h3 : _T_581; // @[Lookup.scala 33:37]
  assign _T_583 = _T_348 ? 4'he : _T_582; // @[Lookup.scala 33:37]
  assign _T_584 = _T_346 ? 4'h6 : _T_583; // @[Lookup.scala 33:37]
  assign _T_585 = _T_344 ? 4'h2 : _T_584; // @[Lookup.scala 33:37]
  assign _T_586 = _T_342 ? 4'hd : _T_585; // @[Lookup.scala 33:37]
  assign _T_587 = _T_340 ? 4'hd : _T_586; // @[Lookup.scala 33:37]
  assign _T_588 = _T_338 ? 4'h5 : _T_587; // @[Lookup.scala 33:37]
  assign _T_589 = _T_336 ? 4'h1 : _T_588; // @[Lookup.scala 33:37]
  assign _T_590 = _T_334 ? 4'hc : _T_589; // @[Lookup.scala 33:37]
  assign _T_591 = _T_332 ? 4'hc : _T_590; // @[Lookup.scala 33:37]
  assign _T_592 = _T_330 ? 4'h4 : _T_591; // @[Lookup.scala 33:37]
  assign _T_593 = _T_328 ? 4'h0 : _T_592; // @[Lookup.scala 33:37]
  assign _T_594 = _T_326 ? 4'h7 : _T_593; // @[Lookup.scala 33:37]
  assign _T_595 = _T_324 ? 4'h3 : _T_594; // @[Lookup.scala 33:37]
  assign _T_596 = _T_322 ? 4'he : _T_595; // @[Lookup.scala 33:37]
  assign _T_597 = _T_320 ? 4'h6 : _T_596; // @[Lookup.scala 33:37]
  assign _T_598 = _T_318 ? 4'h2 : _T_597; // @[Lookup.scala 33:37]
  assign _T_599 = _T_316 ? 4'hd : _T_598; // @[Lookup.scala 33:37]
  assign _T_600 = _T_314 ? 4'hd : _T_599; // @[Lookup.scala 33:37]
  assign _T_601 = _T_312 ? 4'h5 : _T_600; // @[Lookup.scala 33:37]
  assign _T_602 = _T_310 ? 4'h1 : _T_601; // @[Lookup.scala 33:37]
  assign _T_603 = _T_308 ? 4'hc : _T_602; // @[Lookup.scala 33:37]
  assign _T_604 = _T_306 ? 4'hc : _T_603; // @[Lookup.scala 33:37]
  assign _T_605 = _T_304 ? 4'h4 : _T_604; // @[Lookup.scala 33:37]
  assign _T_606 = _T_302 ? 4'h0 : _T_605; // @[Lookup.scala 33:37]
  assign _T_607 = _T_300 ? 4'hd : _T_606; // @[Lookup.scala 33:37]
  assign _T_608 = _T_298 ? 4'hd : _T_607; // @[Lookup.scala 33:37]
  assign _T_609 = _T_296 ? 4'hc : _T_608; // @[Lookup.scala 33:37]
  assign _T_610 = _T_294 ? 4'hc : _T_609; // @[Lookup.scala 33:37]
  assign _T_611 = _T_292 ? 4'he : _T_610; // @[Lookup.scala 33:37]
  assign _T_612 = _T_290 ? 4'h7 : _T_611; // @[Lookup.scala 33:37]
  assign _T_613 = _T_288 ? 4'h6 : _T_612; // @[Lookup.scala 33:37]
  assign _T_614 = _T_286 ? 4'h5 : _T_613; // @[Lookup.scala 33:37]
  assign _T_615 = _T_284 ? 4'h4 : _T_614; // @[Lookup.scala 33:37]
  assign _T_616 = _T_282 ? 4'h3 : _T_615; // @[Lookup.scala 33:37]
  assign _T_617 = _T_280 ? 4'h2 : _T_616; // @[Lookup.scala 33:37]
  assign _T_618 = _T_278 ? 4'h1 : _T_617; // @[Lookup.scala 33:37]
  assign _T_619 = _T_276 ? 4'h0 : _T_618; // @[Lookup.scala 33:37]
  assign _T_620 = _T_274 ? 4'h7 : _T_619; // @[Lookup.scala 33:37]
  assign _T_621 = _T_272 ? 4'h6 : _T_620; // @[Lookup.scala 33:37]
  assign _T_622 = _T_270 ? 4'h5 : _T_621; // @[Lookup.scala 33:37]
  assign _T_623 = _T_268 ? 4'h4 : _T_622; // @[Lookup.scala 33:37]
  assign _T_624 = _T_266 ? 4'h3 : _T_623; // @[Lookup.scala 33:37]
  assign _T_625 = _T_264 ? 4'h2 : _T_624; // @[Lookup.scala 33:37]
  assign _T_626 = _T_262 ? 4'h1 : _T_625; // @[Lookup.scala 33:37]
  assign _T_627 = _T_260 ? 4'h0 : _T_626; // @[Lookup.scala 33:37]
  assign _T_628 = _T_258 ? 4'hf : _T_627; // @[Lookup.scala 33:37]
  assign _T_629 = _T_256 ? 4'h7 : _T_628; // @[Lookup.scala 33:37]
  assign _T_630 = _T_254 ? 4'h6 : _T_629; // @[Lookup.scala 33:37]
  assign _T_631 = _T_252 ? 4'h3 : _T_630; // @[Lookup.scala 33:37]
  assign _T_632 = _T_250 ? 4'h2 : _T_631; // @[Lookup.scala 33:37]
  assign _T_633 = _T_248 ? 4'hf : _T_632; // @[Lookup.scala 33:37]
  assign _T_634 = _T_246 ? 4'h7 : _T_633; // @[Lookup.scala 33:37]
  assign _T_635 = _T_244 ? 4'h6 : _T_634; // @[Lookup.scala 33:37]
  assign _T_636 = _T_242 ? 4'h3 : _T_635; // @[Lookup.scala 33:37]
  assign _T_637 = _T_240 ? 4'h2 : _T_636; // @[Lookup.scala 33:37]
  assign _T_638 = _T_238 ? 4'hf : _T_637; // @[Lookup.scala 33:37]
  assign _T_639 = _T_236 ? 4'h7 : _T_638; // @[Lookup.scala 33:37]
  assign _T_640 = _T_234 ? 4'h6 : _T_639; // @[Lookup.scala 33:37]
  assign _T_641 = _T_232 ? 4'h3 : _T_640; // @[Lookup.scala 33:37]
  assign _T_642 = _T_230 ? 4'h2 : _T_641; // @[Lookup.scala 33:37]
  assign _T_643 = _T_228 ? 4'h1 : _T_642; // @[Lookup.scala 33:37]
  assign _T_644 = _T_226 ? 4'h0 : _T_643; // @[Lookup.scala 33:37]
  assign _T_645 = _T_224 ? 4'h1 : _T_644; // @[Lookup.scala 33:37]
  assign _T_646 = _T_222 ? 4'h0 : _T_645; // @[Lookup.scala 33:37]
  assign _T_647 = _T_220 ? 4'h0 : _T_646; // @[Lookup.scala 33:37]
  assign _T_648 = _T_218 ? 4'h1 : _T_647; // @[Lookup.scala 33:37]
  assign _T_649 = _T_216 ? 4'h0 : _T_648; // @[Lookup.scala 33:37]
  assign _T_650 = _T_214 ? 4'h1 : _T_649; // @[Lookup.scala 33:37]
  assign _T_651 = _T_212 ? 4'h0 : _T_650; // @[Lookup.scala 33:37]
  assign _T_652 = _T_210 ? 4'h0 : _T_651; // @[Lookup.scala 33:37]
  assign _T_653 = _T_208 ? 4'h1 : _T_652; // @[Lookup.scala 33:37]
  assign _T_654 = _T_206 ? 4'h0 : _T_653; // @[Lookup.scala 33:37]
  assign _T_655 = _T_204 ? 4'h1 : _T_654; // @[Lookup.scala 33:37]
  assign _T_656 = _T_202 ? 4'h0 : _T_655; // @[Lookup.scala 33:37]
  assign _T_657 = _T_200 ? 4'h0 : _T_656; // @[Lookup.scala 33:37]
  assign _T_658 = _T_198 ? 4'h3 : _T_657; // @[Lookup.scala 33:37]
  assign _T_659 = _T_196 ? 4'h2 : _T_658; // @[Lookup.scala 33:37]
  assign _T_660 = _T_194 ? 4'h1 : _T_659; // @[Lookup.scala 33:37]
  assign _T_661 = _T_192 ? 4'h0 : _T_660; // @[Lookup.scala 33:37]
  assign _T_662 = _T_190 ? 4'h3 : _T_661; // @[Lookup.scala 33:37]
  assign _T_663 = _T_188 ? 4'h2 : _T_662; // @[Lookup.scala 33:37]
  assign _T_664 = _T_186 ? 4'h1 : _T_663; // @[Lookup.scala 33:37]
  assign _T_665 = _T_184 ? 4'h0 : _T_664; // @[Lookup.scala 33:37]
  assign _T_666 = _T_182 ? 4'h5 : _T_665; // @[Lookup.scala 33:37]
  assign _T_667 = _T_180 ? 4'h4 : _T_666; // @[Lookup.scala 33:37]
  assign _T_668 = _T_178 ? 4'h3 : _T_667; // @[Lookup.scala 33:37]
  assign _T_669 = _T_176 ? 4'h2 : _T_668; // @[Lookup.scala 33:37]
  assign _T_670 = _T_174 ? 4'h1 : _T_669; // @[Lookup.scala 33:37]
  assign _T_671 = _T_172 ? 4'h0 : _T_670; // @[Lookup.scala 33:37]
  assign _T_672 = _T_170 ? 4'h5 : _T_671; // @[Lookup.scala 33:37]
  assign _T_673 = _T_168 ? 4'h4 : _T_672; // @[Lookup.scala 33:37]
  assign _T_674 = _T_166 ? 4'h2 : _T_673; // @[Lookup.scala 33:37]
  assign _T_675 = _T_164 ? 4'h1 : _T_674; // @[Lookup.scala 33:37]
  assign _T_676 = _T_162 ? 4'h0 : _T_675; // @[Lookup.scala 33:37]
  assign _T_677 = _T_160 ? 4'h1 : _T_676; // @[Lookup.scala 33:37]
  assign _T_678 = _T_158 ? 4'h1 : _T_677; // @[Lookup.scala 33:37]
  assign _T_679 = _T_156 ? 4'h0 : _T_678; // @[Lookup.scala 33:37]
  assign _T_680 = _T_154 ? 4'h0 : _T_679; // @[Lookup.scala 33:37]
  assign _T_681 = _T_152 ? 4'h0 : _T_680; // @[Lookup.scala 33:37]
  assign _T_682 = _T_150 ? 4'h1 : _T_681; // @[Lookup.scala 33:37]
  assign _T_683 = _T_148 ? 4'h1 : _T_682; // @[Lookup.scala 33:37]
  assign _T_684 = _T_146 ? 4'h1 : _T_683; // @[Lookup.scala 33:37]
  assign _T_685 = _T_144 ? 4'h0 : _T_684; // @[Lookup.scala 33:37]
  assign _T_686 = _T_142 ? 4'h0 : _T_685; // @[Lookup.scala 33:37]
  assign _T_687 = _T_140 ? 4'h0 : _T_686; // @[Lookup.scala 33:37]
  assign _T_688 = _T_138 ? 4'h1 : _T_687; // @[Lookup.scala 33:37]
  assign _T_689 = _T_136 ? 4'h1 : _T_688; // @[Lookup.scala 33:37]
  assign _T_690 = _T_134 ? 4'h1 : _T_689; // @[Lookup.scala 33:37]
  assign _T_691 = _T_132 ? 4'h0 : _T_690; // @[Lookup.scala 33:37]
  assign _T_692 = _T_130 ? 4'h0 : _T_691; // @[Lookup.scala 33:37]
  assign _T_693 = _T_128 ? 4'h0 : _T_692; // @[Lookup.scala 33:37]
  assign _T_694 = _T_126 ? 4'h1 : _T_693; // @[Lookup.scala 33:37]
  assign _T_695 = _T_124 ? 4'h1 : _T_694; // @[Lookup.scala 33:37]
  assign _T_696 = _T_122 ? 4'h1 : _T_695; // @[Lookup.scala 33:37]
  assign _T_697 = _T_120 ? 4'h0 : _T_696; // @[Lookup.scala 33:37]
  assign _T_698 = _T_118 ? 4'h0 : _T_697; // @[Lookup.scala 33:37]
  assign _T_699 = _T_116 ? 4'h0 : _T_698; // @[Lookup.scala 33:37]
  assign _T_700 = _T_114 ? 4'h1 : _T_699; // @[Lookup.scala 33:37]
  assign _T_701 = _T_112 ? 4'h1 : _T_700; // @[Lookup.scala 33:37]
  assign _T_702 = _T_110 ? 4'h1 : _T_701; // @[Lookup.scala 33:37]
  assign _T_703 = _T_108 ? 4'h0 : _T_702; // @[Lookup.scala 33:37]
  assign _T_704 = _T_106 ? 4'h1 : _T_703; // @[Lookup.scala 33:37]
  assign _T_705 = _T_104 ? 4'h1 : _T_704; // @[Lookup.scala 33:37]
  assign _T_706 = _T_102 ? 4'h0 : _T_705; // @[Lookup.scala 33:37]
  assign _T_707 = _T_100 ? 4'h3 : _T_706; // @[Lookup.scala 33:37]
  assign _T_708 = _T_98 ? 4'h2 : _T_707; // @[Lookup.scala 33:37]
  assign _T_709 = _T_96 ? 4'h1 : _T_708; // @[Lookup.scala 33:37]
  assign _T_710 = _T_94 ? 4'h0 : _T_709; // @[Lookup.scala 33:37]
  assign _T_711 = _T_92 ? 4'h3 : _T_710; // @[Lookup.scala 33:37]
  assign _T_712 = _T_90 ? 4'h2 : _T_711; // @[Lookup.scala 33:37]
  assign _T_713 = _T_88 ? 4'h1 : _T_712; // @[Lookup.scala 33:37]
  assign _T_714 = _T_86 ? 4'h0 : _T_713; // @[Lookup.scala 33:37]
  assign _T_715 = _T_84 ? 4'h2 : _T_714; // @[Lookup.scala 33:37]
  assign _T_716 = _T_82 ? 4'h1 : _T_715; // @[Lookup.scala 33:37]
  assign _T_717 = _T_80 ? 4'h0 : _T_716; // @[Lookup.scala 33:37]
  assign _T_718 = _T_78 ? 4'h2 : _T_717; // @[Lookup.scala 33:37]
  assign _T_719 = _T_76 ? 4'h1 : _T_718; // @[Lookup.scala 33:37]
  assign _T_720 = _T_74 ? 4'h0 : _T_719; // @[Lookup.scala 33:37]
  assign _T_721 = _T_72 ? 4'h2 : _T_720; // @[Lookup.scala 33:37]
  assign _T_722 = _T_70 ? 4'h1 : _T_721; // @[Lookup.scala 33:37]
  assign _T_723 = _T_68 ? 4'h0 : _T_722; // @[Lookup.scala 33:37]
  assign _T_724 = _T_66 ? 4'h2 : _T_723; // @[Lookup.scala 33:37]
  assign _T_725 = _T_64 ? 4'h1 : _T_724; // @[Lookup.scala 33:37]
  assign _T_726 = _T_62 ? 4'h0 : _T_725; // @[Lookup.scala 33:37]
  assign _T_727 = _T_60 ? 4'h0 : _T_726; // @[Lookup.scala 33:37]
  assign _T_728 = _T_58 ? 4'h4 : _T_727; // @[Lookup.scala 33:37]
  assign _T_729 = _T_56 ? 4'h2 : _T_728; // @[Lookup.scala 33:37]
  assign _T_730 = _T_54 ? 4'h0 : _T_729; // @[Lookup.scala 33:37]
  assign _T_731 = _T_52 ? 4'h0 : _T_730; // @[Lookup.scala 33:37]
  assign _T_732 = _T_50 ? 4'h0 : _T_731; // @[Lookup.scala 33:37]
  assign _T_733 = _T_48 ? 4'h4 : _T_732; // @[Lookup.scala 33:37]
  assign _T_734 = _T_46 ? 4'h2 : _T_733; // @[Lookup.scala 33:37]
  assign _T_735 = _T_44 ? 4'h0 : _T_734; // @[Lookup.scala 33:37]
  assign _T_736 = _T_42 ? 4'h0 : _T_735; // @[Lookup.scala 33:37]
  assign _T_737 = _T_40 ? 4'h1 : _T_736; // @[Lookup.scala 33:37]
  assign _T_738 = _T_38 ? 4'h0 : _T_737; // @[Lookup.scala 33:37]
  assign _T_739 = _T_36 ? 4'h5 : _T_738; // @[Lookup.scala 33:37]
  assign _T_740 = _T_34 ? 4'h4 : _T_739; // @[Lookup.scala 33:37]
  assign _T_741 = _T_32 ? 4'h3 : _T_740; // @[Lookup.scala 33:37]
  assign _T_742 = _T_30 ? 4'h2 : _T_741; // @[Lookup.scala 33:37]
  assign _T_743 = _T_28 ? 4'h1 : _T_742; // @[Lookup.scala 33:37]
  assign _T_744 = _T_26 ? 4'h0 : _T_743; // @[Lookup.scala 33:37]
  assign _T_745 = _T_24 ? 4'h0 : _T_744; // @[Lookup.scala 33:37]
  assign _T_746 = _T_22 ? 4'h1 : _T_745; // @[Lookup.scala 33:37]
  assign _T_747 = _T_20 ? 4'h0 : _T_746; // @[Lookup.scala 33:37]
  assign _T_748 = _T_18 ? 4'h5 : _T_747; // @[Lookup.scala 33:37]
  assign _T_749 = _T_16 ? 4'h4 : _T_748; // @[Lookup.scala 33:37]
  assign _T_750 = _T_14 ? 4'h3 : _T_749; // @[Lookup.scala 33:37]
  assign _T_751 = _T_12 ? 4'h2 : _T_750; // @[Lookup.scala 33:37]
  assign _T_752 = _T_10 ? 4'h1 : _T_751; // @[Lookup.scala 33:37]
  assign _T_753 = _T_8 ? 4'h0 : _T_752; // @[Lookup.scala 33:37]
  assign _T_754 = _T_6 ? 4'h0 : _T_753; // @[Lookup.scala 33:37]
  assign _T_755 = _T_4 ? 4'h1 : _T_754; // @[Lookup.scala 33:37]
  assign _T_758 = _T_376 | _T_378; // @[Lookup.scala 33:37]
  assign _T_759 = _T_374 | _T_758; // @[Lookup.scala 33:37]
  assign _T_760 = _T_372 | _T_759; // @[Lookup.scala 33:37]
  assign _T_761 = _T_370 | _T_760; // @[Lookup.scala 33:37]
  assign _T_762 = _T_368 | _T_761; // @[Lookup.scala 33:37]
  assign _T_763 = _T_366 | _T_762; // @[Lookup.scala 33:37]
  assign _T_764 = _T_364 | _T_763; // @[Lookup.scala 33:37]
  assign _T_765 = _T_362 | _T_764; // @[Lookup.scala 33:37]
  assign _T_766 = _T_360 | _T_765; // @[Lookup.scala 33:37]
  assign _T_767 = _T_358 | _T_766; // @[Lookup.scala 33:37]
  assign _T_768 = _T_356 | _T_767; // @[Lookup.scala 33:37]
  assign _T_769 = _T_354 | _T_768; // @[Lookup.scala 33:37]
  assign _T_770 = _T_352 | _T_769; // @[Lookup.scala 33:37]
  assign _T_771 = _T_350 | _T_770; // @[Lookup.scala 33:37]
  assign _T_772 = _T_348 | _T_771; // @[Lookup.scala 33:37]
  assign _T_773 = _T_346 | _T_772; // @[Lookup.scala 33:37]
  assign _T_774 = _T_344 | _T_773; // @[Lookup.scala 33:37]
  assign _T_775 = _T_342 | _T_774; // @[Lookup.scala 33:37]
  assign _T_776 = _T_340 | _T_775; // @[Lookup.scala 33:37]
  assign _T_777 = _T_338 | _T_776; // @[Lookup.scala 33:37]
  assign _T_778 = _T_336 | _T_777; // @[Lookup.scala 33:37]
  assign _T_779 = _T_334 | _T_778; // @[Lookup.scala 33:37]
  assign _T_780 = _T_332 | _T_779; // @[Lookup.scala 33:37]
  assign _T_781 = _T_330 | _T_780; // @[Lookup.scala 33:37]
  assign _T_782 = _T_328 | _T_781; // @[Lookup.scala 33:37]
  assign _T_783 = _T_326 | _T_782; // @[Lookup.scala 33:37]
  assign _T_784 = _T_324 | _T_783; // @[Lookup.scala 33:37]
  assign _T_785 = _T_322 | _T_784; // @[Lookup.scala 33:37]
  assign _T_786 = _T_320 | _T_785; // @[Lookup.scala 33:37]
  assign _T_787 = _T_318 | _T_786; // @[Lookup.scala 33:37]
  assign _T_788 = _T_316 | _T_787; // @[Lookup.scala 33:37]
  assign _T_789 = _T_314 | _T_788; // @[Lookup.scala 33:37]
  assign _T_790 = _T_312 | _T_789; // @[Lookup.scala 33:37]
  assign _T_791 = _T_310 | _T_790; // @[Lookup.scala 33:37]
  assign _T_792 = _T_308 | _T_791; // @[Lookup.scala 33:37]
  assign _T_793 = _T_306 | _T_792; // @[Lookup.scala 33:37]
  assign _T_794 = _T_304 | _T_793; // @[Lookup.scala 33:37]
  assign _T_795 = _T_302 | _T_794; // @[Lookup.scala 33:37]
  assign _T_796 = _T_300 | _T_795; // @[Lookup.scala 33:37]
  assign _T_797 = _T_298 | _T_796; // @[Lookup.scala 33:37]
  assign _T_798 = _T_296 | _T_797; // @[Lookup.scala 33:37]
  assign _T_799 = _T_294 | _T_798; // @[Lookup.scala 33:37]
  assign _T_800 = _T_292 | _T_799; // @[Lookup.scala 33:37]
  assign _T_801 = _T_290 | _T_800; // @[Lookup.scala 33:37]
  assign _T_802 = _T_288 | _T_801; // @[Lookup.scala 33:37]
  assign _T_803 = _T_286 | _T_802; // @[Lookup.scala 33:37]
  assign _T_804 = _T_284 | _T_803; // @[Lookup.scala 33:37]
  assign _T_805 = _T_282 | _T_804; // @[Lookup.scala 33:37]
  assign _T_806 = _T_280 | _T_805; // @[Lookup.scala 33:37]
  assign _T_807 = _T_278 | _T_806; // @[Lookup.scala 33:37]
  assign _T_808 = _T_276 | _T_807; // @[Lookup.scala 33:37]
  assign _T_809 = _T_274 | _T_808; // @[Lookup.scala 33:37]
  assign _T_810 = _T_272 | _T_809; // @[Lookup.scala 33:37]
  assign _T_811 = _T_270 | _T_810; // @[Lookup.scala 33:37]
  assign _T_812 = _T_268 | _T_811; // @[Lookup.scala 33:37]
  assign _T_813 = _T_266 | _T_812; // @[Lookup.scala 33:37]
  assign _T_814 = _T_264 | _T_813; // @[Lookup.scala 33:37]
  assign _T_815 = _T_262 | _T_814; // @[Lookup.scala 33:37]
  assign _T_816 = _T_260 | _T_815; // @[Lookup.scala 33:37]
  assign _T_817 = _T_258 | _T_816; // @[Lookup.scala 33:37]
  assign _T_818 = _T_256 | _T_817; // @[Lookup.scala 33:37]
  assign _T_819 = _T_254 | _T_818; // @[Lookup.scala 33:37]
  assign _T_820 = _T_252 | _T_819; // @[Lookup.scala 33:37]
  assign _T_821 = _T_250 | _T_820; // @[Lookup.scala 33:37]
  assign _T_822 = _T_248 | _T_821; // @[Lookup.scala 33:37]
  assign _T_823 = _T_246 | _T_822; // @[Lookup.scala 33:37]
  assign _T_824 = _T_244 | _T_823; // @[Lookup.scala 33:37]
  assign _T_825 = _T_242 | _T_824; // @[Lookup.scala 33:37]
  assign _T_826 = _T_240 | _T_825; // @[Lookup.scala 33:37]
  assign _T_827 = _T_238 | _T_826; // @[Lookup.scala 33:37]
  assign _T_828 = _T_236 | _T_827; // @[Lookup.scala 33:37]
  assign _T_829 = _T_234 | _T_828; // @[Lookup.scala 33:37]
  assign _T_830 = _T_232 | _T_829; // @[Lookup.scala 33:37]
  assign _T_831 = _T_230 | _T_830; // @[Lookup.scala 33:37]
  assign _T_832 = _T_228 ? 1'h0 : _T_831; // @[Lookup.scala 33:37]
  assign _T_833 = _T_226 ? 1'h0 : _T_832; // @[Lookup.scala 33:37]
  assign _T_834 = _T_224 ? 1'h0 : _T_833; // @[Lookup.scala 33:37]
  assign _T_835 = _T_222 ? 1'h0 : _T_834; // @[Lookup.scala 33:37]
  assign _T_836 = _T_220 ? 1'h0 : _T_835; // @[Lookup.scala 33:37]
  assign _T_837 = _T_218 ? 1'h0 : _T_836; // @[Lookup.scala 33:37]
  assign _T_838 = _T_216 ? 1'h0 : _T_837; // @[Lookup.scala 33:37]
  assign _T_839 = _T_214 ? 1'h0 : _T_838; // @[Lookup.scala 33:37]
  assign _T_840 = _T_212 ? 1'h0 : _T_839; // @[Lookup.scala 33:37]
  assign _T_841 = _T_210 ? 1'h0 : _T_840; // @[Lookup.scala 33:37]
  assign _T_842 = _T_208 ? 1'h0 : _T_841; // @[Lookup.scala 33:37]
  assign _T_843 = _T_206 ? 1'h0 : _T_842; // @[Lookup.scala 33:37]
  assign _T_844 = _T_204 ? 1'h0 : _T_843; // @[Lookup.scala 33:37]
  assign _T_845 = _T_202 ? 1'h0 : _T_844; // @[Lookup.scala 33:37]
  assign _T_846 = _T_200 | _T_845; // @[Lookup.scala 33:37]
  assign _T_847 = _T_198 | _T_846; // @[Lookup.scala 33:37]
  assign _T_848 = _T_196 | _T_847; // @[Lookup.scala 33:37]
  assign _T_849 = _T_194 | _T_848; // @[Lookup.scala 33:37]
  assign _T_850 = _T_192 | _T_849; // @[Lookup.scala 33:37]
  assign _T_851 = _T_190 | _T_850; // @[Lookup.scala 33:37]
  assign _T_852 = _T_188 | _T_851; // @[Lookup.scala 33:37]
  assign _T_853 = _T_186 | _T_852; // @[Lookup.scala 33:37]
  assign _T_854 = _T_184 | _T_853; // @[Lookup.scala 33:37]
  assign _T_855 = _T_182 | _T_854; // @[Lookup.scala 33:37]
  assign _T_856 = _T_180 | _T_855; // @[Lookup.scala 33:37]
  assign _T_857 = _T_178 | _T_856; // @[Lookup.scala 33:37]
  assign _T_858 = _T_176 | _T_857; // @[Lookup.scala 33:37]
  assign _T_859 = _T_174 | _T_858; // @[Lookup.scala 33:37]
  assign _T_860 = _T_172 | _T_859; // @[Lookup.scala 33:37]
  assign _T_861 = _T_170 | _T_860; // @[Lookup.scala 33:37]
  assign _T_862 = _T_168 | _T_861; // @[Lookup.scala 33:37]
  assign _T_863 = _T_166 | _T_862; // @[Lookup.scala 33:37]
  assign _T_864 = _T_164 | _T_863; // @[Lookup.scala 33:37]
  assign _T_865 = _T_162 | _T_864; // @[Lookup.scala 33:37]
  assign _T_866 = _T_160 | _T_865; // @[Lookup.scala 33:37]
  assign _T_867 = _T_158 | _T_866; // @[Lookup.scala 33:37]
  assign _T_868 = _T_156 | _T_867; // @[Lookup.scala 33:37]
  assign _T_869 = _T_154 | _T_868; // @[Lookup.scala 33:37]
  assign _T_870 = _T_152 ? 1'h0 : _T_869; // @[Lookup.scala 33:37]
  assign _T_871 = _T_150 ? 1'h0 : _T_870; // @[Lookup.scala 33:37]
  assign _T_872 = _T_148 | _T_871; // @[Lookup.scala 33:37]
  assign _T_873 = _T_146 | _T_872; // @[Lookup.scala 33:37]
  assign _T_874 = _T_144 | _T_873; // @[Lookup.scala 33:37]
  assign _T_875 = _T_142 | _T_874; // @[Lookup.scala 33:37]
  assign _T_876 = _T_140 ? 1'h0 : _T_875; // @[Lookup.scala 33:37]
  assign _T_877 = _T_138 ? 1'h0 : _T_876; // @[Lookup.scala 33:37]
  assign _T_878 = _T_136 | _T_877; // @[Lookup.scala 33:37]
  assign _T_879 = _T_134 | _T_878; // @[Lookup.scala 33:37]
  assign _T_880 = _T_132 | _T_879; // @[Lookup.scala 33:37]
  assign _T_881 = _T_130 | _T_880; // @[Lookup.scala 33:37]
  assign _T_882 = _T_128 ? 1'h0 : _T_881; // @[Lookup.scala 33:37]
  assign _T_883 = _T_126 ? 1'h0 : _T_882; // @[Lookup.scala 33:37]
  assign _T_884 = _T_124 | _T_883; // @[Lookup.scala 33:37]
  assign _T_885 = _T_122 | _T_884; // @[Lookup.scala 33:37]
  assign _T_886 = _T_120 | _T_885; // @[Lookup.scala 33:37]
  assign _T_887 = _T_118 | _T_886; // @[Lookup.scala 33:37]
  assign _T_888 = _T_116 ? 1'h0 : _T_887; // @[Lookup.scala 33:37]
  assign _T_889 = _T_114 ? 1'h0 : _T_888; // @[Lookup.scala 33:37]
  assign _T_890 = _T_112 ? 1'h0 : _T_889; // @[Lookup.scala 33:37]
  assign _T_891 = _T_110 ? 1'h0 : _T_890; // @[Lookup.scala 33:37]
  assign _T_892 = _T_108 ? 1'h0 : _T_891; // @[Lookup.scala 33:37]
  assign _T_893 = _T_106 ? 1'h0 : _T_892; // @[Lookup.scala 33:37]
  assign _T_894 = _T_104 ? 1'h0 : _T_893; // @[Lookup.scala 33:37]
  assign _T_895 = _T_102 ? 1'h0 : _T_894; // @[Lookup.scala 33:37]
  assign _T_896 = _T_100 | _T_895; // @[Lookup.scala 33:37]
  assign _T_897 = _T_98 | _T_896; // @[Lookup.scala 33:37]
  assign _T_898 = _T_96 | _T_897; // @[Lookup.scala 33:37]
  assign _T_899 = _T_94 | _T_898; // @[Lookup.scala 33:37]
  assign _T_900 = _T_92 | _T_899; // @[Lookup.scala 33:37]
  assign _T_901 = _T_90 | _T_900; // @[Lookup.scala 33:37]
  assign _T_902 = _T_88 | _T_901; // @[Lookup.scala 33:37]
  assign _T_903 = _T_86 | _T_902; // @[Lookup.scala 33:37]
  assign _T_904 = _T_84 | _T_903; // @[Lookup.scala 33:37]
  assign _T_905 = _T_82 | _T_904; // @[Lookup.scala 33:37]
  assign _T_906 = _T_80 | _T_905; // @[Lookup.scala 33:37]
  assign _T_907 = _T_78 | _T_906; // @[Lookup.scala 33:37]
  assign _T_908 = _T_76 | _T_907; // @[Lookup.scala 33:37]
  assign _T_909 = _T_74 | _T_908; // @[Lookup.scala 33:37]
  assign _T_910 = _T_72 | _T_909; // @[Lookup.scala 33:37]
  assign _T_911 = _T_70 | _T_910; // @[Lookup.scala 33:37]
  assign _T_912 = _T_68 | _T_911; // @[Lookup.scala 33:37]
  assign _T_913 = _T_66 | _T_912; // @[Lookup.scala 33:37]
  assign _T_914 = _T_64 | _T_913; // @[Lookup.scala 33:37]
  assign _T_915 = _T_62 | _T_914; // @[Lookup.scala 33:37]
  assign _T_916 = _T_60 | _T_915; // @[Lookup.scala 33:37]
  assign _T_917 = _T_58 | _T_916; // @[Lookup.scala 33:37]
  assign _T_918 = _T_56 | _T_917; // @[Lookup.scala 33:37]
  assign _T_919 = _T_54 | _T_918; // @[Lookup.scala 33:37]
  assign _T_920 = _T_52 ? 1'h0 : _T_919; // @[Lookup.scala 33:37]
  assign _T_921 = _T_50 | _T_920; // @[Lookup.scala 33:37]
  assign _T_922 = _T_48 | _T_921; // @[Lookup.scala 33:37]
  assign _T_923 = _T_46 | _T_922; // @[Lookup.scala 33:37]
  assign _T_924 = _T_44 | _T_923; // @[Lookup.scala 33:37]
  assign _T_925 = _T_42 ? 1'h0 : _T_924; // @[Lookup.scala 33:37]
  assign _T_926 = _T_40 | _T_925; // @[Lookup.scala 33:37]
  assign _T_927 = _T_38 | _T_926; // @[Lookup.scala 33:37]
  assign _T_928 = _T_36 | _T_927; // @[Lookup.scala 33:37]
  assign _T_929 = _T_34 | _T_928; // @[Lookup.scala 33:37]
  assign _T_930 = _T_32 | _T_929; // @[Lookup.scala 33:37]
  assign _T_931 = _T_30 | _T_930; // @[Lookup.scala 33:37]
  assign _T_932 = _T_28 | _T_931; // @[Lookup.scala 33:37]
  assign _T_933 = _T_26 | _T_932; // @[Lookup.scala 33:37]
  assign _T_934 = _T_24 ? 1'h0 : _T_933; // @[Lookup.scala 33:37]
  assign _T_935 = _T_22 | _T_934; // @[Lookup.scala 33:37]
  assign _T_936 = _T_20 | _T_935; // @[Lookup.scala 33:37]
  assign _T_937 = _T_18 | _T_936; // @[Lookup.scala 33:37]
  assign _T_938 = _T_16 | _T_937; // @[Lookup.scala 33:37]
  assign _T_939 = _T_14 | _T_938; // @[Lookup.scala 33:37]
  assign _T_940 = _T_12 | _T_939; // @[Lookup.scala 33:37]
  assign _T_941 = _T_10 | _T_940; // @[Lookup.scala 33:37]
  assign _T_942 = _T_8 | _T_941; // @[Lookup.scala 33:37]
  assign _T_943 = _T_6 ? 1'h0 : _T_942; // @[Lookup.scala 33:37]
  assign _T_944 = _T_4 | _T_943; // @[Lookup.scala 33:37]
  assign _T_1037 = _T_196 | _T_198; // @[Lookup.scala 33:37]
  assign _T_1038 = _T_194 | _T_1037; // @[Lookup.scala 33:37]
  assign _T_1039 = _T_192 | _T_1038; // @[Lookup.scala 33:37]
  assign _T_1040 = _T_190 | _T_1039; // @[Lookup.scala 33:37]
  assign _T_1041 = _T_188 | _T_1040; // @[Lookup.scala 33:37]
  assign _T_1042 = _T_186 | _T_1041; // @[Lookup.scala 33:37]
  assign _T_1043 = _T_184 | _T_1042; // @[Lookup.scala 33:37]
  assign _T_1044 = _T_182 ? 1'h0 : _T_1043; // @[Lookup.scala 33:37]
  assign _T_1045 = _T_180 ? 1'h0 : _T_1044; // @[Lookup.scala 33:37]
  assign _T_1046 = _T_178 ? 1'h0 : _T_1045; // @[Lookup.scala 33:37]
  assign _T_1047 = _T_176 ? 1'h0 : _T_1046; // @[Lookup.scala 33:37]
  assign _T_1048 = _T_174 ? 1'h0 : _T_1047; // @[Lookup.scala 33:37]
  assign _T_1049 = _T_172 ? 1'h0 : _T_1048; // @[Lookup.scala 33:37]
  assign _T_1050 = _T_170 ? 1'h0 : _T_1049; // @[Lookup.scala 33:37]
  assign _T_1051 = _T_168 ? 1'h0 : _T_1050; // @[Lookup.scala 33:37]
  assign _T_1052 = _T_166 ? 1'h0 : _T_1051; // @[Lookup.scala 33:37]
  assign _T_1053 = _T_164 ? 1'h0 : _T_1052; // @[Lookup.scala 33:37]
  assign _T_1054 = _T_162 ? 1'h0 : _T_1053; // @[Lookup.scala 33:37]
  assign _T_1055 = _T_160 | _T_1054; // @[Lookup.scala 33:37]
  assign _T_1056 = _T_158 | _T_1055; // @[Lookup.scala 33:37]
  assign _T_1057 = _T_156 | _T_1056; // @[Lookup.scala 33:37]
  assign _T_1058 = _T_154 | _T_1057; // @[Lookup.scala 33:37]
  assign _T_1059 = _T_152 | _T_1058; // @[Lookup.scala 33:37]
  assign _T_1060 = _T_150 | _T_1059; // @[Lookup.scala 33:37]
  assign _T_1061 = _T_148 | _T_1060; // @[Lookup.scala 33:37]
  assign _T_1062 = _T_146 | _T_1061; // @[Lookup.scala 33:37]
  assign _T_1063 = _T_144 | _T_1062; // @[Lookup.scala 33:37]
  assign _T_1064 = _T_142 | _T_1063; // @[Lookup.scala 33:37]
  assign _T_1065 = _T_140 | _T_1064; // @[Lookup.scala 33:37]
  assign _T_1066 = _T_138 | _T_1065; // @[Lookup.scala 33:37]
  assign _T_1067 = _T_136 | _T_1066; // @[Lookup.scala 33:37]
  assign _T_1068 = _T_134 | _T_1067; // @[Lookup.scala 33:37]
  assign _T_1069 = _T_132 | _T_1068; // @[Lookup.scala 33:37]
  assign _T_1070 = _T_130 | _T_1069; // @[Lookup.scala 33:37]
  assign _T_1071 = _T_128 | _T_1070; // @[Lookup.scala 33:37]
  assign _T_1072 = _T_126 | _T_1071; // @[Lookup.scala 33:37]
  assign _T_1073 = _T_124 | _T_1072; // @[Lookup.scala 33:37]
  assign _T_1074 = _T_122 | _T_1073; // @[Lookup.scala 33:37]
  assign _T_1075 = _T_120 | _T_1074; // @[Lookup.scala 33:37]
  assign _T_1076 = _T_118 | _T_1075; // @[Lookup.scala 33:37]
  assign _T_1077 = _T_116 | _T_1076; // @[Lookup.scala 33:37]
  assign _T_1078 = _T_114 | _T_1077; // @[Lookup.scala 33:37]
  assign _T_1079 = _T_112 ? 1'h0 : _T_1078; // @[Lookup.scala 33:37]
  assign _T_1080 = _T_110 ? 1'h0 : _T_1079; // @[Lookup.scala 33:37]
  assign _T_1081 = _T_108 ? 1'h0 : _T_1080; // @[Lookup.scala 33:37]
  assign _T_1082 = _T_106 ? 1'h0 : _T_1081; // @[Lookup.scala 33:37]
  assign _T_1083 = _T_104 ? 1'h0 : _T_1082; // @[Lookup.scala 33:37]
  assign _T_1084 = _T_102 ? 1'h0 : _T_1083; // @[Lookup.scala 33:37]
  assign _T_1085 = _T_100 ? 1'h0 : _T_1084; // @[Lookup.scala 33:37]
  assign _T_1086 = _T_98 ? 1'h0 : _T_1085; // @[Lookup.scala 33:37]
  assign _T_1087 = _T_96 ? 1'h0 : _T_1086; // @[Lookup.scala 33:37]
  assign _T_1088 = _T_94 ? 1'h0 : _T_1087; // @[Lookup.scala 33:37]
  assign _T_1089 = _T_92 ? 1'h0 : _T_1088; // @[Lookup.scala 33:37]
  assign _T_1090 = _T_90 ? 1'h0 : _T_1089; // @[Lookup.scala 33:37]
  assign _T_1091 = _T_88 ? 1'h0 : _T_1090; // @[Lookup.scala 33:37]
  assign _T_1092 = _T_86 ? 1'h0 : _T_1091; // @[Lookup.scala 33:37]
  assign _T_1093 = _T_84 | _T_1092; // @[Lookup.scala 33:37]
  assign _T_1094 = _T_82 | _T_1093; // @[Lookup.scala 33:37]
  assign _T_1095 = _T_80 | _T_1094; // @[Lookup.scala 33:37]
  assign _T_1096 = _T_78 | _T_1095; // @[Lookup.scala 33:37]
  assign _T_1097 = _T_76 | _T_1096; // @[Lookup.scala 33:37]
  assign _T_1098 = _T_74 | _T_1097; // @[Lookup.scala 33:37]
  assign _T_1099 = _T_72 ? 1'h0 : _T_1098; // @[Lookup.scala 33:37]
  assign _T_1100 = _T_70 ? 1'h0 : _T_1099; // @[Lookup.scala 33:37]
  assign _T_1101 = _T_68 ? 1'h0 : _T_1100; // @[Lookup.scala 33:37]
  assign _T_1102 = _T_66 ? 1'h0 : _T_1101; // @[Lookup.scala 33:37]
  assign _T_1103 = _T_64 ? 1'h0 : _T_1102; // @[Lookup.scala 33:37]
  assign _T_1104 = _T_62 ? 1'h0 : _T_1103; // @[Lookup.scala 33:37]
  assign _T_1105 = _T_60 ? 1'h0 : _T_1104; // @[Lookup.scala 33:37]
  assign _T_1106 = _T_58 ? 1'h0 : _T_1105; // @[Lookup.scala 33:37]
  assign _T_1107 = _T_56 ? 1'h0 : _T_1106; // @[Lookup.scala 33:37]
  assign _T_1108 = _T_54 ? 1'h0 : _T_1107; // @[Lookup.scala 33:37]
  assign _T_1109 = _T_52 ? 1'h0 : _T_1108; // @[Lookup.scala 33:37]
  assign _T_1110 = _T_50 ? 1'h0 : _T_1109; // @[Lookup.scala 33:37]
  assign _T_1111 = _T_48 ? 1'h0 : _T_1110; // @[Lookup.scala 33:37]
  assign _T_1112 = _T_46 ? 1'h0 : _T_1111; // @[Lookup.scala 33:37]
  assign _T_1113 = _T_44 ? 1'h0 : _T_1112; // @[Lookup.scala 33:37]
  assign _T_1114 = _T_42 ? 1'h0 : _T_1113; // @[Lookup.scala 33:37]
  assign _T_1115 = _T_40 | _T_1114; // @[Lookup.scala 33:37]
  assign _T_1116 = _T_38 | _T_1115; // @[Lookup.scala 33:37]
  assign _T_1117 = _T_36 | _T_1116; // @[Lookup.scala 33:37]
  assign _T_1118 = _T_34 | _T_1117; // @[Lookup.scala 33:37]
  assign _T_1119 = _T_32 | _T_1118; // @[Lookup.scala 33:37]
  assign _T_1120 = _T_30 | _T_1119; // @[Lookup.scala 33:37]
  assign _T_1121 = _T_28 | _T_1120; // @[Lookup.scala 33:37]
  assign _T_1122 = _T_26 | _T_1121; // @[Lookup.scala 33:37]
  assign _T_1123 = _T_24 | _T_1122; // @[Lookup.scala 33:37]
  assign _T_1124 = _T_22 | _T_1123; // @[Lookup.scala 33:37]
  assign _T_1125 = _T_20 | _T_1124; // @[Lookup.scala 33:37]
  assign _T_1126 = _T_18 | _T_1125; // @[Lookup.scala 33:37]
  assign _T_1127 = _T_16 | _T_1126; // @[Lookup.scala 33:37]
  assign _T_1128 = _T_14 | _T_1127; // @[Lookup.scala 33:37]
  assign _T_1129 = _T_12 | _T_1128; // @[Lookup.scala 33:37]
  assign _T_1130 = _T_10 | _T_1129; // @[Lookup.scala 33:37]
  assign _T_1131 = _T_8 | _T_1130; // @[Lookup.scala 33:37]
  assign _T_1132 = _T_6 | _T_1131; // @[Lookup.scala 33:37]
  assign _T_1133 = _T_4 ? 1'h0 : _T_1132; // @[Lookup.scala 33:37]
  assign _T_1134 = _T_2 ? 1'h0 : _T_1133; // @[Lookup.scala 33:37]
  assign _T_1215 = _T_218 ? 1'h0 : _T_220; // @[Lookup.scala 33:37]
  assign _T_1216 = _T_216 ? 1'h0 : _T_1215; // @[Lookup.scala 33:37]
  assign _T_1217 = _T_214 ? 1'h0 : _T_1216; // @[Lookup.scala 33:37]
  assign _T_1218 = _T_212 ? 1'h0 : _T_1217; // @[Lookup.scala 33:37]
  assign _T_1219 = _T_210 ? 1'h0 : _T_1218; // @[Lookup.scala 33:37]
  assign _T_1220 = _T_208 ? 1'h0 : _T_1219; // @[Lookup.scala 33:37]
  assign _T_1221 = _T_206 ? 1'h0 : _T_1220; // @[Lookup.scala 33:37]
  assign _T_1222 = _T_204 ? 1'h0 : _T_1221; // @[Lookup.scala 33:37]
  assign _T_1223 = _T_202 ? 1'h0 : _T_1222; // @[Lookup.scala 33:37]
  assign _T_1224 = _T_200 ? 1'h0 : _T_1223; // @[Lookup.scala 33:37]
  assign _T_1225 = _T_198 ? 1'h0 : _T_1224; // @[Lookup.scala 33:37]
  assign _T_1226 = _T_196 ? 1'h0 : _T_1225; // @[Lookup.scala 33:37]
  assign _T_1227 = _T_194 ? 1'h0 : _T_1226; // @[Lookup.scala 33:37]
  assign _T_1228 = _T_192 ? 1'h0 : _T_1227; // @[Lookup.scala 33:37]
  assign _T_1229 = _T_190 ? 1'h0 : _T_1228; // @[Lookup.scala 33:37]
  assign _T_1230 = _T_188 ? 1'h0 : _T_1229; // @[Lookup.scala 33:37]
  assign _T_1231 = _T_186 ? 1'h0 : _T_1230; // @[Lookup.scala 33:37]
  assign _T_1232 = _T_184 ? 1'h0 : _T_1231; // @[Lookup.scala 33:37]
  assign _T_1233 = _T_182 ? 1'h0 : _T_1232; // @[Lookup.scala 33:37]
  assign _T_1234 = _T_180 ? 1'h0 : _T_1233; // @[Lookup.scala 33:37]
  assign _T_1235 = _T_178 ? 1'h0 : _T_1234; // @[Lookup.scala 33:37]
  assign _T_1236 = _T_176 ? 1'h0 : _T_1235; // @[Lookup.scala 33:37]
  assign _T_1237 = _T_174 ? 1'h0 : _T_1236; // @[Lookup.scala 33:37]
  assign _T_1238 = _T_172 ? 1'h0 : _T_1237; // @[Lookup.scala 33:37]
  assign _T_1239 = _T_170 ? 1'h0 : _T_1238; // @[Lookup.scala 33:37]
  assign _T_1240 = _T_168 ? 1'h0 : _T_1239; // @[Lookup.scala 33:37]
  assign _T_1241 = _T_166 ? 1'h0 : _T_1240; // @[Lookup.scala 33:37]
  assign _T_1242 = _T_164 ? 1'h0 : _T_1241; // @[Lookup.scala 33:37]
  assign _T_1243 = _T_162 ? 1'h0 : _T_1242; // @[Lookup.scala 33:37]
  assign _T_1244 = _T_160 ? 1'h0 : _T_1243; // @[Lookup.scala 33:37]
  assign _T_1245 = _T_158 ? 1'h0 : _T_1244; // @[Lookup.scala 33:37]
  assign _T_1246 = _T_156 ? 1'h0 : _T_1245; // @[Lookup.scala 33:37]
  assign _T_1247 = _T_154 ? 1'h0 : _T_1246; // @[Lookup.scala 33:37]
  assign _T_1248 = _T_152 ? 1'h0 : _T_1247; // @[Lookup.scala 33:37]
  assign _T_1249 = _T_150 ? 1'h0 : _T_1248; // @[Lookup.scala 33:37]
  assign _T_1250 = _T_148 ? 1'h0 : _T_1249; // @[Lookup.scala 33:37]
  assign _T_1251 = _T_146 ? 1'h0 : _T_1250; // @[Lookup.scala 33:37]
  assign _T_1252 = _T_144 ? 1'h0 : _T_1251; // @[Lookup.scala 33:37]
  assign _T_1253 = _T_142 ? 1'h0 : _T_1252; // @[Lookup.scala 33:37]
  assign _T_1254 = _T_140 ? 1'h0 : _T_1253; // @[Lookup.scala 33:37]
  assign _T_1255 = _T_138 ? 1'h0 : _T_1254; // @[Lookup.scala 33:37]
  assign _T_1256 = _T_136 ? 1'h0 : _T_1255; // @[Lookup.scala 33:37]
  assign _T_1257 = _T_134 ? 1'h0 : _T_1256; // @[Lookup.scala 33:37]
  assign _T_1258 = _T_132 ? 1'h0 : _T_1257; // @[Lookup.scala 33:37]
  assign _T_1259 = _T_130 ? 1'h0 : _T_1258; // @[Lookup.scala 33:37]
  assign _T_1260 = _T_128 ? 1'h0 : _T_1259; // @[Lookup.scala 33:37]
  assign _T_1261 = _T_126 ? 1'h0 : _T_1260; // @[Lookup.scala 33:37]
  assign _T_1262 = _T_124 ? 1'h0 : _T_1261; // @[Lookup.scala 33:37]
  assign _T_1263 = _T_122 ? 1'h0 : _T_1262; // @[Lookup.scala 33:37]
  assign _T_1264 = _T_120 ? 1'h0 : _T_1263; // @[Lookup.scala 33:37]
  assign _T_1265 = _T_118 ? 1'h0 : _T_1264; // @[Lookup.scala 33:37]
  assign _T_1266 = _T_116 ? 1'h0 : _T_1265; // @[Lookup.scala 33:37]
  assign _T_1267 = _T_114 ? 1'h0 : _T_1266; // @[Lookup.scala 33:37]
  assign _T_1268 = _T_112 | _T_1267; // @[Lookup.scala 33:37]
  assign _T_1269 = _T_110 | _T_1268; // @[Lookup.scala 33:37]
  assign _T_1270 = _T_108 | _T_1269; // @[Lookup.scala 33:37]
  assign _T_1271 = _T_106 | _T_1270; // @[Lookup.scala 33:37]
  assign _T_1272 = _T_104 | _T_1271; // @[Lookup.scala 33:37]
  assign _T_1273 = _T_102 | _T_1272; // @[Lookup.scala 33:37]
  assign _T_1274 = _T_100 | _T_1273; // @[Lookup.scala 33:37]
  assign _T_1275 = _T_98 | _T_1274; // @[Lookup.scala 33:37]
  assign _T_1276 = _T_96 | _T_1275; // @[Lookup.scala 33:37]
  assign _T_1277 = _T_94 | _T_1276; // @[Lookup.scala 33:37]
  assign _T_1278 = _T_92 | _T_1277; // @[Lookup.scala 33:37]
  assign _T_1279 = _T_90 | _T_1278; // @[Lookup.scala 33:37]
  assign _T_1280 = _T_88 | _T_1279; // @[Lookup.scala 33:37]
  assign _T_1281 = _T_86 | _T_1280; // @[Lookup.scala 33:37]
  assign _T_1282 = _T_84 ? 1'h0 : _T_1281; // @[Lookup.scala 33:37]
  assign _T_1283 = _T_82 ? 1'h0 : _T_1282; // @[Lookup.scala 33:37]
  assign _T_1284 = _T_80 ? 1'h0 : _T_1283; // @[Lookup.scala 33:37]
  assign _T_1285 = _T_78 ? 1'h0 : _T_1284; // @[Lookup.scala 33:37]
  assign _T_1286 = _T_76 ? 1'h0 : _T_1285; // @[Lookup.scala 33:37]
  assign _T_1287 = _T_74 ? 1'h0 : _T_1286; // @[Lookup.scala 33:37]
  assign _T_1288 = _T_72 ? 1'h0 : _T_1287; // @[Lookup.scala 33:37]
  assign _T_1289 = _T_70 ? 1'h0 : _T_1288; // @[Lookup.scala 33:37]
  assign _T_1290 = _T_68 ? 1'h0 : _T_1289; // @[Lookup.scala 33:37]
  assign _T_1291 = _T_66 ? 1'h0 : _T_1290; // @[Lookup.scala 33:37]
  assign _T_1292 = _T_64 ? 1'h0 : _T_1291; // @[Lookup.scala 33:37]
  assign _T_1293 = _T_62 ? 1'h0 : _T_1292; // @[Lookup.scala 33:37]
  assign _T_1294 = _T_60 ? 1'h0 : _T_1293; // @[Lookup.scala 33:37]
  assign _T_1295 = _T_58 ? 1'h0 : _T_1294; // @[Lookup.scala 33:37]
  assign _T_1296 = _T_56 ? 1'h0 : _T_1295; // @[Lookup.scala 33:37]
  assign _T_1297 = _T_54 ? 1'h0 : _T_1296; // @[Lookup.scala 33:37]
  assign _T_1298 = _T_52 ? 1'h0 : _T_1297; // @[Lookup.scala 33:37]
  assign _T_1299 = _T_50 ? 1'h0 : _T_1298; // @[Lookup.scala 33:37]
  assign _T_1300 = _T_48 ? 1'h0 : _T_1299; // @[Lookup.scala 33:37]
  assign _T_1301 = _T_46 ? 1'h0 : _T_1300; // @[Lookup.scala 33:37]
  assign _T_1302 = _T_44 ? 1'h0 : _T_1301; // @[Lookup.scala 33:37]
  assign _T_1303 = _T_42 ? 1'h0 : _T_1302; // @[Lookup.scala 33:37]
  assign _T_1304 = _T_40 ? 1'h0 : _T_1303; // @[Lookup.scala 33:37]
  assign _T_1305 = _T_38 ? 1'h0 : _T_1304; // @[Lookup.scala 33:37]
  assign _T_1306 = _T_36 ? 1'h0 : _T_1305; // @[Lookup.scala 33:37]
  assign _T_1307 = _T_34 ? 1'h0 : _T_1306; // @[Lookup.scala 33:37]
  assign _T_1308 = _T_32 ? 1'h0 : _T_1307; // @[Lookup.scala 33:37]
  assign _T_1309 = _T_30 ? 1'h0 : _T_1308; // @[Lookup.scala 33:37]
  assign _T_1310 = _T_28 ? 1'h0 : _T_1309; // @[Lookup.scala 33:37]
  assign _T_1311 = _T_26 ? 1'h0 : _T_1310; // @[Lookup.scala 33:37]
  assign _T_1312 = _T_24 ? 1'h0 : _T_1311; // @[Lookup.scala 33:37]
  assign _T_1313 = _T_22 ? 1'h0 : _T_1312; // @[Lookup.scala 33:37]
  assign _T_1314 = _T_20 ? 1'h0 : _T_1313; // @[Lookup.scala 33:37]
  assign _T_1315 = _T_18 ? 1'h0 : _T_1314; // @[Lookup.scala 33:37]
  assign _T_1316 = _T_16 ? 1'h0 : _T_1315; // @[Lookup.scala 33:37]
  assign _T_1317 = _T_14 ? 1'h0 : _T_1316; // @[Lookup.scala 33:37]
  assign _T_1318 = _T_12 ? 1'h0 : _T_1317; // @[Lookup.scala 33:37]
  assign _T_1319 = _T_10 ? 1'h0 : _T_1318; // @[Lookup.scala 33:37]
  assign _T_1320 = _T_8 ? 1'h0 : _T_1319; // @[Lookup.scala 33:37]
  assign _T_1321 = _T_6 ? 1'h0 : _T_1320; // @[Lookup.scala 33:37]
  assign _T_1322 = _T_4 ? 1'h0 : _T_1321; // @[Lookup.scala 33:37]
  assign _T_1434 = _T_158 ? 1'h0 : _T_160; // @[Lookup.scala 33:37]
  assign _T_1435 = _T_156 | _T_1434; // @[Lookup.scala 33:37]
  assign _T_1436 = _T_154 ? 1'h0 : _T_1435; // @[Lookup.scala 33:37]
  assign _T_1437 = _T_152 | _T_1436; // @[Lookup.scala 33:37]
  assign _T_1438 = _T_150 | _T_1437; // @[Lookup.scala 33:37]
  assign _T_1439 = _T_148 | _T_1438; // @[Lookup.scala 33:37]
  assign _T_1440 = _T_146 ? 1'h0 : _T_1439; // @[Lookup.scala 33:37]
  assign _T_1441 = _T_144 | _T_1440; // @[Lookup.scala 33:37]
  assign _T_1442 = _T_142 ? 1'h0 : _T_1441; // @[Lookup.scala 33:37]
  assign _T_1443 = _T_140 | _T_1442; // @[Lookup.scala 33:37]
  assign _T_1444 = _T_138 | _T_1443; // @[Lookup.scala 33:37]
  assign _T_1445 = _T_136 | _T_1444; // @[Lookup.scala 33:37]
  assign _T_1446 = _T_134 ? 1'h0 : _T_1445; // @[Lookup.scala 33:37]
  assign _T_1447 = _T_132 | _T_1446; // @[Lookup.scala 33:37]
  assign _T_1448 = _T_130 ? 1'h0 : _T_1447; // @[Lookup.scala 33:37]
  assign _T_1449 = _T_128 | _T_1448; // @[Lookup.scala 33:37]
  assign _T_1450 = _T_126 | _T_1449; // @[Lookup.scala 33:37]
  assign _T_1451 = _T_124 | _T_1450; // @[Lookup.scala 33:37]
  assign _T_1452 = _T_122 ? 1'h0 : _T_1451; // @[Lookup.scala 33:37]
  assign _T_1453 = _T_120 | _T_1452; // @[Lookup.scala 33:37]
  assign _T_1454 = _T_118 ? 1'h0 : _T_1453; // @[Lookup.scala 33:37]
  assign _T_1455 = _T_116 | _T_1454; // @[Lookup.scala 33:37]
  assign _T_1456 = _T_114 | _T_1455; // @[Lookup.scala 33:37]
  assign _T_1457 = _T_112 | _T_1456; // @[Lookup.scala 33:37]
  assign _T_1458 = _T_110 | _T_1457; // @[Lookup.scala 33:37]
  assign _T_1459 = _T_108 | _T_1458; // @[Lookup.scala 33:37]
  assign _T_1460 = _T_106 | _T_1459; // @[Lookup.scala 33:37]
  assign _T_1461 = _T_104 | _T_1460; // @[Lookup.scala 33:37]
  assign _T_1462 = _T_102 | _T_1461; // @[Lookup.scala 33:37]
  assign _T_1463 = _T_100 ? 1'h0 : _T_1462; // @[Lookup.scala 33:37]
  assign _T_1464 = _T_98 ? 1'h0 : _T_1463; // @[Lookup.scala 33:37]
  assign _T_1465 = _T_96 ? 1'h0 : _T_1464; // @[Lookup.scala 33:37]
  assign _T_1466 = _T_94 ? 1'h0 : _T_1465; // @[Lookup.scala 33:37]
  assign _T_1467 = _T_92 ? 1'h0 : _T_1466; // @[Lookup.scala 33:37]
  assign _T_1468 = _T_90 ? 1'h0 : _T_1467; // @[Lookup.scala 33:37]
  assign _T_1469 = _T_88 ? 1'h0 : _T_1468; // @[Lookup.scala 33:37]
  assign _T_1470 = _T_86 ? 1'h0 : _T_1469; // @[Lookup.scala 33:37]
  assign _T_1471 = _T_84 ? 1'h0 : _T_1470; // @[Lookup.scala 33:37]
  assign _T_1472 = _T_82 ? 1'h0 : _T_1471; // @[Lookup.scala 33:37]
  assign _T_1473 = _T_80 ? 1'h0 : _T_1472; // @[Lookup.scala 33:37]
  assign _T_1474 = _T_78 ? 1'h0 : _T_1473; // @[Lookup.scala 33:37]
  assign _T_1475 = _T_76 ? 1'h0 : _T_1474; // @[Lookup.scala 33:37]
  assign _T_1476 = _T_74 ? 1'h0 : _T_1475; // @[Lookup.scala 33:37]
  assign _T_1477 = _T_72 ? 1'h0 : _T_1476; // @[Lookup.scala 33:37]
  assign _T_1478 = _T_70 ? 1'h0 : _T_1477; // @[Lookup.scala 33:37]
  assign _T_1479 = _T_68 ? 1'h0 : _T_1478; // @[Lookup.scala 33:37]
  assign _T_1480 = _T_66 ? 1'h0 : _T_1479; // @[Lookup.scala 33:37]
  assign _T_1481 = _T_64 ? 1'h0 : _T_1480; // @[Lookup.scala 33:37]
  assign _T_1482 = _T_62 ? 1'h0 : _T_1481; // @[Lookup.scala 33:37]
  assign _T_1483 = _T_60 | _T_1482; // @[Lookup.scala 33:37]
  assign _T_1484 = _T_58 ? 1'h0 : _T_1483; // @[Lookup.scala 33:37]
  assign _T_1485 = _T_56 ? 1'h0 : _T_1484; // @[Lookup.scala 33:37]
  assign _T_1486 = _T_54 ? 1'h0 : _T_1485; // @[Lookup.scala 33:37]
  assign _T_1487 = _T_52 | _T_1486; // @[Lookup.scala 33:37]
  assign _T_1488 = _T_50 | _T_1487; // @[Lookup.scala 33:37]
  assign _T_1489 = _T_48 ? 1'h0 : _T_1488; // @[Lookup.scala 33:37]
  assign _T_1490 = _T_46 ? 1'h0 : _T_1489; // @[Lookup.scala 33:37]
  assign _T_1491 = _T_44 ? 1'h0 : _T_1490; // @[Lookup.scala 33:37]
  assign _T_1492 = _T_42 | _T_1491; // @[Lookup.scala 33:37]
  assign _T_1493 = _T_40 | _T_1492; // @[Lookup.scala 33:37]
  assign _T_1494 = _T_38 | _T_1493; // @[Lookup.scala 33:37]
  assign _T_1495 = _T_36 ? 1'h0 : _T_1494; // @[Lookup.scala 33:37]
  assign _T_1496 = _T_34 ? 1'h0 : _T_1495; // @[Lookup.scala 33:37]
  assign _T_1497 = _T_32 ? 1'h0 : _T_1496; // @[Lookup.scala 33:37]
  assign _T_1498 = _T_30 ? 1'h0 : _T_1497; // @[Lookup.scala 33:37]
  assign _T_1499 = _T_28 ? 1'h0 : _T_1498; // @[Lookup.scala 33:37]
  assign _T_1500 = _T_26 ? 1'h0 : _T_1499; // @[Lookup.scala 33:37]
  assign _T_1501 = _T_24 | _T_1500; // @[Lookup.scala 33:37]
  assign _T_1502 = _T_22 | _T_1501; // @[Lookup.scala 33:37]
  assign _T_1503 = _T_20 | _T_1502; // @[Lookup.scala 33:37]
  assign _T_1504 = _T_18 ? 1'h0 : _T_1503; // @[Lookup.scala 33:37]
  assign _T_1505 = _T_16 ? 1'h0 : _T_1504; // @[Lookup.scala 33:37]
  assign _T_1506 = _T_14 ? 1'h0 : _T_1505; // @[Lookup.scala 33:37]
  assign _T_1507 = _T_12 ? 1'h0 : _T_1506; // @[Lookup.scala 33:37]
  assign _T_1508 = _T_10 ? 1'h0 : _T_1507; // @[Lookup.scala 33:37]
  assign _T_1509 = _T_8 ? 1'h0 : _T_1508; // @[Lookup.scala 33:37]
  assign _T_1510 = _T_6 | _T_1509; // @[Lookup.scala 33:37]
  assign _T_1511 = _T_4 ? 1'h0 : _T_1510; // @[Lookup.scala 33:37]
  assign _T_1517 = _T_370 | _T_372; // @[Lookup.scala 33:37]
  assign _T_1518 = _T_368 | _T_1517; // @[Lookup.scala 33:37]
  assign _T_1519 = _T_366 ? 1'h0 : _T_1518; // @[Lookup.scala 33:37]
  assign _T_1520 = _T_364 ? 1'h0 : _T_1519; // @[Lookup.scala 33:37]
  assign _T_1521 = _T_362 ? 1'h0 : _T_1520; // @[Lookup.scala 33:37]
  assign _T_1522 = _T_360 | _T_1521; // @[Lookup.scala 33:37]
  assign _T_1523 = _T_358 ? 1'h0 : _T_1522; // @[Lookup.scala 33:37]
  assign _T_1524 = _T_356 ? 1'h0 : _T_1523; // @[Lookup.scala 33:37]
  assign _T_1525 = _T_354 ? 1'h0 : _T_1524; // @[Lookup.scala 33:37]
  assign _T_1526 = _T_352 ? 1'h0 : _T_1525; // @[Lookup.scala 33:37]
  assign _T_1527 = _T_350 ? 1'h0 : _T_1526; // @[Lookup.scala 33:37]
  assign _T_1528 = _T_348 ? 1'h0 : _T_1527; // @[Lookup.scala 33:37]
  assign _T_1529 = _T_346 | _T_1528; // @[Lookup.scala 33:37]
  assign _T_1530 = _T_344 | _T_1529; // @[Lookup.scala 33:37]
  assign _T_1531 = _T_342 | _T_1530; // @[Lookup.scala 33:37]
  assign _T_1532 = _T_340 ? 1'h0 : _T_1531; // @[Lookup.scala 33:37]
  assign _T_1533 = _T_338 ? 1'h0 : _T_1532; // @[Lookup.scala 33:37]
  assign _T_1534 = _T_336 ? 1'h0 : _T_1533; // @[Lookup.scala 33:37]
  assign _T_1535 = _T_334 | _T_1534; // @[Lookup.scala 33:37]
  assign _T_1536 = _T_332 ? 1'h0 : _T_1535; // @[Lookup.scala 33:37]
  assign _T_1537 = _T_330 ? 1'h0 : _T_1536; // @[Lookup.scala 33:37]
  assign _T_1538 = _T_328 ? 1'h0 : _T_1537; // @[Lookup.scala 33:37]
  assign _T_1539 = _T_326 ? 1'h0 : _T_1538; // @[Lookup.scala 33:37]
  assign _T_1540 = _T_324 ? 1'h0 : _T_1539; // @[Lookup.scala 33:37]
  assign _T_1541 = _T_322 ? 1'h0 : _T_1540; // @[Lookup.scala 33:37]
  assign _T_1542 = _T_320 | _T_1541; // @[Lookup.scala 33:37]
  assign _T_1543 = _T_318 | _T_1542; // @[Lookup.scala 33:37]
  assign _T_1544 = _T_316 | _T_1543; // @[Lookup.scala 33:37]
  assign _T_1545 = _T_314 ? 1'h0 : _T_1544; // @[Lookup.scala 33:37]
  assign _T_1546 = _T_312 ? 1'h0 : _T_1545; // @[Lookup.scala 33:37]
  assign _T_1547 = _T_310 ? 1'h0 : _T_1546; // @[Lookup.scala 33:37]
  assign _T_1548 = _T_308 | _T_1547; // @[Lookup.scala 33:37]
  assign _T_1549 = _T_306 ? 1'h0 : _T_1548; // @[Lookup.scala 33:37]
  assign _T_1550 = _T_304 ? 1'h0 : _T_1549; // @[Lookup.scala 33:37]
  assign _T_1551 = _T_302 ? 1'h0 : _T_1550; // @[Lookup.scala 33:37]
  assign _T_1552 = _T_300 | _T_1551; // @[Lookup.scala 33:37]
  assign _T_1553 = _T_298 ? 1'h0 : _T_1552; // @[Lookup.scala 33:37]
  assign _T_1554 = _T_296 | _T_1553; // @[Lookup.scala 33:37]
  assign _T_1555 = _T_294 ? 1'h0 : _T_1554; // @[Lookup.scala 33:37]
  assign _T_1556 = _T_292 ? 1'h0 : _T_1555; // @[Lookup.scala 33:37]
  assign _T_1557 = _T_290 ? 1'h0 : _T_1556; // @[Lookup.scala 33:37]
  assign _T_1558 = _T_288 | _T_1557; // @[Lookup.scala 33:37]
  assign _T_1559 = _T_286 | _T_1558; // @[Lookup.scala 33:37]
  assign _T_1560 = _T_284 | _T_1559; // @[Lookup.scala 33:37]
  assign _T_1561 = _T_282 ? 1'h0 : _T_1560; // @[Lookup.scala 33:37]
  assign _T_1562 = _T_280 | _T_1561; // @[Lookup.scala 33:37]
  assign _T_1563 = _T_278 | _T_1562; // @[Lookup.scala 33:37]
  assign _T_1564 = _T_276 | _T_1563; // @[Lookup.scala 33:37]
  assign _T_1565 = _T_274 ? 1'h0 : _T_1564; // @[Lookup.scala 33:37]
  assign _T_1566 = _T_272 | _T_1565; // @[Lookup.scala 33:37]
  assign _T_1567 = _T_270 | _T_1566; // @[Lookup.scala 33:37]
  assign _T_1568 = _T_268 | _T_1567; // @[Lookup.scala 33:37]
  assign _T_1569 = _T_266 ? 1'h0 : _T_1568; // @[Lookup.scala 33:37]
  assign _T_1570 = _T_264 | _T_1569; // @[Lookup.scala 33:37]
  assign _T_1571 = _T_262 | _T_1570; // @[Lookup.scala 33:37]
  assign _T_1572 = _T_260 | _T_1571; // @[Lookup.scala 33:37]
  assign _T_1573 = _T_258 ? 1'h0 : _T_1572; // @[Lookup.scala 33:37]
  assign _T_1574 = _T_256 ? 1'h0 : _T_1573; // @[Lookup.scala 33:37]
  assign _T_1575 = _T_254 | _T_1574; // @[Lookup.scala 33:37]
  assign _T_1576 = _T_252 ? 1'h0 : _T_1575; // @[Lookup.scala 33:37]
  assign _T_1577 = _T_250 | _T_1576; // @[Lookup.scala 33:37]
  assign _T_1578 = _T_248 ? 1'h0 : _T_1577; // @[Lookup.scala 33:37]
  assign _T_1579 = _T_246 ? 1'h0 : _T_1578; // @[Lookup.scala 33:37]
  assign _T_1580 = _T_244 | _T_1579; // @[Lookup.scala 33:37]
  assign _T_1581 = _T_242 ? 1'h0 : _T_1580; // @[Lookup.scala 33:37]
  assign _T_1582 = _T_240 | _T_1581; // @[Lookup.scala 33:37]
  assign _T_1583 = _T_238 ? 1'h0 : _T_1582; // @[Lookup.scala 33:37]
  assign _T_1584 = _T_236 ? 1'h0 : _T_1583; // @[Lookup.scala 33:37]
  assign _T_1585 = _T_234 | _T_1584; // @[Lookup.scala 33:37]
  assign _T_1586 = _T_232 ? 1'h0 : _T_1585; // @[Lookup.scala 33:37]
  assign _T_1587 = _T_230 | _T_1586; // @[Lookup.scala 33:37]
  assign _T_1588 = _T_228 ? 1'h0 : _T_1587; // @[Lookup.scala 33:37]
  assign _T_1589 = _T_226 ? 1'h0 : _T_1588; // @[Lookup.scala 33:37]
  assign _T_1590 = _T_224 | _T_1589; // @[Lookup.scala 33:37]
  assign _T_1591 = _T_222 | _T_1590; // @[Lookup.scala 33:37]
  assign _T_1592 = _T_220 ? 1'h0 : _T_1591; // @[Lookup.scala 33:37]
  assign _T_1593 = _T_218 ? 1'h0 : _T_1592; // @[Lookup.scala 33:37]
  assign _T_1594 = _T_216 ? 1'h0 : _T_1593; // @[Lookup.scala 33:37]
  assign _T_1595 = _T_214 | _T_1594; // @[Lookup.scala 33:37]
  assign _T_1596 = _T_212 | _T_1595; // @[Lookup.scala 33:37]
  assign _T_1597 = _T_210 ? 1'h0 : _T_1596; // @[Lookup.scala 33:37]
  assign _T_1598 = _T_208 ? 1'h0 : _T_1597; // @[Lookup.scala 33:37]
  assign _T_1599 = _T_206 ? 1'h0 : _T_1598; // @[Lookup.scala 33:37]
  assign _T_1600 = _T_204 ? 1'h0 : _T_1599; // @[Lookup.scala 33:37]
  assign _T_1601 = _T_202 ? 1'h0 : _T_1600; // @[Lookup.scala 33:37]
  assign _T_1602 = _T_200 | _T_1601; // @[Lookup.scala 33:37]
  assign _T_1603 = _T_198 ? 1'h0 : _T_1602; // @[Lookup.scala 33:37]
  assign _T_1604 = _T_196 ? 1'h0 : _T_1603; // @[Lookup.scala 33:37]
  assign _T_1605 = _T_194 ? 1'h0 : _T_1604; // @[Lookup.scala 33:37]
  assign _T_1606 = _T_192 ? 1'h0 : _T_1605; // @[Lookup.scala 33:37]
  assign _T_1607 = _T_190 | _T_1606; // @[Lookup.scala 33:37]
  assign _T_1608 = _T_188 | _T_1607; // @[Lookup.scala 33:37]
  assign _T_1609 = _T_186 | _T_1608; // @[Lookup.scala 33:37]
  assign _T_1610 = _T_184 | _T_1609; // @[Lookup.scala 33:37]
  assign _T_1611 = _T_182 ? 1'h0 : _T_1610; // @[Lookup.scala 33:37]
  assign _T_1612 = _T_180 ? 1'h0 : _T_1611; // @[Lookup.scala 33:37]
  assign _T_1613 = _T_178 ? 1'h0 : _T_1612; // @[Lookup.scala 33:37]
  assign _T_1614 = _T_176 ? 1'h0 : _T_1613; // @[Lookup.scala 33:37]
  assign _T_1615 = _T_174 ? 1'h0 : _T_1614; // @[Lookup.scala 33:37]
  assign _T_1616 = _T_172 ? 1'h0 : _T_1615; // @[Lookup.scala 33:37]
  assign _T_1617 = _T_170 | _T_1616; // @[Lookup.scala 33:37]
  assign _T_1618 = _T_168 | _T_1617; // @[Lookup.scala 33:37]
  assign _T_1619 = _T_166 | _T_1618; // @[Lookup.scala 33:37]
  assign _T_1620 = _T_164 | _T_1619; // @[Lookup.scala 33:37]
  assign _T_1621 = _T_162 | _T_1620; // @[Lookup.scala 33:37]
  assign _T_1622 = _T_160 ? 1'h0 : _T_1621; // @[Lookup.scala 33:37]
  assign _T_1623 = _T_158 ? 1'h0 : _T_1622; // @[Lookup.scala 33:37]
  assign _T_1624 = _T_156 ? 1'h0 : _T_1623; // @[Lookup.scala 33:37]
  assign _T_1625 = _T_154 ? 1'h0 : _T_1624; // @[Lookup.scala 33:37]
  assign _T_1626 = _T_152 ? 1'h0 : _T_1625; // @[Lookup.scala 33:37]
  assign _T_1627 = _T_150 ? 1'h0 : _T_1626; // @[Lookup.scala 33:37]
  assign _T_1628 = _T_148 | _T_1627; // @[Lookup.scala 33:37]
  assign _T_1629 = _T_146 | _T_1628; // @[Lookup.scala 33:37]
  assign _T_1630 = _T_144 | _T_1629; // @[Lookup.scala 33:37]
  assign _T_1631 = _T_142 | _T_1630; // @[Lookup.scala 33:37]
  assign _T_1632 = _T_140 | _T_1631; // @[Lookup.scala 33:37]
  assign _T_1633 = _T_138 | _T_1632; // @[Lookup.scala 33:37]
  assign _T_1634 = _T_136 ? 1'h0 : _T_1633; // @[Lookup.scala 33:37]
  assign _T_1635 = _T_134 ? 1'h0 : _T_1634; // @[Lookup.scala 33:37]
  assign _T_1636 = _T_132 ? 1'h0 : _T_1635; // @[Lookup.scala 33:37]
  assign _T_1637 = _T_130 ? 1'h0 : _T_1636; // @[Lookup.scala 33:37]
  assign _T_1638 = _T_128 ? 1'h0 : _T_1637; // @[Lookup.scala 33:37]
  assign _T_1639 = _T_126 ? 1'h0 : _T_1638; // @[Lookup.scala 33:37]
  assign _T_1640 = _T_124 | _T_1639; // @[Lookup.scala 33:37]
  assign _T_1641 = _T_122 | _T_1640; // @[Lookup.scala 33:37]
  assign _T_1642 = _T_120 | _T_1641; // @[Lookup.scala 33:37]
  assign _T_1643 = _T_118 | _T_1642; // @[Lookup.scala 33:37]
  assign _T_1644 = _T_116 | _T_1643; // @[Lookup.scala 33:37]
  assign _T_1645 = _T_114 | _T_1644; // @[Lookup.scala 33:37]
  assign _T_1646 = _T_112 | _T_1645; // @[Lookup.scala 33:37]
  assign _T_1647 = _T_110 ? 1'h0 : _T_1646; // @[Lookup.scala 33:37]
  assign _T_1648 = _T_108 ? 1'h0 : _T_1647; // @[Lookup.scala 33:37]
  assign _T_1649 = _T_106 | _T_1648; // @[Lookup.scala 33:37]
  assign _T_1650 = _T_104 ? 1'h0 : _T_1649; // @[Lookup.scala 33:37]
  assign _T_1651 = _T_102 ? 1'h0 : _T_1650; // @[Lookup.scala 33:37]
  assign _T_1652 = _T_100 ? 1'h0 : _T_1651; // @[Lookup.scala 33:37]
  assign _T_1653 = _T_98 ? 1'h0 : _T_1652; // @[Lookup.scala 33:37]
  assign _T_1654 = _T_96 ? 1'h0 : _T_1653; // @[Lookup.scala 33:37]
  assign _T_1655 = _T_94 ? 1'h0 : _T_1654; // @[Lookup.scala 33:37]
  assign _T_1656 = _T_92 | _T_1655; // @[Lookup.scala 33:37]
  assign _T_1657 = _T_90 | _T_1656; // @[Lookup.scala 33:37]
  assign _T_1658 = _T_88 | _T_1657; // @[Lookup.scala 33:37]
  assign _T_1659 = _T_86 | _T_1658; // @[Lookup.scala 33:37]
  assign _T_1660 = _T_84 ? 1'h0 : _T_1659; // @[Lookup.scala 33:37]
  assign _T_1661 = _T_82 ? 1'h0 : _T_1660; // @[Lookup.scala 33:37]
  assign _T_1662 = _T_80 ? 1'h0 : _T_1661; // @[Lookup.scala 33:37]
  assign _T_1663 = _T_78 | _T_1662; // @[Lookup.scala 33:37]
  assign _T_1664 = _T_76 | _T_1663; // @[Lookup.scala 33:37]
  assign _T_1665 = _T_74 | _T_1664; // @[Lookup.scala 33:37]
  assign _T_1666 = _T_72 ? 1'h0 : _T_1665; // @[Lookup.scala 33:37]
  assign _T_1667 = _T_70 ? 1'h0 : _T_1666; // @[Lookup.scala 33:37]
  assign _T_1668 = _T_68 ? 1'h0 : _T_1667; // @[Lookup.scala 33:37]
  assign _T_1669 = _T_66 | _T_1668; // @[Lookup.scala 33:37]
  assign _T_1670 = _T_64 | _T_1669; // @[Lookup.scala 33:37]
  assign _T_1671 = _T_62 | _T_1670; // @[Lookup.scala 33:37]
  assign _T_1672 = _T_60 ? 1'h0 : _T_1671; // @[Lookup.scala 33:37]
  assign _T_1673 = _T_58 ? 1'h0 : _T_1672; // @[Lookup.scala 33:37]
  assign _T_1674 = _T_56 ? 1'h0 : _T_1673; // @[Lookup.scala 33:37]
  assign _T_1675 = _T_54 ? 1'h0 : _T_1674; // @[Lookup.scala 33:37]
  assign _T_1676 = _T_52 ? 1'h0 : _T_1675; // @[Lookup.scala 33:37]
  assign _T_1677 = _T_50 | _T_1676; // @[Lookup.scala 33:37]
  assign _T_1678 = _T_48 | _T_1677; // @[Lookup.scala 33:37]
  assign _T_1679 = _T_46 | _T_1678; // @[Lookup.scala 33:37]
  assign _T_1680 = _T_44 | _T_1679; // @[Lookup.scala 33:37]
  assign _T_1681 = _T_42 | _T_1680; // @[Lookup.scala 33:37]
  assign _T_1682 = _T_40 ? 1'h0 : _T_1681; // @[Lookup.scala 33:37]
  assign _T_1683 = _T_38 ? 1'h0 : _T_1682; // @[Lookup.scala 33:37]
  assign _T_1684 = _T_36 ? 1'h0 : _T_1683; // @[Lookup.scala 33:37]
  assign _T_1685 = _T_34 ? 1'h0 : _T_1684; // @[Lookup.scala 33:37]
  assign _T_1686 = _T_32 ? 1'h0 : _T_1685; // @[Lookup.scala 33:37]
  assign _T_1687 = _T_30 ? 1'h0 : _T_1686; // @[Lookup.scala 33:37]
  assign _T_1688 = _T_28 ? 1'h0 : _T_1687; // @[Lookup.scala 33:37]
  assign _T_1689 = _T_26 ? 1'h0 : _T_1688; // @[Lookup.scala 33:37]
  assign _T_1690 = _T_24 ? 1'h0 : _T_1689; // @[Lookup.scala 33:37]
  assign _T_1691 = _T_22 | _T_1690; // @[Lookup.scala 33:37]
  assign _T_1692 = _T_20 | _T_1691; // @[Lookup.scala 33:37]
  assign _T_1693 = _T_18 | _T_1692; // @[Lookup.scala 33:37]
  assign _T_1694 = _T_16 | _T_1693; // @[Lookup.scala 33:37]
  assign _T_1695 = _T_14 | _T_1694; // @[Lookup.scala 33:37]
  assign _T_1696 = _T_12 | _T_1695; // @[Lookup.scala 33:37]
  assign _T_1697 = _T_10 | _T_1696; // @[Lookup.scala 33:37]
  assign _T_1698 = _T_8 | _T_1697; // @[Lookup.scala 33:37]
  assign _T_1699 = _T_6 | _T_1698; // @[Lookup.scala 33:37]
  assign _T_1700 = _T_4 ? 1'h0 : _T_1699; // @[Lookup.scala 33:37]
  assign _T_1722 = 5'h3 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1723 = _T_1722 ? io_finst_inst[4:0] : 5'h0; // @[Mux.scala 80:57]
  assign _T_1725 = 5'hb == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1726 = _T_1725 ? io_finst_inst[4:0] : _T_1723; // @[Mux.scala 80:57]
  assign _T_1727 = 5'hc == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1728 = _T_1727 ? io_finst_inst[4:0] : _T_1726; // @[Mux.scala 80:57]
  assign _T_1729 = 5'hd == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1730 = _T_1729 ? io_finst_inst[4:0] : _T_1728; // @[Mux.scala 80:57]
  assign _T_1731 = 5'he == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1732 = _T_1731 ? io_finst_inst[4:0] : _T_1730; // @[Mux.scala 80:57]
  assign _T_1733 = 5'h1 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1734 = _T_1733 ? io_finst_inst[4:0] : _T_1732; // @[Mux.scala 80:57]
  assign _T_1735 = 5'h2 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1736 = _T_1735 ? io_finst_inst[4:0] : _T_1734; // @[Mux.scala 80:57]
  assign _T_1737 = 5'ha == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1738 = _T_1737 ? io_finst_inst[4:0] : _T_1736; // @[Mux.scala 80:57]
  assign _T_1739 = 5'h8 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1740 = _T_1739 ? io_finst_inst[4:0] : _T_1738; // @[Mux.scala 80:57]
  assign _T_1741 = 5'h9 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1742 = _T_1741 ? io_finst_inst[4:0] : _T_1740; // @[Mux.scala 80:57]
  assign _T_1744 = _T_1741 ? io_finst_inst[4:0] : _T_1742; // @[Mux.scala 80:57]
  assign _T_1745 = 5'h6 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1746 = _T_1745 ? io_finst_inst[4:0] : _T_1744; // @[Mux.scala 80:57]
  assign _T_1747 = 5'h11 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1748 = _T_1747 ? io_finst_inst[4:0] : _T_1746; // @[Mux.scala 80:57]
  assign _T_1749 = 5'h12 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1750 = _T_1749 ? io_finst_inst[4:0] : _T_1748; // @[Mux.scala 80:57]
  assign _T_1751 = 5'h13 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1752 = _T_1751 ? io_finst_inst[4:0] : _T_1750; // @[Mux.scala 80:57]
  assign _T_1753 = 5'h10 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1754 = _T_1753 ? io_finst_inst[4:0] : _T_1752; // @[Mux.scala 80:57]
  assign _T_1755 = 5'h15 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1756 = _T_1755 ? io_finst_inst[4:0] : _T_1754; // @[Mux.scala 80:57]
  assign _T_1757 = 5'h16 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1758 = _T_1757 ? io_finst_inst[4:0] : _T_1756; // @[Mux.scala 80:57]
  assign _T_1759 = 5'h17 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1760 = _T_1759 ? io_finst_inst[4:0] : _T_1758; // @[Mux.scala 80:57]
  assign _T_1761 = 5'h14 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1783 = 5'h1c == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1784 = _T_1783 ? io_finst_inst[9:5] : 5'h0; // @[Mux.scala 80:57]
  assign _T_1787 = _T_1725 ? io_finst_inst[9:5] : _T_1784; // @[Mux.scala 80:57]
  assign _T_1789 = _T_1727 ? io_finst_inst[9:5] : _T_1787; // @[Mux.scala 80:57]
  assign _T_1791 = _T_1729 ? io_finst_inst[9:5] : _T_1789; // @[Mux.scala 80:57]
  assign _T_1793 = _T_1731 ? io_finst_inst[9:5] : _T_1791; // @[Mux.scala 80:57]
  assign _T_1795 = _T_1733 ? io_finst_inst[9:5] : _T_1793; // @[Mux.scala 80:57]
  assign _T_1797 = _T_1735 ? io_finst_inst[9:5] : _T_1795; // @[Mux.scala 80:57]
  assign _T_1799 = _T_1741 ? io_finst_inst[9:5] : _T_1797; // @[Mux.scala 80:57]
  assign _T_1801 = _T_1739 ? io_finst_inst[9:5] : _T_1799; // @[Mux.scala 80:57]
  assign _T_1802 = 5'h4 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1803 = _T_1802 ? io_finst_inst[9:5] : _T_1801; // @[Mux.scala 80:57]
  assign _T_1804 = 5'h5 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1805 = _T_1804 ? io_finst_inst[9:5] : _T_1803; // @[Mux.scala 80:57]
  assign _T_1807 = _T_1745 ? io_finst_inst[9:5] : _T_1805; // @[Mux.scala 80:57]
  assign _T_1809 = _T_1747 ? io_finst_inst[9:5] : _T_1807; // @[Mux.scala 80:57]
  assign _T_1811 = _T_1749 ? io_finst_inst[9:5] : _T_1809; // @[Mux.scala 80:57]
  assign _T_1813 = _T_1751 ? io_finst_inst[9:5] : _T_1811; // @[Mux.scala 80:57]
  assign _T_1815 = _T_1753 ? io_finst_inst[9:5] : _T_1813; // @[Mux.scala 80:57]
  assign _T_1817 = _T_1755 ? io_finst_inst[9:5] : _T_1815; // @[Mux.scala 80:57]
  assign _T_1819 = _T_1757 ? io_finst_inst[9:5] : _T_1817; // @[Mux.scala 80:57]
  assign _T_1821 = _T_1759 ? io_finst_inst[9:5] : _T_1819; // @[Mux.scala 80:57]
  assign _T_1840 = _T_1733 ? io_finst_inst[20:16] : 5'h0; // @[Mux.scala 80:57]
  assign _T_1843 = _T_1741 ? io_finst_inst[20:16] : _T_1840; // @[Mux.scala 80:57]
  assign _T_1845 = _T_1745 ? io_finst_inst[20:16] : _T_1843; // @[Mux.scala 80:57]
  assign _T_1847 = _T_1804 ? io_finst_inst[20:16] : _T_1845; // @[Mux.scala 80:57]
  assign _T_1848 = 5'h1a == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1849 = _T_1848 ? io_finst_inst[4:0] : _T_1847; // @[Mux.scala 80:57]
  assign _T_1851 = _T_1725 ? io_finst_inst[4:0] : _T_1849; // @[Mux.scala 80:57]
  assign _T_1853 = _T_1729 ? io_finst_inst[20:16] : _T_1851; // @[Mux.scala 80:57]
  assign _T_1855 = _T_1731 ? io_finst_inst[20:16] : _T_1853; // @[Mux.scala 80:57]
  assign _T_1857 = _T_1737 ? io_finst_inst[4:0] : _T_1855; // @[Mux.scala 80:57]
  assign _T_1858 = 5'h1b == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1859 = _T_1858 ? io_finst_inst[4:0] : _T_1857; // @[Mux.scala 80:57]
  assign _T_1861 = _T_1755 ? io_finst_inst[14:10] : _T_1859; // @[Mux.scala 80:57]
  assign _T_1863 = _T_1757 ? io_finst_inst[14:10] : _T_1861; // @[Mux.scala 80:57]
  assign _T_1865 = _T_1759 ? io_finst_inst[14:10] : _T_1863; // @[Mux.scala 80:57]
  assign _T_1867 = _T_1749 ? io_finst_inst[20:16] : _T_1865; // @[Mux.scala 80:57]
  assign _T_1879 = {io_finst_inst[23:5],io_finst_inst[30:29]}; // @[Cat.scala 29:58]
  assign _T_1891 = _T_1725 ? io_finst_inst[22:10] : 13'h0; // @[Mux.scala 80:57]
  assign _T_1894 = _T_1735 ? io_finst_inst[22:10] : _T_1891; // @[Mux.scala 80:57]
  assign _T_1896 = _T_1737 ? io_finst_inst[22:5] : {{5'd0}, _T_1894}; // @[Mux.scala 80:57]
  assign _T_1898 = _T_1848 ? io_finst_inst[23:5] : {{1'd0}, _T_1896}; // @[Mux.scala 80:57]
  assign _T_1900 = _T_1802 ? {{13'd0}, io_finst_inst[21:16]} : _T_1898; // @[Mux.scala 80:57]
  assign _T_1902 = _T_1731 ? {{14'd0}, io_finst_inst[14:10]} : _T_1900; // @[Mux.scala 80:57]
  assign _T_1903 = 5'h18 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1904 = _T_1903 ? io_finst_inst[25:0] : {{7'd0}, _T_1902}; // @[Mux.scala 80:57]
  assign _T_1906 = _T_1722 ? {{5'd0}, _T_1879} : _T_1904; // @[Mux.scala 80:57]
  assign _T_1907 = 5'h19 == dinst_itype; // @[Mux.scala 80:60]
  assign _T_1908 = _T_1907 ? {{7'd0}, io_finst_inst[23:5]} : _T_1906; // @[Mux.scala 80:57]
  assign _T_1910 = _T_1858 ? {{7'd0}, io_finst_inst[23:5]} : _T_1908; // @[Mux.scala 80:57]
  assign _T_1912 = _T_1739 ? {{14'd0}, io_finst_inst[21:10]} : _T_1910; // @[Mux.scala 80:57]
  assign _T_1914 = _T_1747 ? {{17'd0}, io_finst_inst[20:12]} : _T_1912; // @[Mux.scala 80:57]
  assign _T_1916 = _T_1751 ? {{17'd0}, io_finst_inst[20:12]} : _T_1914; // @[Mux.scala 80:57]
  assign _T_1918 = _T_1753 ? {{16'd0}, io_finst_inst[21:12]} : _T_1916; // @[Mux.scala 80:57]
  assign _T_1920 = _T_1755 ? {{19'd0}, io_finst_inst[21:15]} : _T_1918; // @[Mux.scala 80:57]
  assign _T_1922 = _T_1757 ? {{19'd0}, io_finst_inst[21:15]} : _T_1920; // @[Mux.scala 80:57]
  assign _T_1924 = _T_1759 ? {{19'd0}, io_finst_inst[21:15]} : _T_1922; // @[Mux.scala 80:57]
  assign _T_1930 = io_finst_inst[22] ? 4'hc : 4'h0; // @[Decode.scala 131:21]
  assign _T_1933 = _T_1733 ? io_finst_inst[15:10] : 6'h0; // @[Mux.scala 80:57]
  assign _T_1936 = _T_1741 ? io_finst_inst[15:10] : _T_1933; // @[Mux.scala 80:57]
  assign _T_1938 = _T_1739 ? {{2'd0}, _T_1930} : _T_1936; // @[Mux.scala 80:57]
  assign _T_1940 = _T_1725 ? io_finst_inst[21:16] : _T_1938; // @[Mux.scala 80:57]
  assign _T_1945 = _T_1729 ? io_finst_inst[11:10] : 2'h0; // @[Mux.scala 80:57]
  assign _T_1948 = _T_1733 ? io_finst_inst[23:22] : _T_1945; // @[Mux.scala 80:57]
  assign _T_1950 = _T_1741 ? io_finst_inst[23:22] : _T_1948; // @[Mux.scala 80:57]
  assign _T_1952 = _T_1739 ? 2'h0 : _T_1950; // @[Mux.scala 80:57]
  assign _T_1960 = _T_1745 ? io_finst_inst[15:12] : 4'h0; // @[Mux.scala 80:57]
  assign _T_1963 = _T_1802 ? io_finst_inst[15:12] : _T_1960; // @[Mux.scala 80:57]
  assign _T_1965 = _T_1804 ? io_finst_inst[15:12] : _T_1963; // @[Mux.scala 80:57]
  assign _T_1971 = _T_1802 ? io_finst_inst[3:0] : 4'h0; // @[Mux.scala 80:57]
  assign _T_1976 = dinst_itype == 5'h12; // @[Decode.scala 164:16]
  assign io_dinst_rd_valid = _T_2 | _T_944; // @[Decode.scala 226:12]
  assign io_dinst_rd_bits = _T_1761 ? io_finst_inst[4:0] : _T_1760; // @[Decode.scala 226:12]
  assign io_dinst_rs1 = _T_1761 ? io_finst_inst[9:5] : _T_1821; // @[Decode.scala 226:12]
  assign io_dinst_rs2 = _T_1761 ? io_finst_inst[4:0] : _T_1867; // @[Decode.scala 226:12]
  assign io_dinst_imm = _T_1761 ? {{14'd0}, io_finst_inst[21:10]} : _T_1924; // @[Decode.scala 226:12]
  assign io_dinst_shift_val_valid = _T_1976 ? io_finst_inst[12] : _T_1134; // @[Decode.scala 226:12]
  assign io_dinst_shift_val_bits = _T_1976 ? {{3'd0}, io_finst_inst[15:13]} : _T_1940; // @[Decode.scala 226:12]
  assign io_dinst_shift_type = _T_1725 ? 2'h3 : _T_1952; // @[Decode.scala 226:12]
  assign io_dinst_cond_valid = _T_2 ? 1'h0 : _T_1322; // @[Decode.scala 226:12]
  assign io_dinst_cond_bits = _T_1907 ? io_finst_inst[3:0] : _T_1965; // @[Decode.scala 226:12]
  assign io_dinst_is32bit = _T_2 ? 1'h0 : _T_1700; // @[Decode.scala 226:12]
  assign io_dinst_itype = _T_2 ? 5'h3 : _T_566; // @[Decode.scala 226:12]
  assign io_dinst_op = _T_2 ? 4'h0 : _T_755; // @[Decode.scala 226:12]
  assign io_dinst_nzcv_valid = _T_2 ? 1'h0 : _T_1511; // @[Decode.scala 226:12]
  assign io_dinst_nzcv_bits = _T_1804 ? io_finst_inst[3:0] : _T_1971; // @[Decode.scala 226:12]
  assign io_dinst_tag = io_finst_tag; // @[Decode.scala 226:12]
  assign io_dinst_inst32_valid = dinst_itype != 5'h0; // @[Decode.scala 226:12]
  assign io_dinst_inst32_bits = io_finst_inst; // @[Decode.scala 226:12]
  assign io_dinst_pc = io_finst_pc; // @[Decode.scala 226:12]
endmodule
