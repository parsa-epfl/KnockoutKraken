
module DevteroFlexTopLevel (
`ifdef DEBUG
    output         dbg_bits_fetch_valid,
    output [4:0]   dbg_bits_fetch_tag,
    output         dbg_bits_issue_valid,
    output [4:0]   dbg_bits_issue_tag,
    output         dbg_bits_issuingMem,
    output         dbg_bits_issuingTransplant,
    output         dbg_bits_commit_valid,
    output [4:0]   dbg_bits_commit_tag,
    output         dbg_bits_transplant_valid,
    output [4:0]   dbg_bits_transplant_tag,
    output [31:0] [31:0] [63:0]  dbg_bits_stateVec_rfile,
    output [31:0] [63:0] dbg_bits_stateVec_regs_PC,
    output [31:0] [3:0] dbg_bits_stateVec_regs_NZCV,
`endif
    input          clock,
    input          reset,
    input  [5:0]   S_AXI_awid,
    input  [6:0]   S_AXI_awaddr,
    input  [7:0]   S_AXI_awlen,
    input  [2:0]   S_AXI_awsize,
    input  [1:0]   S_AXI_awburst,
    input          S_AXI_awlock,
    input  [3:0]   S_AXI_awcache,
    input  [2:0]   S_AXI_awprot,
    input  [3:0]   S_AXI_awqos,
    input          S_AXI_awvalid,
    output         S_AXI_awready,
    input  [511:0] S_AXI_wdata,
    input  [63:0]  S_AXI_wstrb,
    input          S_AXI_wlast,
    input          S_AXI_wvalid,
    output         S_AXI_wready,
    output [5:0]   S_AXI_bid,
    output [1:0]   S_AXI_bresp,
    output         S_AXI_bvalid,
    input          S_AXI_bready,
    input  [5:0]   S_AXI_arid,
    input  [6:0]   S_AXI_araddr,
    input  [7:0]   S_AXI_arlen,
    input  [2:0]   S_AXI_arsize,
    input  [1:0]   S_AXI_arburst,
    input          S_AXI_arlock,
    input  [3:0]   S_AXI_arcache,
    input  [2:0]   S_AXI_arprot,
    input  [3:0]   S_AXI_arqos,
    input          S_AXI_arvalid,
    output         S_AXI_arready,
    output [5:0]   S_AXI_rid,
    output [511:0] S_AXI_rdata,
    output [1:0]   S_AXI_rresp,
    output         S_AXI_rlast,
    output         S_AXI_rvalid,
    input          S_AXI_rready,
    input  [31:0]  S_AXIL_awaddr,
    input  [2:0]   S_AXIL_awprot,
    input          S_AXIL_awvalid,
    output         S_AXIL_awready,
    input  [31:0]  S_AXIL_wdata,
    input  [3:0]   S_AXIL_wstrb,
    input          S_AXIL_wvalid,
    output         S_AXIL_wready,
    output [1:0]   S_AXIL_bresp,
    output         S_AXIL_bvalid,
    input          S_AXIL_bready,
    input  [31:0]  S_AXIL_araddr,
    input  [2:0]   S_AXIL_arprot,
    input          S_AXIL_arvalid,
    output         S_AXIL_arready,
    output [31:0]  S_AXIL_rdata,
    output [1:0]   S_AXIL_rresp,
    output         S_AXIL_rvalid,
    input          S_AXIL_rready,
    output [5:0]   M_AXI_awid,
    output [23:0]  M_AXI_awaddr,
    output [7:0]   M_AXI_awlen,
    output [2:0]   M_AXI_awsize,
    output [1:0]   M_AXI_awburst,
    output         M_AXI_awlock,
    output [3:0]   M_AXI_awcache,
    output [2:0]   M_AXI_awprot,
    output [3:0]   M_AXI_awqos,
    output         M_AXI_awvalid,
    input          M_AXI_awready,
    output [511:0] M_AXI_wdata,
    output [63:0]  M_AXI_wstrb,
    output         M_AXI_wlast,
    output         M_AXI_wvalid,
    input          M_AXI_wready,
    input  [5:0]   M_AXI_bid,
    input  [1:0]   M_AXI_bresp,
    input          M_AXI_bvalid,
    output         M_AXI_bready,
    output [5:0]   M_AXI_arid,
    output [23:0]  M_AXI_araddr,
    output [7:0]   M_AXI_arlen,
    output [2:0]   M_AXI_arsize,
    output [1:0]   M_AXI_arburst,
    output         M_AXI_arlock,
    output [3:0]   M_AXI_arcache,
    output [2:0]   M_AXI_arprot,
    output [3:0]   M_AXI_arqos,
    output         M_AXI_arvalid,
    input          M_AXI_arready,
    input  [5:0]   M_AXI_rid,
    input  [511:0] M_AXI_rdata,
    input  [1:0]   M_AXI_rresp,
    input          M_AXI_rlast,
    input          M_AXI_rvalid,
    output         M_AXI_rready

);
`ifdef DEVTEROFLEX_INSTRUMENTED
    ARMFlexTopInstrumented DevteroFlexInstance (
`else
    ARMFlexTopSimulator DevteroFlexInstance (
`endif
        .clock              (clock        ),
        .reset              (reset        ),
        .S_AXI_aw_awid      (S_AXI_awid   ),
        .S_AXI_aw_awaddr    (S_AXI_awaddr ),
        .S_AXI_aw_awlen     (S_AXI_awlen  ),
        .S_AXI_aw_awsize    (S_AXI_awsize ),
        .S_AXI_aw_awburst   (S_AXI_awburst),
        .S_AXI_aw_awlock    (S_AXI_awlock ),
        .S_AXI_aw_awcache   (S_AXI_awcache),
        .S_AXI_aw_awprot    (S_AXI_awprot ),
        .S_AXI_aw_awqos     (S_AXI_awqos  ),
        .S_AXI_aw_awvalid   (S_AXI_awvalid),
        .S_AXI_aw_awready   (S_AXI_awready),
        .S_AXI_w_wdata      (S_AXI_wdata  ),
        .S_AXI_w_wstrb      (S_AXI_wstrb  ),
        .S_AXI_w_wlast      (S_AXI_wlast  ),
        .S_AXI_w_wvalid     (S_AXI_wvalid ),
        .S_AXI_w_wready     (S_AXI_wready ),
        .S_AXI_b_bid        (S_AXI_bid    ),
        .S_AXI_b_bresp      (S_AXI_bresp  ),
        .S_AXI_b_bvalid     (S_AXI_bvalid ),
        .S_AXI_b_bready     (S_AXI_bready ),
        .S_AXI_ar_arid      (S_AXI_arid   ),
        .S_AXI_ar_araddr    (S_AXI_araddr ),
        .S_AXI_ar_arlen     (S_AXI_arlen  ),
        .S_AXI_ar_arsize    (S_AXI_arsize ),
        .S_AXI_ar_arburst   (S_AXI_arburst),
        .S_AXI_ar_arlock    (S_AXI_arlock ),
        .S_AXI_ar_arcache   (S_AXI_arcache),
        .S_AXI_ar_arprot    (S_AXI_arprot ),
        .S_AXI_ar_arqos     (S_AXI_arqos  ),
        .S_AXI_ar_arvalid   (S_AXI_arvalid),
        .S_AXI_ar_arready   (S_AXI_arready),
        .S_AXI_r_rid        (S_AXI_rid    ),
        .S_AXI_r_rdata      (S_AXI_rdata  ),
        .S_AXI_r_rresp      (S_AXI_rresp  ),
        .S_AXI_r_rlast      (S_AXI_rlast  ),
        .S_AXI_r_rvalid     (S_AXI_rvalid ),
        .S_AXI_r_rready     (S_AXI_rready ),
        .S_AXIL_aw_awaddr   (S_AXIL_awaddr),
        .S_AXIL_aw_awprot   (S_AXIL_awprot),
        .S_AXIL_aw_awvalid  (S_AXIL_awvalid),
        .S_AXIL_aw_awready  (S_AXIL_awready),
        .S_AXIL_w_wdata     (S_AXIL_wdata ),
        .S_AXIL_w_wstrb     (S_AXIL_wstrb ),
        .S_AXIL_w_wvalid    (S_AXIL_wvalid),
        .S_AXIL_w_wready    (S_AXIL_wready),
        .S_AXIL_b_bresp     (S_AXIL_bresp ),
        .S_AXIL_b_bvalid    (S_AXIL_bvalid),
        .S_AXIL_b_bready    (S_AXIL_bready),
        .S_AXIL_ar_araddr   (S_AXIL_araddr),
        .S_AXIL_ar_arprot   (S_AXIL_arprot),
        .S_AXIL_ar_arvalid  (S_AXIL_arvalid),
        .S_AXIL_ar_arready  (S_AXIL_arready),
        .S_AXIL_r_rdata     (S_AXIL_rdata ),
        .S_AXIL_r_rresp     (S_AXIL_rresp ),
        .S_AXIL_r_rvalid    (S_AXIL_rvalid),
        .S_AXIL_r_rready    (S_AXIL_rready),
        .M_AXI_aw_awid      (M_AXI_awid   ),
        .M_AXI_aw_awaddr    (M_AXI_awaddr ),
        .M_AXI_aw_awlen     (M_AXI_awlen  ),
        .M_AXI_aw_awsize    (M_AXI_awsize ),
        .M_AXI_aw_awburst   (M_AXI_awburst),
        .M_AXI_aw_awlock    (M_AXI_awlock ),
        .M_AXI_aw_awcache   (M_AXI_awcache),
        .M_AXI_aw_awprot    (M_AXI_awprot ),
        .M_AXI_aw_awqos     (M_AXI_awqos  ),
        .M_AXI_aw_awvalid   (M_AXI_awvalid),
        .M_AXI_aw_awready   (M_AXI_awready),
        .M_AXI_w_wdata      (M_AXI_wdata  ),
        .M_AXI_w_wstrb      (M_AXI_wstrb  ),
        .M_AXI_w_wlast      (M_AXI_wlast  ),
        .M_AXI_w_wvalid     (M_AXI_wvalid ),
        .M_AXI_w_wready     (M_AXI_wready ),
        .M_AXI_b_bid        (M_AXI_bid    ),
        .M_AXI_b_bresp      (M_AXI_bresp  ),
        .M_AXI_b_bvalid     (M_AXI_bvalid ),
        .M_AXI_b_bready     (M_AXI_bready ),
        .M_AXI_ar_arid      (M_AXI_arid   ),
        .M_AXI_ar_araddr    (M_AXI_araddr ),
        .M_AXI_ar_arlen     (M_AXI_arlen  ),
        .M_AXI_ar_arsize    (M_AXI_arsize ),
        .M_AXI_ar_arburst   (M_AXI_arburst),
        .M_AXI_ar_arlock    (M_AXI_arlock ),
        .M_AXI_ar_arcache   (M_AXI_arcache),
        .M_AXI_ar_arprot    (M_AXI_arprot ),
        .M_AXI_ar_arqos     (M_AXI_arqos  ),
        .M_AXI_ar_arvalid   (M_AXI_arvalid),
        .M_AXI_ar_arready   (M_AXI_arready),
        .M_AXI_r_rid        (M_AXI_rid    ),
        .M_AXI_r_rdata      (M_AXI_rdata  ),
        .M_AXI_r_rresp      (M_AXI_rresp  ),
        .M_AXI_r_rlast      (M_AXI_rlast  ),
        .M_AXI_r_rvalid     (M_AXI_rvalid ),
        .M_AXI_r_rready     (M_AXI_rready ),
`ifdef DEBUG
    .dbg_bits_fetch_valid              (dbg_bits_fetch_valid       ),
    .dbg_bits_fetch_tag                (dbg_bits_fetch_tag),
    .dbg_bits_issue_valid              (dbg_bits_issue_valid),
    .dbg_bits_issue_tag                (dbg_bits_issue_tag),
    .dbg_bits_issuingMem               (dbg_bits_issuingMem),
    .dbg_bits_issuingTransplant        (dbg_bits_issuingTransplant),
    .dbg_bits_commit_valid             (dbg_bits_commit_valid),
    .dbg_bits_commit_tag               (dbg_bits_commit_tag),
    .dbg_bits_transplant_valid         (dbg_bits_transplant_valid),
    .dbg_bits_transplant_tag           (dbg_bits_transplant_tag),
    .dbg_bits_stateVec_0_rfile_0       (dbg_bits_stateVec_rfile[0][0 ]),
    .dbg_bits_stateVec_0_rfile_1       (dbg_bits_stateVec_rfile[0][1 ]),
    .dbg_bits_stateVec_0_rfile_2       (dbg_bits_stateVec_rfile[0][2 ]),
    .dbg_bits_stateVec_0_rfile_3       (dbg_bits_stateVec_rfile[0][3 ]),
    .dbg_bits_stateVec_0_rfile_4       (dbg_bits_stateVec_rfile[0][4 ]),
    .dbg_bits_stateVec_0_rfile_5       (dbg_bits_stateVec_rfile[0][5 ]),
    .dbg_bits_stateVec_0_rfile_6       (dbg_bits_stateVec_rfile[0][6 ]),
    .dbg_bits_stateVec_0_rfile_7       (dbg_bits_stateVec_rfile[0][7 ]),
    .dbg_bits_stateVec_0_rfile_8       (dbg_bits_stateVec_rfile[0][8 ]),
    .dbg_bits_stateVec_0_rfile_9       (dbg_bits_stateVec_rfile[0][9 ]),
    .dbg_bits_stateVec_0_rfile_10      (dbg_bits_stateVec_rfile[0][10]),
    .dbg_bits_stateVec_0_rfile_11      (dbg_bits_stateVec_rfile[0][11]),
    .dbg_bits_stateVec_0_rfile_12      (dbg_bits_stateVec_rfile[0][12]),
    .dbg_bits_stateVec_0_rfile_13      (dbg_bits_stateVec_rfile[0][13]),
    .dbg_bits_stateVec_0_rfile_14      (dbg_bits_stateVec_rfile[0][14]),
    .dbg_bits_stateVec_0_rfile_15      (dbg_bits_stateVec_rfile[0][15]),
    .dbg_bits_stateVec_0_rfile_16      (dbg_bits_stateVec_rfile[0][16]),
    .dbg_bits_stateVec_0_rfile_17      (dbg_bits_stateVec_rfile[0][17]),
    .dbg_bits_stateVec_0_rfile_18      (dbg_bits_stateVec_rfile[0][18]),
    .dbg_bits_stateVec_0_rfile_19      (dbg_bits_stateVec_rfile[0][19]),
    .dbg_bits_stateVec_0_rfile_20      (dbg_bits_stateVec_rfile[0][20]),
    .dbg_bits_stateVec_0_rfile_21      (dbg_bits_stateVec_rfile[0][21]),
    .dbg_bits_stateVec_0_rfile_22      (dbg_bits_stateVec_rfile[0][22]),
    .dbg_bits_stateVec_0_rfile_23      (dbg_bits_stateVec_rfile[0][23]),
    .dbg_bits_stateVec_0_rfile_24      (dbg_bits_stateVec_rfile[0][24]),
    .dbg_bits_stateVec_0_rfile_25      (dbg_bits_stateVec_rfile[0][25]),
    .dbg_bits_stateVec_0_rfile_26      (dbg_bits_stateVec_rfile[0][26]),
    .dbg_bits_stateVec_0_rfile_27      (dbg_bits_stateVec_rfile[0][27]),
    .dbg_bits_stateVec_0_rfile_28      (dbg_bits_stateVec_rfile[0][28]),
    .dbg_bits_stateVec_0_rfile_29      (dbg_bits_stateVec_rfile[0][29]),
    .dbg_bits_stateVec_0_rfile_30      (dbg_bits_stateVec_rfile[0][30]),
    .dbg_bits_stateVec_0_rfile_31      (dbg_bits_stateVec_rfile[0][31]),
    .dbg_bits_stateVec_0_regs_PC       (dbg_bits_stateVec_regs_PC[0]),
    .dbg_bits_stateVec_0_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[0]),
    .dbg_bits_stateVec_1_rfile_0       (dbg_bits_stateVec_rfile[1][0 ]),
    .dbg_bits_stateVec_1_rfile_1       (dbg_bits_stateVec_rfile[1][1 ]),
    .dbg_bits_stateVec_1_rfile_2       (dbg_bits_stateVec_rfile[1][2 ]),
    .dbg_bits_stateVec_1_rfile_3       (dbg_bits_stateVec_rfile[1][3 ]),
    .dbg_bits_stateVec_1_rfile_4       (dbg_bits_stateVec_rfile[1][4 ]),
    .dbg_bits_stateVec_1_rfile_5       (dbg_bits_stateVec_rfile[1][5 ]),
    .dbg_bits_stateVec_1_rfile_6       (dbg_bits_stateVec_rfile[1][6 ]),
    .dbg_bits_stateVec_1_rfile_7       (dbg_bits_stateVec_rfile[1][7 ]),
    .dbg_bits_stateVec_1_rfile_8       (dbg_bits_stateVec_rfile[1][8 ]),
    .dbg_bits_stateVec_1_rfile_9       (dbg_bits_stateVec_rfile[1][9 ]),
    .dbg_bits_stateVec_1_rfile_10      (dbg_bits_stateVec_rfile[1][10]),
    .dbg_bits_stateVec_1_rfile_11      (dbg_bits_stateVec_rfile[1][11]),
    .dbg_bits_stateVec_1_rfile_12      (dbg_bits_stateVec_rfile[1][12]),
    .dbg_bits_stateVec_1_rfile_13      (dbg_bits_stateVec_rfile[1][13]),
    .dbg_bits_stateVec_1_rfile_14      (dbg_bits_stateVec_rfile[1][14]),
    .dbg_bits_stateVec_1_rfile_15      (dbg_bits_stateVec_rfile[1][15]),
    .dbg_bits_stateVec_1_rfile_16      (dbg_bits_stateVec_rfile[1][16]),
    .dbg_bits_stateVec_1_rfile_17      (dbg_bits_stateVec_rfile[1][17]),
    .dbg_bits_stateVec_1_rfile_18      (dbg_bits_stateVec_rfile[1][18]),
    .dbg_bits_stateVec_1_rfile_19      (dbg_bits_stateVec_rfile[1][19]),
    .dbg_bits_stateVec_1_rfile_20      (dbg_bits_stateVec_rfile[1][20]),
    .dbg_bits_stateVec_1_rfile_21      (dbg_bits_stateVec_rfile[1][21]),
    .dbg_bits_stateVec_1_rfile_22      (dbg_bits_stateVec_rfile[1][22]),
    .dbg_bits_stateVec_1_rfile_23      (dbg_bits_stateVec_rfile[1][23]),
    .dbg_bits_stateVec_1_rfile_24      (dbg_bits_stateVec_rfile[1][24]),
    .dbg_bits_stateVec_1_rfile_25      (dbg_bits_stateVec_rfile[1][25]),
    .dbg_bits_stateVec_1_rfile_26      (dbg_bits_stateVec_rfile[1][26]),
    .dbg_bits_stateVec_1_rfile_27      (dbg_bits_stateVec_rfile[1][27]),
    .dbg_bits_stateVec_1_rfile_28      (dbg_bits_stateVec_rfile[1][28]),
    .dbg_bits_stateVec_1_rfile_29      (dbg_bits_stateVec_rfile[1][29]),
    .dbg_bits_stateVec_1_rfile_30      (dbg_bits_stateVec_rfile[1][30]),
    .dbg_bits_stateVec_1_rfile_31      (dbg_bits_stateVec_rfile[1][31]),
    .dbg_bits_stateVec_1_regs_PC       (dbg_bits_stateVec_regs_PC[1]),
    .dbg_bits_stateVec_1_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[1]),
    .dbg_bits_stateVec_2_rfile_0       (dbg_bits_stateVec_rfile[2][0 ]),
    .dbg_bits_stateVec_2_rfile_1       (dbg_bits_stateVec_rfile[2][1 ]),
    .dbg_bits_stateVec_2_rfile_2       (dbg_bits_stateVec_rfile[2][2 ]),
    .dbg_bits_stateVec_2_rfile_3       (dbg_bits_stateVec_rfile[2][3 ]),
    .dbg_bits_stateVec_2_rfile_4       (dbg_bits_stateVec_rfile[2][4 ]),
    .dbg_bits_stateVec_2_rfile_5       (dbg_bits_stateVec_rfile[2][5 ]),
    .dbg_bits_stateVec_2_rfile_6       (dbg_bits_stateVec_rfile[2][6 ]),
    .dbg_bits_stateVec_2_rfile_7       (dbg_bits_stateVec_rfile[2][7 ]),
    .dbg_bits_stateVec_2_rfile_8       (dbg_bits_stateVec_rfile[2][8 ]),
    .dbg_bits_stateVec_2_rfile_9       (dbg_bits_stateVec_rfile[2][9 ]),
    .dbg_bits_stateVec_2_rfile_10      (dbg_bits_stateVec_rfile[2][10]),
    .dbg_bits_stateVec_2_rfile_11      (dbg_bits_stateVec_rfile[2][11]),
    .dbg_bits_stateVec_2_rfile_12      (dbg_bits_stateVec_rfile[2][12]),
    .dbg_bits_stateVec_2_rfile_13      (dbg_bits_stateVec_rfile[2][13]),
    .dbg_bits_stateVec_2_rfile_14      (dbg_bits_stateVec_rfile[2][14]),
    .dbg_bits_stateVec_2_rfile_15      (dbg_bits_stateVec_rfile[2][15]),
    .dbg_bits_stateVec_2_rfile_16      (dbg_bits_stateVec_rfile[2][16]),
    .dbg_bits_stateVec_2_rfile_17      (dbg_bits_stateVec_rfile[2][17]),
    .dbg_bits_stateVec_2_rfile_18      (dbg_bits_stateVec_rfile[2][18]),
    .dbg_bits_stateVec_2_rfile_19      (dbg_bits_stateVec_rfile[2][19]),
    .dbg_bits_stateVec_2_rfile_20      (dbg_bits_stateVec_rfile[2][20]),
    .dbg_bits_stateVec_2_rfile_21      (dbg_bits_stateVec_rfile[2][21]),
    .dbg_bits_stateVec_2_rfile_22      (dbg_bits_stateVec_rfile[2][22]),
    .dbg_bits_stateVec_2_rfile_23      (dbg_bits_stateVec_rfile[2][23]),
    .dbg_bits_stateVec_2_rfile_24      (dbg_bits_stateVec_rfile[2][24]),
    .dbg_bits_stateVec_2_rfile_25      (dbg_bits_stateVec_rfile[2][25]),
    .dbg_bits_stateVec_2_rfile_26      (dbg_bits_stateVec_rfile[2][26]),
    .dbg_bits_stateVec_2_rfile_27      (dbg_bits_stateVec_rfile[2][27]),
    .dbg_bits_stateVec_2_rfile_28      (dbg_bits_stateVec_rfile[2][28]),
    .dbg_bits_stateVec_2_rfile_29      (dbg_bits_stateVec_rfile[2][29]),
    .dbg_bits_stateVec_2_rfile_30      (dbg_bits_stateVec_rfile[2][30]),
    .dbg_bits_stateVec_2_rfile_31      (dbg_bits_stateVec_rfile[2][31]),
    .dbg_bits_stateVec_2_regs_PC       (dbg_bits_stateVec_regs_PC[2]),
    .dbg_bits_stateVec_2_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[2]),
    .dbg_bits_stateVec_3_rfile_0       (dbg_bits_stateVec_rfile[3][0 ]),
    .dbg_bits_stateVec_3_rfile_1       (dbg_bits_stateVec_rfile[3][1 ]),
    .dbg_bits_stateVec_3_rfile_2       (dbg_bits_stateVec_rfile[3][2 ]),
    .dbg_bits_stateVec_3_rfile_3       (dbg_bits_stateVec_rfile[3][3 ]),
    .dbg_bits_stateVec_3_rfile_4       (dbg_bits_stateVec_rfile[3][4 ]),
    .dbg_bits_stateVec_3_rfile_5       (dbg_bits_stateVec_rfile[3][5 ]),
    .dbg_bits_stateVec_3_rfile_6       (dbg_bits_stateVec_rfile[3][6 ]),
    .dbg_bits_stateVec_3_rfile_7       (dbg_bits_stateVec_rfile[3][7 ]),
    .dbg_bits_stateVec_3_rfile_8       (dbg_bits_stateVec_rfile[3][8 ]),
    .dbg_bits_stateVec_3_rfile_9       (dbg_bits_stateVec_rfile[3][9 ]),
    .dbg_bits_stateVec_3_rfile_10      (dbg_bits_stateVec_rfile[3][10]),
    .dbg_bits_stateVec_3_rfile_11      (dbg_bits_stateVec_rfile[3][11]),
    .dbg_bits_stateVec_3_rfile_12      (dbg_bits_stateVec_rfile[3][12]),
    .dbg_bits_stateVec_3_rfile_13      (dbg_bits_stateVec_rfile[3][13]),
    .dbg_bits_stateVec_3_rfile_14      (dbg_bits_stateVec_rfile[3][14]),
    .dbg_bits_stateVec_3_rfile_15      (dbg_bits_stateVec_rfile[3][15]),
    .dbg_bits_stateVec_3_rfile_16      (dbg_bits_stateVec_rfile[3][16]),
    .dbg_bits_stateVec_3_rfile_17      (dbg_bits_stateVec_rfile[3][17]),
    .dbg_bits_stateVec_3_rfile_18      (dbg_bits_stateVec_rfile[3][18]),
    .dbg_bits_stateVec_3_rfile_19      (dbg_bits_stateVec_rfile[3][19]),
    .dbg_bits_stateVec_3_rfile_20      (dbg_bits_stateVec_rfile[3][20]),
    .dbg_bits_stateVec_3_rfile_21      (dbg_bits_stateVec_rfile[3][21]),
    .dbg_bits_stateVec_3_rfile_22      (dbg_bits_stateVec_rfile[3][22]),
    .dbg_bits_stateVec_3_rfile_23      (dbg_bits_stateVec_rfile[3][23]),
    .dbg_bits_stateVec_3_rfile_24      (dbg_bits_stateVec_rfile[3][24]),
    .dbg_bits_stateVec_3_rfile_25      (dbg_bits_stateVec_rfile[3][25]),
    .dbg_bits_stateVec_3_rfile_26      (dbg_bits_stateVec_rfile[3][26]),
    .dbg_bits_stateVec_3_rfile_27      (dbg_bits_stateVec_rfile[3][27]),
    .dbg_bits_stateVec_3_rfile_28      (dbg_bits_stateVec_rfile[3][28]),
    .dbg_bits_stateVec_3_rfile_29      (dbg_bits_stateVec_rfile[3][29]),
    .dbg_bits_stateVec_3_rfile_30      (dbg_bits_stateVec_rfile[3][30]),
    .dbg_bits_stateVec_3_rfile_31      (dbg_bits_stateVec_rfile[3][31]),
    .dbg_bits_stateVec_3_regs_PC       (dbg_bits_stateVec_regs_PC[3]),
    .dbg_bits_stateVec_3_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[3]),
    .dbg_bits_stateVec_4_rfile_0       (dbg_bits_stateVec_rfile[4][0 ]),
    .dbg_bits_stateVec_4_rfile_1       (dbg_bits_stateVec_rfile[4][1 ]),
    .dbg_bits_stateVec_4_rfile_2       (dbg_bits_stateVec_rfile[4][2 ]),
    .dbg_bits_stateVec_4_rfile_3       (dbg_bits_stateVec_rfile[4][3 ]),
    .dbg_bits_stateVec_4_rfile_4       (dbg_bits_stateVec_rfile[4][4 ]),
    .dbg_bits_stateVec_4_rfile_5       (dbg_bits_stateVec_rfile[4][5 ]),
    .dbg_bits_stateVec_4_rfile_6       (dbg_bits_stateVec_rfile[4][6 ]),
    .dbg_bits_stateVec_4_rfile_7       (dbg_bits_stateVec_rfile[4][7 ]),
    .dbg_bits_stateVec_4_rfile_8       (dbg_bits_stateVec_rfile[4][8 ]),
    .dbg_bits_stateVec_4_rfile_9       (dbg_bits_stateVec_rfile[4][9 ]),
    .dbg_bits_stateVec_4_rfile_10      (dbg_bits_stateVec_rfile[4][10]),
    .dbg_bits_stateVec_4_rfile_11      (dbg_bits_stateVec_rfile[4][11]),
    .dbg_bits_stateVec_4_rfile_12      (dbg_bits_stateVec_rfile[4][12]),
    .dbg_bits_stateVec_4_rfile_13      (dbg_bits_stateVec_rfile[4][13]),
    .dbg_bits_stateVec_4_rfile_14      (dbg_bits_stateVec_rfile[4][14]),
    .dbg_bits_stateVec_4_rfile_15      (dbg_bits_stateVec_rfile[4][15]),
    .dbg_bits_stateVec_4_rfile_16      (dbg_bits_stateVec_rfile[4][16]),
    .dbg_bits_stateVec_4_rfile_17      (dbg_bits_stateVec_rfile[4][17]),
    .dbg_bits_stateVec_4_rfile_18      (dbg_bits_stateVec_rfile[4][18]),
    .dbg_bits_stateVec_4_rfile_19      (dbg_bits_stateVec_rfile[4][19]),
    .dbg_bits_stateVec_4_rfile_20      (dbg_bits_stateVec_rfile[4][20]),
    .dbg_bits_stateVec_4_rfile_21      (dbg_bits_stateVec_rfile[4][21]),
    .dbg_bits_stateVec_4_rfile_22      (dbg_bits_stateVec_rfile[4][22]),
    .dbg_bits_stateVec_4_rfile_23      (dbg_bits_stateVec_rfile[4][23]),
    .dbg_bits_stateVec_4_rfile_24      (dbg_bits_stateVec_rfile[4][24]),
    .dbg_bits_stateVec_4_rfile_25      (dbg_bits_stateVec_rfile[4][25]),
    .dbg_bits_stateVec_4_rfile_26      (dbg_bits_stateVec_rfile[4][26]),
    .dbg_bits_stateVec_4_rfile_27      (dbg_bits_stateVec_rfile[4][27]),
    .dbg_bits_stateVec_4_rfile_28      (dbg_bits_stateVec_rfile[4][28]),
    .dbg_bits_stateVec_4_rfile_29      (dbg_bits_stateVec_rfile[4][29]),
    .dbg_bits_stateVec_4_rfile_30      (dbg_bits_stateVec_rfile[4][30]),
    .dbg_bits_stateVec_4_rfile_31      (dbg_bits_stateVec_rfile[4][31]),
    .dbg_bits_stateVec_4_regs_PC       (dbg_bits_stateVec_regs_PC[4]),
    .dbg_bits_stateVec_4_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[4]),
    .dbg_bits_stateVec_5_rfile_0       (dbg_bits_stateVec_rfile[5][0 ]),
    .dbg_bits_stateVec_5_rfile_1       (dbg_bits_stateVec_rfile[5][1 ]),
    .dbg_bits_stateVec_5_rfile_2       (dbg_bits_stateVec_rfile[5][2 ]),
    .dbg_bits_stateVec_5_rfile_3       (dbg_bits_stateVec_rfile[5][3 ]),
    .dbg_bits_stateVec_5_rfile_4       (dbg_bits_stateVec_rfile[5][4 ]),
    .dbg_bits_stateVec_5_rfile_5       (dbg_bits_stateVec_rfile[5][5 ]),
    .dbg_bits_stateVec_5_rfile_6       (dbg_bits_stateVec_rfile[5][6 ]),
    .dbg_bits_stateVec_5_rfile_7       (dbg_bits_stateVec_rfile[5][7 ]),
    .dbg_bits_stateVec_5_rfile_8       (dbg_bits_stateVec_rfile[5][8 ]),
    .dbg_bits_stateVec_5_rfile_9       (dbg_bits_stateVec_rfile[5][9 ]),
    .dbg_bits_stateVec_5_rfile_10      (dbg_bits_stateVec_rfile[5][10]),
    .dbg_bits_stateVec_5_rfile_11      (dbg_bits_stateVec_rfile[5][11]),
    .dbg_bits_stateVec_5_rfile_12      (dbg_bits_stateVec_rfile[5][12]),
    .dbg_bits_stateVec_5_rfile_13      (dbg_bits_stateVec_rfile[5][13]),
    .dbg_bits_stateVec_5_rfile_14      (dbg_bits_stateVec_rfile[5][14]),
    .dbg_bits_stateVec_5_rfile_15      (dbg_bits_stateVec_rfile[5][15]),
    .dbg_bits_stateVec_5_rfile_16      (dbg_bits_stateVec_rfile[5][16]),
    .dbg_bits_stateVec_5_rfile_17      (dbg_bits_stateVec_rfile[5][17]),
    .dbg_bits_stateVec_5_rfile_18      (dbg_bits_stateVec_rfile[5][18]),
    .dbg_bits_stateVec_5_rfile_19      (dbg_bits_stateVec_rfile[5][19]),
    .dbg_bits_stateVec_5_rfile_20      (dbg_bits_stateVec_rfile[5][20]),
    .dbg_bits_stateVec_5_rfile_21      (dbg_bits_stateVec_rfile[5][21]),
    .dbg_bits_stateVec_5_rfile_22      (dbg_bits_stateVec_rfile[5][22]),
    .dbg_bits_stateVec_5_rfile_23      (dbg_bits_stateVec_rfile[5][23]),
    .dbg_bits_stateVec_5_rfile_24      (dbg_bits_stateVec_rfile[5][24]),
    .dbg_bits_stateVec_5_rfile_25      (dbg_bits_stateVec_rfile[5][25]),
    .dbg_bits_stateVec_5_rfile_26      (dbg_bits_stateVec_rfile[5][26]),
    .dbg_bits_stateVec_5_rfile_27      (dbg_bits_stateVec_rfile[5][27]),
    .dbg_bits_stateVec_5_rfile_28      (dbg_bits_stateVec_rfile[5][28]),
    .dbg_bits_stateVec_5_rfile_29      (dbg_bits_stateVec_rfile[5][29]),
    .dbg_bits_stateVec_5_rfile_30      (dbg_bits_stateVec_rfile[5][30]),
    .dbg_bits_stateVec_5_rfile_31      (dbg_bits_stateVec_rfile[5][31]),
    .dbg_bits_stateVec_5_regs_PC       (dbg_bits_stateVec_regs_PC[5]),
    .dbg_bits_stateVec_5_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[5]),
    .dbg_bits_stateVec_6_rfile_0       (dbg_bits_stateVec_rfile[6][0 ]),
    .dbg_bits_stateVec_6_rfile_1       (dbg_bits_stateVec_rfile[6][1 ]),
    .dbg_bits_stateVec_6_rfile_2       (dbg_bits_stateVec_rfile[6][2 ]),
    .dbg_bits_stateVec_6_rfile_3       (dbg_bits_stateVec_rfile[6][3 ]),
    .dbg_bits_stateVec_6_rfile_4       (dbg_bits_stateVec_rfile[6][4 ]),
    .dbg_bits_stateVec_6_rfile_5       (dbg_bits_stateVec_rfile[6][5 ]),
    .dbg_bits_stateVec_6_rfile_6       (dbg_bits_stateVec_rfile[6][6 ]),
    .dbg_bits_stateVec_6_rfile_7       (dbg_bits_stateVec_rfile[6][7 ]),
    .dbg_bits_stateVec_6_rfile_8       (dbg_bits_stateVec_rfile[6][8 ]),
    .dbg_bits_stateVec_6_rfile_9       (dbg_bits_stateVec_rfile[6][9 ]),
    .dbg_bits_stateVec_6_rfile_10      (dbg_bits_stateVec_rfile[6][10]),
    .dbg_bits_stateVec_6_rfile_11      (dbg_bits_stateVec_rfile[6][11]),
    .dbg_bits_stateVec_6_rfile_12      (dbg_bits_stateVec_rfile[6][12]),
    .dbg_bits_stateVec_6_rfile_13      (dbg_bits_stateVec_rfile[6][13]),
    .dbg_bits_stateVec_6_rfile_14      (dbg_bits_stateVec_rfile[6][14]),
    .dbg_bits_stateVec_6_rfile_15      (dbg_bits_stateVec_rfile[6][15]),
    .dbg_bits_stateVec_6_rfile_16      (dbg_bits_stateVec_rfile[6][16]),
    .dbg_bits_stateVec_6_rfile_17      (dbg_bits_stateVec_rfile[6][17]),
    .dbg_bits_stateVec_6_rfile_18      (dbg_bits_stateVec_rfile[6][18]),
    .dbg_bits_stateVec_6_rfile_19      (dbg_bits_stateVec_rfile[6][19]),
    .dbg_bits_stateVec_6_rfile_20      (dbg_bits_stateVec_rfile[6][20]),
    .dbg_bits_stateVec_6_rfile_21      (dbg_bits_stateVec_rfile[6][21]),
    .dbg_bits_stateVec_6_rfile_22      (dbg_bits_stateVec_rfile[6][22]),
    .dbg_bits_stateVec_6_rfile_23      (dbg_bits_stateVec_rfile[6][23]),
    .dbg_bits_stateVec_6_rfile_24      (dbg_bits_stateVec_rfile[6][24]),
    .dbg_bits_stateVec_6_rfile_25      (dbg_bits_stateVec_rfile[6][25]),
    .dbg_bits_stateVec_6_rfile_26      (dbg_bits_stateVec_rfile[6][26]),
    .dbg_bits_stateVec_6_rfile_27      (dbg_bits_stateVec_rfile[6][27]),
    .dbg_bits_stateVec_6_rfile_28      (dbg_bits_stateVec_rfile[6][28]),
    .dbg_bits_stateVec_6_rfile_29      (dbg_bits_stateVec_rfile[6][29]),
    .dbg_bits_stateVec_6_rfile_30      (dbg_bits_stateVec_rfile[6][30]),
    .dbg_bits_stateVec_6_rfile_31      (dbg_bits_stateVec_rfile[6][31]),
    .dbg_bits_stateVec_6_regs_PC       (dbg_bits_stateVec_regs_PC[6]),
    .dbg_bits_stateVec_6_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[6]),
    .dbg_bits_stateVec_7_rfile_0       (dbg_bits_stateVec_rfile[7][0 ]),
    .dbg_bits_stateVec_7_rfile_1       (dbg_bits_stateVec_rfile[7][1 ]),
    .dbg_bits_stateVec_7_rfile_2       (dbg_bits_stateVec_rfile[7][2 ]),
    .dbg_bits_stateVec_7_rfile_3       (dbg_bits_stateVec_rfile[7][3 ]),
    .dbg_bits_stateVec_7_rfile_4       (dbg_bits_stateVec_rfile[7][4 ]),
    .dbg_bits_stateVec_7_rfile_5       (dbg_bits_stateVec_rfile[7][5 ]),
    .dbg_bits_stateVec_7_rfile_6       (dbg_bits_stateVec_rfile[7][6 ]),
    .dbg_bits_stateVec_7_rfile_7       (dbg_bits_stateVec_rfile[7][7 ]),
    .dbg_bits_stateVec_7_rfile_8       (dbg_bits_stateVec_rfile[7][8 ]),
    .dbg_bits_stateVec_7_rfile_9       (dbg_bits_stateVec_rfile[7][9 ]),
    .dbg_bits_stateVec_7_rfile_10      (dbg_bits_stateVec_rfile[7][10]),
    .dbg_bits_stateVec_7_rfile_11      (dbg_bits_stateVec_rfile[7][11]),
    .dbg_bits_stateVec_7_rfile_12      (dbg_bits_stateVec_rfile[7][12]),
    .dbg_bits_stateVec_7_rfile_13      (dbg_bits_stateVec_rfile[7][13]),
    .dbg_bits_stateVec_7_rfile_14      (dbg_bits_stateVec_rfile[7][14]),
    .dbg_bits_stateVec_7_rfile_15      (dbg_bits_stateVec_rfile[7][15]),
    .dbg_bits_stateVec_7_rfile_16      (dbg_bits_stateVec_rfile[7][16]),
    .dbg_bits_stateVec_7_rfile_17      (dbg_bits_stateVec_rfile[7][17]),
    .dbg_bits_stateVec_7_rfile_18      (dbg_bits_stateVec_rfile[7][18]),
    .dbg_bits_stateVec_7_rfile_19      (dbg_bits_stateVec_rfile[7][19]),
    .dbg_bits_stateVec_7_rfile_20      (dbg_bits_stateVec_rfile[7][20]),
    .dbg_bits_stateVec_7_rfile_21      (dbg_bits_stateVec_rfile[7][21]),
    .dbg_bits_stateVec_7_rfile_22      (dbg_bits_stateVec_rfile[7][22]),
    .dbg_bits_stateVec_7_rfile_23      (dbg_bits_stateVec_rfile[7][23]),
    .dbg_bits_stateVec_7_rfile_24      (dbg_bits_stateVec_rfile[7][24]),
    .dbg_bits_stateVec_7_rfile_25      (dbg_bits_stateVec_rfile[7][25]),
    .dbg_bits_stateVec_7_rfile_26      (dbg_bits_stateVec_rfile[7][26]),
    .dbg_bits_stateVec_7_rfile_27      (dbg_bits_stateVec_rfile[7][27]),
    .dbg_bits_stateVec_7_rfile_28      (dbg_bits_stateVec_rfile[7][28]),
    .dbg_bits_stateVec_7_rfile_29      (dbg_bits_stateVec_rfile[7][29]),
    .dbg_bits_stateVec_7_rfile_30      (dbg_bits_stateVec_rfile[7][30]),
    .dbg_bits_stateVec_7_rfile_31      (dbg_bits_stateVec_rfile[7][31]),
    .dbg_bits_stateVec_7_regs_PC       (dbg_bits_stateVec_regs_PC[7]),
    .dbg_bits_stateVec_7_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[7]),
    .dbg_bits_stateVec_8_rfile_0       (dbg_bits_stateVec_rfile[8][0 ]),
    .dbg_bits_stateVec_8_rfile_1       (dbg_bits_stateVec_rfile[8][1 ]),
    .dbg_bits_stateVec_8_rfile_2       (dbg_bits_stateVec_rfile[8][2 ]),
    .dbg_bits_stateVec_8_rfile_3       (dbg_bits_stateVec_rfile[8][3 ]),
    .dbg_bits_stateVec_8_rfile_4       (dbg_bits_stateVec_rfile[8][4 ]),
    .dbg_bits_stateVec_8_rfile_5       (dbg_bits_stateVec_rfile[8][5 ]),
    .dbg_bits_stateVec_8_rfile_6       (dbg_bits_stateVec_rfile[8][6 ]),
    .dbg_bits_stateVec_8_rfile_7       (dbg_bits_stateVec_rfile[8][7 ]),
    .dbg_bits_stateVec_8_rfile_8       (dbg_bits_stateVec_rfile[8][8 ]),
    .dbg_bits_stateVec_8_rfile_9       (dbg_bits_stateVec_rfile[8][9 ]),
    .dbg_bits_stateVec_8_rfile_10      (dbg_bits_stateVec_rfile[8][10]),
    .dbg_bits_stateVec_8_rfile_11      (dbg_bits_stateVec_rfile[8][11]),
    .dbg_bits_stateVec_8_rfile_12      (dbg_bits_stateVec_rfile[8][12]),
    .dbg_bits_stateVec_8_rfile_13      (dbg_bits_stateVec_rfile[8][13]),
    .dbg_bits_stateVec_8_rfile_14      (dbg_bits_stateVec_rfile[8][14]),
    .dbg_bits_stateVec_8_rfile_15      (dbg_bits_stateVec_rfile[8][15]),
    .dbg_bits_stateVec_8_rfile_16      (dbg_bits_stateVec_rfile[8][16]),
    .dbg_bits_stateVec_8_rfile_17      (dbg_bits_stateVec_rfile[8][17]),
    .dbg_bits_stateVec_8_rfile_18      (dbg_bits_stateVec_rfile[8][18]),
    .dbg_bits_stateVec_8_rfile_19      (dbg_bits_stateVec_rfile[8][19]),
    .dbg_bits_stateVec_8_rfile_20      (dbg_bits_stateVec_rfile[8][20]),
    .dbg_bits_stateVec_8_rfile_21      (dbg_bits_stateVec_rfile[8][21]),
    .dbg_bits_stateVec_8_rfile_22      (dbg_bits_stateVec_rfile[8][22]),
    .dbg_bits_stateVec_8_rfile_23      (dbg_bits_stateVec_rfile[8][23]),
    .dbg_bits_stateVec_8_rfile_24      (dbg_bits_stateVec_rfile[8][24]),
    .dbg_bits_stateVec_8_rfile_25      (dbg_bits_stateVec_rfile[8][25]),
    .dbg_bits_stateVec_8_rfile_26      (dbg_bits_stateVec_rfile[8][26]),
    .dbg_bits_stateVec_8_rfile_27      (dbg_bits_stateVec_rfile[8][27]),
    .dbg_bits_stateVec_8_rfile_28      (dbg_bits_stateVec_rfile[8][28]),
    .dbg_bits_stateVec_8_rfile_29      (dbg_bits_stateVec_rfile[8][29]),
    .dbg_bits_stateVec_8_rfile_30      (dbg_bits_stateVec_rfile[8][30]),
    .dbg_bits_stateVec_8_rfile_31      (dbg_bits_stateVec_rfile[8][31]),
    .dbg_bits_stateVec_8_regs_PC       (dbg_bits_stateVec_regs_PC[8]),
    .dbg_bits_stateVec_8_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[8]),
    .dbg_bits_stateVec_9_rfile_0       (dbg_bits_stateVec_rfile[9][0 ]),
    .dbg_bits_stateVec_9_rfile_1       (dbg_bits_stateVec_rfile[9][1 ]),
    .dbg_bits_stateVec_9_rfile_2       (dbg_bits_stateVec_rfile[9][2 ]),
    .dbg_bits_stateVec_9_rfile_3       (dbg_bits_stateVec_rfile[9][3 ]),
    .dbg_bits_stateVec_9_rfile_4       (dbg_bits_stateVec_rfile[9][4 ]),
    .dbg_bits_stateVec_9_rfile_5       (dbg_bits_stateVec_rfile[9][5 ]),
    .dbg_bits_stateVec_9_rfile_6       (dbg_bits_stateVec_rfile[9][6 ]),
    .dbg_bits_stateVec_9_rfile_7       (dbg_bits_stateVec_rfile[9][7 ]),
    .dbg_bits_stateVec_9_rfile_8       (dbg_bits_stateVec_rfile[9][8 ]),
    .dbg_bits_stateVec_9_rfile_9       (dbg_bits_stateVec_rfile[9][9 ]),
    .dbg_bits_stateVec_9_rfile_10      (dbg_bits_stateVec_rfile[9][10]),
    .dbg_bits_stateVec_9_rfile_11      (dbg_bits_stateVec_rfile[9][11]),
    .dbg_bits_stateVec_9_rfile_12      (dbg_bits_stateVec_rfile[9][12]),
    .dbg_bits_stateVec_9_rfile_13      (dbg_bits_stateVec_rfile[9][13]),
    .dbg_bits_stateVec_9_rfile_14      (dbg_bits_stateVec_rfile[9][14]),
    .dbg_bits_stateVec_9_rfile_15      (dbg_bits_stateVec_rfile[9][15]),
    .dbg_bits_stateVec_9_rfile_16      (dbg_bits_stateVec_rfile[9][16]),
    .dbg_bits_stateVec_9_rfile_17      (dbg_bits_stateVec_rfile[9][17]),
    .dbg_bits_stateVec_9_rfile_18      (dbg_bits_stateVec_rfile[9][18]),
    .dbg_bits_stateVec_9_rfile_19      (dbg_bits_stateVec_rfile[9][19]),
    .dbg_bits_stateVec_9_rfile_20      (dbg_bits_stateVec_rfile[9][20]),
    .dbg_bits_stateVec_9_rfile_21      (dbg_bits_stateVec_rfile[9][21]),
    .dbg_bits_stateVec_9_rfile_22      (dbg_bits_stateVec_rfile[9][22]),
    .dbg_bits_stateVec_9_rfile_23      (dbg_bits_stateVec_rfile[9][23]),
    .dbg_bits_stateVec_9_rfile_24      (dbg_bits_stateVec_rfile[9][24]),
    .dbg_bits_stateVec_9_rfile_25      (dbg_bits_stateVec_rfile[9][25]),
    .dbg_bits_stateVec_9_rfile_26      (dbg_bits_stateVec_rfile[9][26]),
    .dbg_bits_stateVec_9_rfile_27      (dbg_bits_stateVec_rfile[9][27]),
    .dbg_bits_stateVec_9_rfile_28      (dbg_bits_stateVec_rfile[9][28]),
    .dbg_bits_stateVec_9_rfile_29      (dbg_bits_stateVec_rfile[9][29]),
    .dbg_bits_stateVec_9_rfile_30      (dbg_bits_stateVec_rfile[9][30]),
    .dbg_bits_stateVec_9_rfile_31      (dbg_bits_stateVec_rfile[9][31]),
    .dbg_bits_stateVec_9_regs_PC       (dbg_bits_stateVec_regs_PC[9]),
    .dbg_bits_stateVec_9_regs_NZCV     (dbg_bits_stateVec_regs_NZCV[9]),
    .dbg_bits_stateVec_10_rfile_0      (dbg_bits_stateVec_rfile[10][0 ]),
    .dbg_bits_stateVec_10_rfile_1      (dbg_bits_stateVec_rfile[10][1 ]),
    .dbg_bits_stateVec_10_rfile_2      (dbg_bits_stateVec_rfile[10][2 ]),
    .dbg_bits_stateVec_10_rfile_3      (dbg_bits_stateVec_rfile[10][3 ]),
    .dbg_bits_stateVec_10_rfile_4      (dbg_bits_stateVec_rfile[10][4 ]),
    .dbg_bits_stateVec_10_rfile_5      (dbg_bits_stateVec_rfile[10][5 ]),
    .dbg_bits_stateVec_10_rfile_6      (dbg_bits_stateVec_rfile[10][6 ]),
    .dbg_bits_stateVec_10_rfile_7      (dbg_bits_stateVec_rfile[10][7 ]),
    .dbg_bits_stateVec_10_rfile_8      (dbg_bits_stateVec_rfile[10][8 ]),
    .dbg_bits_stateVec_10_rfile_9      (dbg_bits_stateVec_rfile[10][9 ]),
    .dbg_bits_stateVec_10_rfile_10     (dbg_bits_stateVec_rfile[10][10]),
    .dbg_bits_stateVec_10_rfile_11     (dbg_bits_stateVec_rfile[10][11]),
    .dbg_bits_stateVec_10_rfile_12     (dbg_bits_stateVec_rfile[10][12]),
    .dbg_bits_stateVec_10_rfile_13     (dbg_bits_stateVec_rfile[10][13]),
    .dbg_bits_stateVec_10_rfile_14     (dbg_bits_stateVec_rfile[10][14]),
    .dbg_bits_stateVec_10_rfile_15     (dbg_bits_stateVec_rfile[10][15]),
    .dbg_bits_stateVec_10_rfile_16     (dbg_bits_stateVec_rfile[10][16]),
    .dbg_bits_stateVec_10_rfile_17     (dbg_bits_stateVec_rfile[10][17]),
    .dbg_bits_stateVec_10_rfile_18     (dbg_bits_stateVec_rfile[10][18]),
    .dbg_bits_stateVec_10_rfile_19     (dbg_bits_stateVec_rfile[10][19]),
    .dbg_bits_stateVec_10_rfile_20     (dbg_bits_stateVec_rfile[10][20]),
    .dbg_bits_stateVec_10_rfile_21     (dbg_bits_stateVec_rfile[10][21]),
    .dbg_bits_stateVec_10_rfile_22     (dbg_bits_stateVec_rfile[10][22]),
    .dbg_bits_stateVec_10_rfile_23     (dbg_bits_stateVec_rfile[10][23]),
    .dbg_bits_stateVec_10_rfile_24     (dbg_bits_stateVec_rfile[10][24]),
    .dbg_bits_stateVec_10_rfile_25     (dbg_bits_stateVec_rfile[10][25]),
    .dbg_bits_stateVec_10_rfile_26     (dbg_bits_stateVec_rfile[10][26]),
    .dbg_bits_stateVec_10_rfile_27     (dbg_bits_stateVec_rfile[10][27]),
    .dbg_bits_stateVec_10_rfile_28     (dbg_bits_stateVec_rfile[10][28]),
    .dbg_bits_stateVec_10_rfile_29     (dbg_bits_stateVec_rfile[10][29]),
    .dbg_bits_stateVec_10_rfile_30     (dbg_bits_stateVec_rfile[10][30]),
    .dbg_bits_stateVec_10_rfile_31     (dbg_bits_stateVec_rfile[10][31]),
    .dbg_bits_stateVec_10_regs_PC      (dbg_bits_stateVec_regs_PC  [10]),
    .dbg_bits_stateVec_10_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[10]),
    .dbg_bits_stateVec_11_rfile_0      (dbg_bits_stateVec_rfile[11][0 ]),
    .dbg_bits_stateVec_11_rfile_1      (dbg_bits_stateVec_rfile[11][1 ]),
    .dbg_bits_stateVec_11_rfile_2      (dbg_bits_stateVec_rfile[11][2 ]),
    .dbg_bits_stateVec_11_rfile_3      (dbg_bits_stateVec_rfile[11][3 ]),
    .dbg_bits_stateVec_11_rfile_4      (dbg_bits_stateVec_rfile[11][4 ]),
    .dbg_bits_stateVec_11_rfile_5      (dbg_bits_stateVec_rfile[11][5 ]),
    .dbg_bits_stateVec_11_rfile_6      (dbg_bits_stateVec_rfile[11][6 ]),
    .dbg_bits_stateVec_11_rfile_7      (dbg_bits_stateVec_rfile[11][7 ]),
    .dbg_bits_stateVec_11_rfile_8      (dbg_bits_stateVec_rfile[11][8 ]),
    .dbg_bits_stateVec_11_rfile_9      (dbg_bits_stateVec_rfile[11][9 ]),
    .dbg_bits_stateVec_11_rfile_10     (dbg_bits_stateVec_rfile[11][10]),
    .dbg_bits_stateVec_11_rfile_11     (dbg_bits_stateVec_rfile[11][11]),
    .dbg_bits_stateVec_11_rfile_12     (dbg_bits_stateVec_rfile[11][12]),
    .dbg_bits_stateVec_11_rfile_13     (dbg_bits_stateVec_rfile[11][13]),
    .dbg_bits_stateVec_11_rfile_14     (dbg_bits_stateVec_rfile[11][14]),
    .dbg_bits_stateVec_11_rfile_15     (dbg_bits_stateVec_rfile[11][15]),
    .dbg_bits_stateVec_11_rfile_16     (dbg_bits_stateVec_rfile[11][16]),
    .dbg_bits_stateVec_11_rfile_17     (dbg_bits_stateVec_rfile[11][17]),
    .dbg_bits_stateVec_11_rfile_18     (dbg_bits_stateVec_rfile[11][18]),
    .dbg_bits_stateVec_11_rfile_19     (dbg_bits_stateVec_rfile[11][19]),
    .dbg_bits_stateVec_11_rfile_20     (dbg_bits_stateVec_rfile[11][20]),
    .dbg_bits_stateVec_11_rfile_21     (dbg_bits_stateVec_rfile[11][21]),
    .dbg_bits_stateVec_11_rfile_22     (dbg_bits_stateVec_rfile[11][22]),
    .dbg_bits_stateVec_11_rfile_23     (dbg_bits_stateVec_rfile[11][23]),
    .dbg_bits_stateVec_11_rfile_24     (dbg_bits_stateVec_rfile[11][24]),
    .dbg_bits_stateVec_11_rfile_25     (dbg_bits_stateVec_rfile[11][25]),
    .dbg_bits_stateVec_11_rfile_26     (dbg_bits_stateVec_rfile[11][26]),
    .dbg_bits_stateVec_11_rfile_27     (dbg_bits_stateVec_rfile[11][27]),
    .dbg_bits_stateVec_11_rfile_28     (dbg_bits_stateVec_rfile[11][28]),
    .dbg_bits_stateVec_11_rfile_29     (dbg_bits_stateVec_rfile[11][29]),
    .dbg_bits_stateVec_11_rfile_30     (dbg_bits_stateVec_rfile[11][30]),
    .dbg_bits_stateVec_11_rfile_31     (dbg_bits_stateVec_rfile[11][31]),
    .dbg_bits_stateVec_11_regs_PC      (dbg_bits_stateVec_regs_PC  [11]),
    .dbg_bits_stateVec_11_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[11]),
    .dbg_bits_stateVec_12_rfile_0      (dbg_bits_stateVec_rfile[12][0 ]),
    .dbg_bits_stateVec_12_rfile_1      (dbg_bits_stateVec_rfile[12][1 ]),
    .dbg_bits_stateVec_12_rfile_2      (dbg_bits_stateVec_rfile[12][2 ]),
    .dbg_bits_stateVec_12_rfile_3      (dbg_bits_stateVec_rfile[12][3 ]),
    .dbg_bits_stateVec_12_rfile_4      (dbg_bits_stateVec_rfile[12][4 ]),
    .dbg_bits_stateVec_12_rfile_5      (dbg_bits_stateVec_rfile[12][5 ]),
    .dbg_bits_stateVec_12_rfile_6      (dbg_bits_stateVec_rfile[12][6 ]),
    .dbg_bits_stateVec_12_rfile_7      (dbg_bits_stateVec_rfile[12][7 ]),
    .dbg_bits_stateVec_12_rfile_8      (dbg_bits_stateVec_rfile[12][8 ]),
    .dbg_bits_stateVec_12_rfile_9      (dbg_bits_stateVec_rfile[12][9 ]),
    .dbg_bits_stateVec_12_rfile_10     (dbg_bits_stateVec_rfile[12][10]),
    .dbg_bits_stateVec_12_rfile_11     (dbg_bits_stateVec_rfile[12][11]),
    .dbg_bits_stateVec_12_rfile_12     (dbg_bits_stateVec_rfile[12][12]),
    .dbg_bits_stateVec_12_rfile_13     (dbg_bits_stateVec_rfile[12][13]),
    .dbg_bits_stateVec_12_rfile_14     (dbg_bits_stateVec_rfile[12][14]),
    .dbg_bits_stateVec_12_rfile_15     (dbg_bits_stateVec_rfile[12][15]),
    .dbg_bits_stateVec_12_rfile_16     (dbg_bits_stateVec_rfile[12][16]),
    .dbg_bits_stateVec_12_rfile_17     (dbg_bits_stateVec_rfile[12][17]),
    .dbg_bits_stateVec_12_rfile_18     (dbg_bits_stateVec_rfile[12][18]),
    .dbg_bits_stateVec_12_rfile_19     (dbg_bits_stateVec_rfile[12][19]),
    .dbg_bits_stateVec_12_rfile_20     (dbg_bits_stateVec_rfile[12][20]),
    .dbg_bits_stateVec_12_rfile_21     (dbg_bits_stateVec_rfile[12][21]),
    .dbg_bits_stateVec_12_rfile_22     (dbg_bits_stateVec_rfile[12][22]),
    .dbg_bits_stateVec_12_rfile_23     (dbg_bits_stateVec_rfile[12][23]),
    .dbg_bits_stateVec_12_rfile_24     (dbg_bits_stateVec_rfile[12][24]),
    .dbg_bits_stateVec_12_rfile_25     (dbg_bits_stateVec_rfile[12][25]),
    .dbg_bits_stateVec_12_rfile_26     (dbg_bits_stateVec_rfile[12][26]),
    .dbg_bits_stateVec_12_rfile_27     (dbg_bits_stateVec_rfile[12][27]),
    .dbg_bits_stateVec_12_rfile_28     (dbg_bits_stateVec_rfile[12][28]),
    .dbg_bits_stateVec_12_rfile_29     (dbg_bits_stateVec_rfile[12][29]),
    .dbg_bits_stateVec_12_rfile_30     (dbg_bits_stateVec_rfile[12][30]),
    .dbg_bits_stateVec_12_rfile_31     (dbg_bits_stateVec_rfile[12][31]),
    .dbg_bits_stateVec_12_regs_PC      (dbg_bits_stateVec_regs_PC  [12]),
    .dbg_bits_stateVec_12_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[12]),
    .dbg_bits_stateVec_13_rfile_0      (dbg_bits_stateVec_rfile[13][0 ]),
    .dbg_bits_stateVec_13_rfile_1      (dbg_bits_stateVec_rfile[13][1 ]),
    .dbg_bits_stateVec_13_rfile_2      (dbg_bits_stateVec_rfile[13][2 ]),
    .dbg_bits_stateVec_13_rfile_3      (dbg_bits_stateVec_rfile[13][3 ]),
    .dbg_bits_stateVec_13_rfile_4      (dbg_bits_stateVec_rfile[13][4 ]),
    .dbg_bits_stateVec_13_rfile_5      (dbg_bits_stateVec_rfile[13][5 ]),
    .dbg_bits_stateVec_13_rfile_6      (dbg_bits_stateVec_rfile[13][6 ]),
    .dbg_bits_stateVec_13_rfile_7      (dbg_bits_stateVec_rfile[13][7 ]),
    .dbg_bits_stateVec_13_rfile_8      (dbg_bits_stateVec_rfile[13][8 ]),
    .dbg_bits_stateVec_13_rfile_9      (dbg_bits_stateVec_rfile[13][9 ]),
    .dbg_bits_stateVec_13_rfile_10     (dbg_bits_stateVec_rfile[13][10]),
    .dbg_bits_stateVec_13_rfile_11     (dbg_bits_stateVec_rfile[13][11]),
    .dbg_bits_stateVec_13_rfile_12     (dbg_bits_stateVec_rfile[13][12]),
    .dbg_bits_stateVec_13_rfile_13     (dbg_bits_stateVec_rfile[13][13]),
    .dbg_bits_stateVec_13_rfile_14     (dbg_bits_stateVec_rfile[13][14]),
    .dbg_bits_stateVec_13_rfile_15     (dbg_bits_stateVec_rfile[13][15]),
    .dbg_bits_stateVec_13_rfile_16     (dbg_bits_stateVec_rfile[13][16]),
    .dbg_bits_stateVec_13_rfile_17     (dbg_bits_stateVec_rfile[13][17]),
    .dbg_bits_stateVec_13_rfile_18     (dbg_bits_stateVec_rfile[13][18]),
    .dbg_bits_stateVec_13_rfile_19     (dbg_bits_stateVec_rfile[13][19]),
    .dbg_bits_stateVec_13_rfile_20     (dbg_bits_stateVec_rfile[13][20]),
    .dbg_bits_stateVec_13_rfile_21     (dbg_bits_stateVec_rfile[13][21]),
    .dbg_bits_stateVec_13_rfile_22     (dbg_bits_stateVec_rfile[13][22]),
    .dbg_bits_stateVec_13_rfile_23     (dbg_bits_stateVec_rfile[13][23]),
    .dbg_bits_stateVec_13_rfile_24     (dbg_bits_stateVec_rfile[13][24]),
    .dbg_bits_stateVec_13_rfile_25     (dbg_bits_stateVec_rfile[13][25]),
    .dbg_bits_stateVec_13_rfile_26     (dbg_bits_stateVec_rfile[13][26]),
    .dbg_bits_stateVec_13_rfile_27     (dbg_bits_stateVec_rfile[13][27]),
    .dbg_bits_stateVec_13_rfile_28     (dbg_bits_stateVec_rfile[13][28]),
    .dbg_bits_stateVec_13_rfile_29     (dbg_bits_stateVec_rfile[13][29]),
    .dbg_bits_stateVec_13_rfile_30     (dbg_bits_stateVec_rfile[13][30]),
    .dbg_bits_stateVec_13_rfile_31     (dbg_bits_stateVec_rfile[13][31]),
    .dbg_bits_stateVec_13_regs_PC      (dbg_bits_stateVec_regs_PC  [13]),
    .dbg_bits_stateVec_13_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[13]),
    .dbg_bits_stateVec_14_rfile_0      (dbg_bits_stateVec_rfile[14][0 ]),
    .dbg_bits_stateVec_14_rfile_1      (dbg_bits_stateVec_rfile[14][1 ]),
    .dbg_bits_stateVec_14_rfile_2      (dbg_bits_stateVec_rfile[14][2 ]),
    .dbg_bits_stateVec_14_rfile_3      (dbg_bits_stateVec_rfile[14][3 ]),
    .dbg_bits_stateVec_14_rfile_4      (dbg_bits_stateVec_rfile[14][4 ]),
    .dbg_bits_stateVec_14_rfile_5      (dbg_bits_stateVec_rfile[14][5 ]),
    .dbg_bits_stateVec_14_rfile_6      (dbg_bits_stateVec_rfile[14][6 ]),
    .dbg_bits_stateVec_14_rfile_7      (dbg_bits_stateVec_rfile[14][7 ]),
    .dbg_bits_stateVec_14_rfile_8      (dbg_bits_stateVec_rfile[14][8 ]),
    .dbg_bits_stateVec_14_rfile_9      (dbg_bits_stateVec_rfile[14][9 ]),
    .dbg_bits_stateVec_14_rfile_10     (dbg_bits_stateVec_rfile[14][10]),
    .dbg_bits_stateVec_14_rfile_11     (dbg_bits_stateVec_rfile[14][11]),
    .dbg_bits_stateVec_14_rfile_12     (dbg_bits_stateVec_rfile[14][12]),
    .dbg_bits_stateVec_14_rfile_13     (dbg_bits_stateVec_rfile[14][13]),
    .dbg_bits_stateVec_14_rfile_14     (dbg_bits_stateVec_rfile[14][14]),
    .dbg_bits_stateVec_14_rfile_15     (dbg_bits_stateVec_rfile[14][15]),
    .dbg_bits_stateVec_14_rfile_16     (dbg_bits_stateVec_rfile[14][16]),
    .dbg_bits_stateVec_14_rfile_17     (dbg_bits_stateVec_rfile[14][17]),
    .dbg_bits_stateVec_14_rfile_18     (dbg_bits_stateVec_rfile[14][18]),
    .dbg_bits_stateVec_14_rfile_19     (dbg_bits_stateVec_rfile[14][19]),
    .dbg_bits_stateVec_14_rfile_20     (dbg_bits_stateVec_rfile[14][20]),
    .dbg_bits_stateVec_14_rfile_21     (dbg_bits_stateVec_rfile[14][21]),
    .dbg_bits_stateVec_14_rfile_22     (dbg_bits_stateVec_rfile[14][22]),
    .dbg_bits_stateVec_14_rfile_23     (dbg_bits_stateVec_rfile[14][23]),
    .dbg_bits_stateVec_14_rfile_24     (dbg_bits_stateVec_rfile[14][24]),
    .dbg_bits_stateVec_14_rfile_25     (dbg_bits_stateVec_rfile[14][25]),
    .dbg_bits_stateVec_14_rfile_26     (dbg_bits_stateVec_rfile[14][26]),
    .dbg_bits_stateVec_14_rfile_27     (dbg_bits_stateVec_rfile[14][27]),
    .dbg_bits_stateVec_14_rfile_28     (dbg_bits_stateVec_rfile[14][28]),
    .dbg_bits_stateVec_14_rfile_29     (dbg_bits_stateVec_rfile[14][29]),
    .dbg_bits_stateVec_14_rfile_30     (dbg_bits_stateVec_rfile[14][30]),
    .dbg_bits_stateVec_14_rfile_31     (dbg_bits_stateVec_rfile[14][31]),
    .dbg_bits_stateVec_14_regs_PC      (dbg_bits_stateVec_regs_PC  [14]),
    .dbg_bits_stateVec_14_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[14]),
    .dbg_bits_stateVec_15_rfile_0      (dbg_bits_stateVec_rfile[15][0 ]),
    .dbg_bits_stateVec_15_rfile_1      (dbg_bits_stateVec_rfile[15][1 ]),
    .dbg_bits_stateVec_15_rfile_2      (dbg_bits_stateVec_rfile[15][2 ]),
    .dbg_bits_stateVec_15_rfile_3      (dbg_bits_stateVec_rfile[15][3 ]),
    .dbg_bits_stateVec_15_rfile_4      (dbg_bits_stateVec_rfile[15][4 ]),
    .dbg_bits_stateVec_15_rfile_5      (dbg_bits_stateVec_rfile[15][5 ]),
    .dbg_bits_stateVec_15_rfile_6      (dbg_bits_stateVec_rfile[15][6 ]),
    .dbg_bits_stateVec_15_rfile_7      (dbg_bits_stateVec_rfile[15][7 ]),
    .dbg_bits_stateVec_15_rfile_8      (dbg_bits_stateVec_rfile[15][8 ]),
    .dbg_bits_stateVec_15_rfile_9      (dbg_bits_stateVec_rfile[15][9 ]),
    .dbg_bits_stateVec_15_rfile_10     (dbg_bits_stateVec_rfile[15][10]),
    .dbg_bits_stateVec_15_rfile_11     (dbg_bits_stateVec_rfile[15][11]),
    .dbg_bits_stateVec_15_rfile_12     (dbg_bits_stateVec_rfile[15][12]),
    .dbg_bits_stateVec_15_rfile_13     (dbg_bits_stateVec_rfile[15][13]),
    .dbg_bits_stateVec_15_rfile_14     (dbg_bits_stateVec_rfile[15][14]),
    .dbg_bits_stateVec_15_rfile_15     (dbg_bits_stateVec_rfile[15][15]),
    .dbg_bits_stateVec_15_rfile_16     (dbg_bits_stateVec_rfile[15][16]),
    .dbg_bits_stateVec_15_rfile_17     (dbg_bits_stateVec_rfile[15][17]),
    .dbg_bits_stateVec_15_rfile_18     (dbg_bits_stateVec_rfile[15][18]),
    .dbg_bits_stateVec_15_rfile_19     (dbg_bits_stateVec_rfile[15][19]),
    .dbg_bits_stateVec_15_rfile_20     (dbg_bits_stateVec_rfile[15][20]),
    .dbg_bits_stateVec_15_rfile_21     (dbg_bits_stateVec_rfile[15][21]),
    .dbg_bits_stateVec_15_rfile_22     (dbg_bits_stateVec_rfile[15][22]),
    .dbg_bits_stateVec_15_rfile_23     (dbg_bits_stateVec_rfile[15][23]),
    .dbg_bits_stateVec_15_rfile_24     (dbg_bits_stateVec_rfile[15][24]),
    .dbg_bits_stateVec_15_rfile_25     (dbg_bits_stateVec_rfile[15][25]),
    .dbg_bits_stateVec_15_rfile_26     (dbg_bits_stateVec_rfile[15][26]),
    .dbg_bits_stateVec_15_rfile_27     (dbg_bits_stateVec_rfile[15][27]),
    .dbg_bits_stateVec_15_rfile_28     (dbg_bits_stateVec_rfile[15][28]),
    .dbg_bits_stateVec_15_rfile_29     (dbg_bits_stateVec_rfile[15][29]),
    .dbg_bits_stateVec_15_rfile_30     (dbg_bits_stateVec_rfile[15][30]),
    .dbg_bits_stateVec_15_rfile_31     (dbg_bits_stateVec_rfile[15][31]),
    .dbg_bits_stateVec_15_regs_PC      (dbg_bits_stateVec_regs_PC  [15]),
    .dbg_bits_stateVec_15_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[15]),
    .dbg_bits_stateVec_16_rfile_0      (dbg_bits_stateVec_rfile[16][0 ]),
    .dbg_bits_stateVec_16_rfile_1      (dbg_bits_stateVec_rfile[16][1 ]),
    .dbg_bits_stateVec_16_rfile_2      (dbg_bits_stateVec_rfile[16][2 ]),
    .dbg_bits_stateVec_16_rfile_3      (dbg_bits_stateVec_rfile[16][3 ]),
    .dbg_bits_stateVec_16_rfile_4      (dbg_bits_stateVec_rfile[16][4 ]),
    .dbg_bits_stateVec_16_rfile_5      (dbg_bits_stateVec_rfile[16][5 ]),
    .dbg_bits_stateVec_16_rfile_6      (dbg_bits_stateVec_rfile[16][6 ]),
    .dbg_bits_stateVec_16_rfile_7      (dbg_bits_stateVec_rfile[16][7 ]),
    .dbg_bits_stateVec_16_rfile_8      (dbg_bits_stateVec_rfile[16][8 ]),
    .dbg_bits_stateVec_16_rfile_9      (dbg_bits_stateVec_rfile[16][9 ]),
    .dbg_bits_stateVec_16_rfile_10     (dbg_bits_stateVec_rfile[16][10]),
    .dbg_bits_stateVec_16_rfile_11     (dbg_bits_stateVec_rfile[16][11]),
    .dbg_bits_stateVec_16_rfile_12     (dbg_bits_stateVec_rfile[16][12]),
    .dbg_bits_stateVec_16_rfile_13     (dbg_bits_stateVec_rfile[16][13]),
    .dbg_bits_stateVec_16_rfile_14     (dbg_bits_stateVec_rfile[16][14]),
    .dbg_bits_stateVec_16_rfile_15     (dbg_bits_stateVec_rfile[16][15]),
    .dbg_bits_stateVec_16_rfile_16     (dbg_bits_stateVec_rfile[16][16]),
    .dbg_bits_stateVec_16_rfile_17     (dbg_bits_stateVec_rfile[16][17]),
    .dbg_bits_stateVec_16_rfile_18     (dbg_bits_stateVec_rfile[16][18]),
    .dbg_bits_stateVec_16_rfile_19     (dbg_bits_stateVec_rfile[16][19]),
    .dbg_bits_stateVec_16_rfile_20     (dbg_bits_stateVec_rfile[16][20]),
    .dbg_bits_stateVec_16_rfile_21     (dbg_bits_stateVec_rfile[16][21]),
    .dbg_bits_stateVec_16_rfile_22     (dbg_bits_stateVec_rfile[16][22]),
    .dbg_bits_stateVec_16_rfile_23     (dbg_bits_stateVec_rfile[16][23]),
    .dbg_bits_stateVec_16_rfile_24     (dbg_bits_stateVec_rfile[16][24]),
    .dbg_bits_stateVec_16_rfile_25     (dbg_bits_stateVec_rfile[16][25]),
    .dbg_bits_stateVec_16_rfile_26     (dbg_bits_stateVec_rfile[16][26]),
    .dbg_bits_stateVec_16_rfile_27     (dbg_bits_stateVec_rfile[16][27]),
    .dbg_bits_stateVec_16_rfile_28     (dbg_bits_stateVec_rfile[16][28]),
    .dbg_bits_stateVec_16_rfile_29     (dbg_bits_stateVec_rfile[16][29]),
    .dbg_bits_stateVec_16_rfile_30     (dbg_bits_stateVec_rfile[16][30]),
    .dbg_bits_stateVec_16_rfile_31     (dbg_bits_stateVec_rfile[16][31]),
    .dbg_bits_stateVec_16_regs_PC      (dbg_bits_stateVec_regs_PC  [16]),
    .dbg_bits_stateVec_16_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[16]),
    .dbg_bits_stateVec_17_rfile_0      (dbg_bits_stateVec_rfile[17][0 ]),
    .dbg_bits_stateVec_17_rfile_1      (dbg_bits_stateVec_rfile[17][1 ]),
    .dbg_bits_stateVec_17_rfile_2      (dbg_bits_stateVec_rfile[17][2 ]),
    .dbg_bits_stateVec_17_rfile_3      (dbg_bits_stateVec_rfile[17][3 ]),
    .dbg_bits_stateVec_17_rfile_4      (dbg_bits_stateVec_rfile[17][4 ]),
    .dbg_bits_stateVec_17_rfile_5      (dbg_bits_stateVec_rfile[17][5 ]),
    .dbg_bits_stateVec_17_rfile_6      (dbg_bits_stateVec_rfile[17][6 ]),
    .dbg_bits_stateVec_17_rfile_7      (dbg_bits_stateVec_rfile[17][7 ]),
    .dbg_bits_stateVec_17_rfile_8      (dbg_bits_stateVec_rfile[17][8 ]),
    .dbg_bits_stateVec_17_rfile_9      (dbg_bits_stateVec_rfile[17][9 ]),
    .dbg_bits_stateVec_17_rfile_10     (dbg_bits_stateVec_rfile[17][10]),
    .dbg_bits_stateVec_17_rfile_11     (dbg_bits_stateVec_rfile[17][11]),
    .dbg_bits_stateVec_17_rfile_12     (dbg_bits_stateVec_rfile[17][12]),
    .dbg_bits_stateVec_17_rfile_13     (dbg_bits_stateVec_rfile[17][13]),
    .dbg_bits_stateVec_17_rfile_14     (dbg_bits_stateVec_rfile[17][14]),
    .dbg_bits_stateVec_17_rfile_15     (dbg_bits_stateVec_rfile[17][15]),
    .dbg_bits_stateVec_17_rfile_16     (dbg_bits_stateVec_rfile[17][16]),
    .dbg_bits_stateVec_17_rfile_17     (dbg_bits_stateVec_rfile[17][17]),
    .dbg_bits_stateVec_17_rfile_18     (dbg_bits_stateVec_rfile[17][18]),
    .dbg_bits_stateVec_17_rfile_19     (dbg_bits_stateVec_rfile[17][19]),
    .dbg_bits_stateVec_17_rfile_20     (dbg_bits_stateVec_rfile[17][20]),
    .dbg_bits_stateVec_17_rfile_21     (dbg_bits_stateVec_rfile[17][21]),
    .dbg_bits_stateVec_17_rfile_22     (dbg_bits_stateVec_rfile[17][22]),
    .dbg_bits_stateVec_17_rfile_23     (dbg_bits_stateVec_rfile[17][23]),
    .dbg_bits_stateVec_17_rfile_24     (dbg_bits_stateVec_rfile[17][24]),
    .dbg_bits_stateVec_17_rfile_25     (dbg_bits_stateVec_rfile[17][25]),
    .dbg_bits_stateVec_17_rfile_26     (dbg_bits_stateVec_rfile[17][26]),
    .dbg_bits_stateVec_17_rfile_27     (dbg_bits_stateVec_rfile[17][27]),
    .dbg_bits_stateVec_17_rfile_28     (dbg_bits_stateVec_rfile[17][28]),
    .dbg_bits_stateVec_17_rfile_29     (dbg_bits_stateVec_rfile[17][29]),
    .dbg_bits_stateVec_17_rfile_30     (dbg_bits_stateVec_rfile[17][30]),
    .dbg_bits_stateVec_17_rfile_31     (dbg_bits_stateVec_rfile[17][31]),
    .dbg_bits_stateVec_17_regs_PC      (dbg_bits_stateVec_regs_PC  [17]),
    .dbg_bits_stateVec_17_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[17]),
    .dbg_bits_stateVec_18_rfile_0      (dbg_bits_stateVec_rfile[18][0 ]),
    .dbg_bits_stateVec_18_rfile_1      (dbg_bits_stateVec_rfile[18][1 ]),
    .dbg_bits_stateVec_18_rfile_2      (dbg_bits_stateVec_rfile[18][2 ]),
    .dbg_bits_stateVec_18_rfile_3      (dbg_bits_stateVec_rfile[18][3 ]),
    .dbg_bits_stateVec_18_rfile_4      (dbg_bits_stateVec_rfile[18][4 ]),
    .dbg_bits_stateVec_18_rfile_5      (dbg_bits_stateVec_rfile[18][5 ]),
    .dbg_bits_stateVec_18_rfile_6      (dbg_bits_stateVec_rfile[18][6 ]),
    .dbg_bits_stateVec_18_rfile_7      (dbg_bits_stateVec_rfile[18][7 ]),
    .dbg_bits_stateVec_18_rfile_8      (dbg_bits_stateVec_rfile[18][8 ]),
    .dbg_bits_stateVec_18_rfile_9      (dbg_bits_stateVec_rfile[18][9 ]),
    .dbg_bits_stateVec_18_rfile_10     (dbg_bits_stateVec_rfile[18][10]),
    .dbg_bits_stateVec_18_rfile_11     (dbg_bits_stateVec_rfile[18][11]),
    .dbg_bits_stateVec_18_rfile_12     (dbg_bits_stateVec_rfile[18][12]),
    .dbg_bits_stateVec_18_rfile_13     (dbg_bits_stateVec_rfile[18][13]),
    .dbg_bits_stateVec_18_rfile_14     (dbg_bits_stateVec_rfile[18][14]),
    .dbg_bits_stateVec_18_rfile_15     (dbg_bits_stateVec_rfile[18][15]),
    .dbg_bits_stateVec_18_rfile_16     (dbg_bits_stateVec_rfile[18][16]),
    .dbg_bits_stateVec_18_rfile_17     (dbg_bits_stateVec_rfile[18][17]),
    .dbg_bits_stateVec_18_rfile_18     (dbg_bits_stateVec_rfile[18][18]),
    .dbg_bits_stateVec_18_rfile_19     (dbg_bits_stateVec_rfile[18][19]),
    .dbg_bits_stateVec_18_rfile_20     (dbg_bits_stateVec_rfile[18][20]),
    .dbg_bits_stateVec_18_rfile_21     (dbg_bits_stateVec_rfile[18][21]),
    .dbg_bits_stateVec_18_rfile_22     (dbg_bits_stateVec_rfile[18][22]),
    .dbg_bits_stateVec_18_rfile_23     (dbg_bits_stateVec_rfile[18][23]),
    .dbg_bits_stateVec_18_rfile_24     (dbg_bits_stateVec_rfile[18][24]),
    .dbg_bits_stateVec_18_rfile_25     (dbg_bits_stateVec_rfile[18][25]),
    .dbg_bits_stateVec_18_rfile_26     (dbg_bits_stateVec_rfile[18][26]),
    .dbg_bits_stateVec_18_rfile_27     (dbg_bits_stateVec_rfile[18][27]),
    .dbg_bits_stateVec_18_rfile_28     (dbg_bits_stateVec_rfile[18][28]),
    .dbg_bits_stateVec_18_rfile_29     (dbg_bits_stateVec_rfile[18][29]),
    .dbg_bits_stateVec_18_rfile_30     (dbg_bits_stateVec_rfile[18][30]),
    .dbg_bits_stateVec_18_rfile_31     (dbg_bits_stateVec_rfile[18][31]),
    .dbg_bits_stateVec_18_regs_PC      (dbg_bits_stateVec_regs_PC  [18]),
    .dbg_bits_stateVec_18_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[18]),
    .dbg_bits_stateVec_19_rfile_0      (dbg_bits_stateVec_rfile[19][0 ]),
    .dbg_bits_stateVec_19_rfile_1      (dbg_bits_stateVec_rfile[19][1 ]),
    .dbg_bits_stateVec_19_rfile_2      (dbg_bits_stateVec_rfile[19][2 ]),
    .dbg_bits_stateVec_19_rfile_3      (dbg_bits_stateVec_rfile[19][3 ]),
    .dbg_bits_stateVec_19_rfile_4      (dbg_bits_stateVec_rfile[19][4 ]),
    .dbg_bits_stateVec_19_rfile_5      (dbg_bits_stateVec_rfile[19][5 ]),
    .dbg_bits_stateVec_19_rfile_6      (dbg_bits_stateVec_rfile[19][6 ]),
    .dbg_bits_stateVec_19_rfile_7      (dbg_bits_stateVec_rfile[19][7 ]),
    .dbg_bits_stateVec_19_rfile_8      (dbg_bits_stateVec_rfile[19][8 ]),
    .dbg_bits_stateVec_19_rfile_9      (dbg_bits_stateVec_rfile[19][9 ]),
    .dbg_bits_stateVec_19_rfile_10     (dbg_bits_stateVec_rfile[19][10]),
    .dbg_bits_stateVec_19_rfile_11     (dbg_bits_stateVec_rfile[19][11]),
    .dbg_bits_stateVec_19_rfile_12     (dbg_bits_stateVec_rfile[19][12]),
    .dbg_bits_stateVec_19_rfile_13     (dbg_bits_stateVec_rfile[19][13]),
    .dbg_bits_stateVec_19_rfile_14     (dbg_bits_stateVec_rfile[19][14]),
    .dbg_bits_stateVec_19_rfile_15     (dbg_bits_stateVec_rfile[19][15]),
    .dbg_bits_stateVec_19_rfile_16     (dbg_bits_stateVec_rfile[19][16]),
    .dbg_bits_stateVec_19_rfile_17     (dbg_bits_stateVec_rfile[19][17]),
    .dbg_bits_stateVec_19_rfile_18     (dbg_bits_stateVec_rfile[19][18]),
    .dbg_bits_stateVec_19_rfile_19     (dbg_bits_stateVec_rfile[19][19]),
    .dbg_bits_stateVec_19_rfile_20     (dbg_bits_stateVec_rfile[19][20]),
    .dbg_bits_stateVec_19_rfile_21     (dbg_bits_stateVec_rfile[19][21]),
    .dbg_bits_stateVec_19_rfile_22     (dbg_bits_stateVec_rfile[19][22]),
    .dbg_bits_stateVec_19_rfile_23     (dbg_bits_stateVec_rfile[19][23]),
    .dbg_bits_stateVec_19_rfile_24     (dbg_bits_stateVec_rfile[19][24]),
    .dbg_bits_stateVec_19_rfile_25     (dbg_bits_stateVec_rfile[19][25]),
    .dbg_bits_stateVec_19_rfile_26     (dbg_bits_stateVec_rfile[19][26]),
    .dbg_bits_stateVec_19_rfile_27     (dbg_bits_stateVec_rfile[19][27]),
    .dbg_bits_stateVec_19_rfile_28     (dbg_bits_stateVec_rfile[19][28]),
    .dbg_bits_stateVec_19_rfile_29     (dbg_bits_stateVec_rfile[19][29]),
    .dbg_bits_stateVec_19_rfile_30     (dbg_bits_stateVec_rfile[19][30]),
    .dbg_bits_stateVec_19_rfile_31     (dbg_bits_stateVec_rfile[19][31]),
    .dbg_bits_stateVec_19_regs_PC      (dbg_bits_stateVec_regs_PC  [19]),
    .dbg_bits_stateVec_19_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[19]),
    .dbg_bits_stateVec_20_rfile_0      (dbg_bits_stateVec_rfile[20][0 ]),
    .dbg_bits_stateVec_20_rfile_1      (dbg_bits_stateVec_rfile[20][1 ]),
    .dbg_bits_stateVec_20_rfile_2      (dbg_bits_stateVec_rfile[20][2 ]),
    .dbg_bits_stateVec_20_rfile_3      (dbg_bits_stateVec_rfile[20][3 ]),
    .dbg_bits_stateVec_20_rfile_4      (dbg_bits_stateVec_rfile[20][4 ]),
    .dbg_bits_stateVec_20_rfile_5      (dbg_bits_stateVec_rfile[20][5 ]),
    .dbg_bits_stateVec_20_rfile_6      (dbg_bits_stateVec_rfile[20][6 ]),
    .dbg_bits_stateVec_20_rfile_7      (dbg_bits_stateVec_rfile[20][7 ]),
    .dbg_bits_stateVec_20_rfile_8      (dbg_bits_stateVec_rfile[20][8 ]),
    .dbg_bits_stateVec_20_rfile_9      (dbg_bits_stateVec_rfile[20][9 ]),
    .dbg_bits_stateVec_20_rfile_10     (dbg_bits_stateVec_rfile[20][10]),
    .dbg_bits_stateVec_20_rfile_11     (dbg_bits_stateVec_rfile[20][11]),
    .dbg_bits_stateVec_20_rfile_12     (dbg_bits_stateVec_rfile[20][12]),
    .dbg_bits_stateVec_20_rfile_13     (dbg_bits_stateVec_rfile[20][13]),
    .dbg_bits_stateVec_20_rfile_14     (dbg_bits_stateVec_rfile[20][14]),
    .dbg_bits_stateVec_20_rfile_15     (dbg_bits_stateVec_rfile[20][15]),
    .dbg_bits_stateVec_20_rfile_16     (dbg_bits_stateVec_rfile[20][16]),
    .dbg_bits_stateVec_20_rfile_17     (dbg_bits_stateVec_rfile[20][17]),
    .dbg_bits_stateVec_20_rfile_18     (dbg_bits_stateVec_rfile[20][18]),
    .dbg_bits_stateVec_20_rfile_19     (dbg_bits_stateVec_rfile[20][19]),
    .dbg_bits_stateVec_20_rfile_20     (dbg_bits_stateVec_rfile[20][20]),
    .dbg_bits_stateVec_20_rfile_21     (dbg_bits_stateVec_rfile[20][21]),
    .dbg_bits_stateVec_20_rfile_22     (dbg_bits_stateVec_rfile[20][22]),
    .dbg_bits_stateVec_20_rfile_23     (dbg_bits_stateVec_rfile[20][23]),
    .dbg_bits_stateVec_20_rfile_24     (dbg_bits_stateVec_rfile[20][24]),
    .dbg_bits_stateVec_20_rfile_25     (dbg_bits_stateVec_rfile[20][25]),
    .dbg_bits_stateVec_20_rfile_26     (dbg_bits_stateVec_rfile[20][26]),
    .dbg_bits_stateVec_20_rfile_27     (dbg_bits_stateVec_rfile[20][27]),
    .dbg_bits_stateVec_20_rfile_28     (dbg_bits_stateVec_rfile[20][28]),
    .dbg_bits_stateVec_20_rfile_29     (dbg_bits_stateVec_rfile[20][29]),
    .dbg_bits_stateVec_20_rfile_30     (dbg_bits_stateVec_rfile[20][30]),
    .dbg_bits_stateVec_20_rfile_31     (dbg_bits_stateVec_rfile[20][31]),
    .dbg_bits_stateVec_20_regs_PC      (dbg_bits_stateVec_regs_PC  [20]),
    .dbg_bits_stateVec_20_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[20]),
    .dbg_bits_stateVec_21_rfile_0      (dbg_bits_stateVec_rfile[21][0 ]),
    .dbg_bits_stateVec_21_rfile_1      (dbg_bits_stateVec_rfile[21][1 ]),
    .dbg_bits_stateVec_21_rfile_2      (dbg_bits_stateVec_rfile[21][2 ]),
    .dbg_bits_stateVec_21_rfile_3      (dbg_bits_stateVec_rfile[21][3 ]),
    .dbg_bits_stateVec_21_rfile_4      (dbg_bits_stateVec_rfile[21][4 ]),
    .dbg_bits_stateVec_21_rfile_5      (dbg_bits_stateVec_rfile[21][5 ]),
    .dbg_bits_stateVec_21_rfile_6      (dbg_bits_stateVec_rfile[21][6 ]),
    .dbg_bits_stateVec_21_rfile_7      (dbg_bits_stateVec_rfile[21][7 ]),
    .dbg_bits_stateVec_21_rfile_8      (dbg_bits_stateVec_rfile[21][8 ]),
    .dbg_bits_stateVec_21_rfile_9      (dbg_bits_stateVec_rfile[21][9 ]),
    .dbg_bits_stateVec_21_rfile_10     (dbg_bits_stateVec_rfile[21][10]),
    .dbg_bits_stateVec_21_rfile_11     (dbg_bits_stateVec_rfile[21][11]),
    .dbg_bits_stateVec_21_rfile_12     (dbg_bits_stateVec_rfile[21][12]),
    .dbg_bits_stateVec_21_rfile_13     (dbg_bits_stateVec_rfile[21][13]),
    .dbg_bits_stateVec_21_rfile_14     (dbg_bits_stateVec_rfile[21][14]),
    .dbg_bits_stateVec_21_rfile_15     (dbg_bits_stateVec_rfile[21][15]),
    .dbg_bits_stateVec_21_rfile_16     (dbg_bits_stateVec_rfile[21][16]),
    .dbg_bits_stateVec_21_rfile_17     (dbg_bits_stateVec_rfile[21][17]),
    .dbg_bits_stateVec_21_rfile_18     (dbg_bits_stateVec_rfile[21][18]),
    .dbg_bits_stateVec_21_rfile_19     (dbg_bits_stateVec_rfile[21][19]),
    .dbg_bits_stateVec_21_rfile_20     (dbg_bits_stateVec_rfile[21][20]),
    .dbg_bits_stateVec_21_rfile_21     (dbg_bits_stateVec_rfile[21][21]),
    .dbg_bits_stateVec_21_rfile_22     (dbg_bits_stateVec_rfile[21][22]),
    .dbg_bits_stateVec_21_rfile_23     (dbg_bits_stateVec_rfile[21][23]),
    .dbg_bits_stateVec_21_rfile_24     (dbg_bits_stateVec_rfile[21][24]),
    .dbg_bits_stateVec_21_rfile_25     (dbg_bits_stateVec_rfile[21][25]),
    .dbg_bits_stateVec_21_rfile_26     (dbg_bits_stateVec_rfile[21][26]),
    .dbg_bits_stateVec_21_rfile_27     (dbg_bits_stateVec_rfile[21][27]),
    .dbg_bits_stateVec_21_rfile_28     (dbg_bits_stateVec_rfile[21][28]),
    .dbg_bits_stateVec_21_rfile_29     (dbg_bits_stateVec_rfile[21][29]),
    .dbg_bits_stateVec_21_rfile_30     (dbg_bits_stateVec_rfile[21][30]),
    .dbg_bits_stateVec_21_rfile_31     (dbg_bits_stateVec_rfile[21][31]),
    .dbg_bits_stateVec_21_regs_PC      (dbg_bits_stateVec_regs_PC  [21]),
    .dbg_bits_stateVec_21_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[21]),
    .dbg_bits_stateVec_22_rfile_0      (dbg_bits_stateVec_rfile[22][0 ]),
    .dbg_bits_stateVec_22_rfile_1      (dbg_bits_stateVec_rfile[22][1 ]),
    .dbg_bits_stateVec_22_rfile_2      (dbg_bits_stateVec_rfile[22][2 ]),
    .dbg_bits_stateVec_22_rfile_3      (dbg_bits_stateVec_rfile[22][3 ]),
    .dbg_bits_stateVec_22_rfile_4      (dbg_bits_stateVec_rfile[22][4 ]),
    .dbg_bits_stateVec_22_rfile_5      (dbg_bits_stateVec_rfile[22][5 ]),
    .dbg_bits_stateVec_22_rfile_6      (dbg_bits_stateVec_rfile[22][6 ]),
    .dbg_bits_stateVec_22_rfile_7      (dbg_bits_stateVec_rfile[22][7 ]),
    .dbg_bits_stateVec_22_rfile_8      (dbg_bits_stateVec_rfile[22][8 ]),
    .dbg_bits_stateVec_22_rfile_9      (dbg_bits_stateVec_rfile[22][9 ]),
    .dbg_bits_stateVec_22_rfile_10     (dbg_bits_stateVec_rfile[22][10]),
    .dbg_bits_stateVec_22_rfile_11     (dbg_bits_stateVec_rfile[22][11]),
    .dbg_bits_stateVec_22_rfile_12     (dbg_bits_stateVec_rfile[22][12]),
    .dbg_bits_stateVec_22_rfile_13     (dbg_bits_stateVec_rfile[22][13]),
    .dbg_bits_stateVec_22_rfile_14     (dbg_bits_stateVec_rfile[22][14]),
    .dbg_bits_stateVec_22_rfile_15     (dbg_bits_stateVec_rfile[22][15]),
    .dbg_bits_stateVec_22_rfile_16     (dbg_bits_stateVec_rfile[22][16]),
    .dbg_bits_stateVec_22_rfile_17     (dbg_bits_stateVec_rfile[22][17]),
    .dbg_bits_stateVec_22_rfile_18     (dbg_bits_stateVec_rfile[22][18]),
    .dbg_bits_stateVec_22_rfile_19     (dbg_bits_stateVec_rfile[22][19]),
    .dbg_bits_stateVec_22_rfile_20     (dbg_bits_stateVec_rfile[22][20]),
    .dbg_bits_stateVec_22_rfile_21     (dbg_bits_stateVec_rfile[22][21]),
    .dbg_bits_stateVec_22_rfile_22     (dbg_bits_stateVec_rfile[22][22]),
    .dbg_bits_stateVec_22_rfile_23     (dbg_bits_stateVec_rfile[22][23]),
    .dbg_bits_stateVec_22_rfile_24     (dbg_bits_stateVec_rfile[22][24]),
    .dbg_bits_stateVec_22_rfile_25     (dbg_bits_stateVec_rfile[22][25]),
    .dbg_bits_stateVec_22_rfile_26     (dbg_bits_stateVec_rfile[22][26]),
    .dbg_bits_stateVec_22_rfile_27     (dbg_bits_stateVec_rfile[22][27]),
    .dbg_bits_stateVec_22_rfile_28     (dbg_bits_stateVec_rfile[22][28]),
    .dbg_bits_stateVec_22_rfile_29     (dbg_bits_stateVec_rfile[22][29]),
    .dbg_bits_stateVec_22_rfile_30     (dbg_bits_stateVec_rfile[22][30]),
    .dbg_bits_stateVec_22_rfile_31     (dbg_bits_stateVec_rfile[22][31]),
    .dbg_bits_stateVec_22_regs_PC      (dbg_bits_stateVec_regs_PC  [22]),
    .dbg_bits_stateVec_22_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[22]),
    .dbg_bits_stateVec_23_rfile_0      (dbg_bits_stateVec_rfile[23][0 ]),
    .dbg_bits_stateVec_23_rfile_1      (dbg_bits_stateVec_rfile[23][1 ]),
    .dbg_bits_stateVec_23_rfile_2      (dbg_bits_stateVec_rfile[23][2 ]),
    .dbg_bits_stateVec_23_rfile_3      (dbg_bits_stateVec_rfile[23][3 ]),
    .dbg_bits_stateVec_23_rfile_4      (dbg_bits_stateVec_rfile[23][4 ]),
    .dbg_bits_stateVec_23_rfile_5      (dbg_bits_stateVec_rfile[23][5 ]),
    .dbg_bits_stateVec_23_rfile_6      (dbg_bits_stateVec_rfile[23][6 ]),
    .dbg_bits_stateVec_23_rfile_7      (dbg_bits_stateVec_rfile[23][7 ]),
    .dbg_bits_stateVec_23_rfile_8      (dbg_bits_stateVec_rfile[23][8 ]),
    .dbg_bits_stateVec_23_rfile_9      (dbg_bits_stateVec_rfile[23][9 ]),
    .dbg_bits_stateVec_23_rfile_10     (dbg_bits_stateVec_rfile[23][10]),
    .dbg_bits_stateVec_23_rfile_11     (dbg_bits_stateVec_rfile[23][11]),
    .dbg_bits_stateVec_23_rfile_12     (dbg_bits_stateVec_rfile[23][12]),
    .dbg_bits_stateVec_23_rfile_13     (dbg_bits_stateVec_rfile[23][13]),
    .dbg_bits_stateVec_23_rfile_14     (dbg_bits_stateVec_rfile[23][14]),
    .dbg_bits_stateVec_23_rfile_15     (dbg_bits_stateVec_rfile[23][15]),
    .dbg_bits_stateVec_23_rfile_16     (dbg_bits_stateVec_rfile[23][16]),
    .dbg_bits_stateVec_23_rfile_17     (dbg_bits_stateVec_rfile[23][17]),
    .dbg_bits_stateVec_23_rfile_18     (dbg_bits_stateVec_rfile[23][18]),
    .dbg_bits_stateVec_23_rfile_19     (dbg_bits_stateVec_rfile[23][19]),
    .dbg_bits_stateVec_23_rfile_20     (dbg_bits_stateVec_rfile[23][20]),
    .dbg_bits_stateVec_23_rfile_21     (dbg_bits_stateVec_rfile[23][21]),
    .dbg_bits_stateVec_23_rfile_22     (dbg_bits_stateVec_rfile[23][22]),
    .dbg_bits_stateVec_23_rfile_23     (dbg_bits_stateVec_rfile[23][23]),
    .dbg_bits_stateVec_23_rfile_24     (dbg_bits_stateVec_rfile[23][24]),
    .dbg_bits_stateVec_23_rfile_25     (dbg_bits_stateVec_rfile[23][25]),
    .dbg_bits_stateVec_23_rfile_26     (dbg_bits_stateVec_rfile[23][26]),
    .dbg_bits_stateVec_23_rfile_27     (dbg_bits_stateVec_rfile[23][27]),
    .dbg_bits_stateVec_23_rfile_28     (dbg_bits_stateVec_rfile[23][28]),
    .dbg_bits_stateVec_23_rfile_29     (dbg_bits_stateVec_rfile[23][29]),
    .dbg_bits_stateVec_23_rfile_30     (dbg_bits_stateVec_rfile[23][30]),
    .dbg_bits_stateVec_23_rfile_31     (dbg_bits_stateVec_rfile[23][31]),
    .dbg_bits_stateVec_23_regs_PC      (dbg_bits_stateVec_regs_PC  [23]),
    .dbg_bits_stateVec_23_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[23]),
    .dbg_bits_stateVec_24_rfile_0      (dbg_bits_stateVec_rfile[24][0 ]),
    .dbg_bits_stateVec_24_rfile_1      (dbg_bits_stateVec_rfile[24][1 ]),
    .dbg_bits_stateVec_24_rfile_2      (dbg_bits_stateVec_rfile[24][2 ]),
    .dbg_bits_stateVec_24_rfile_3      (dbg_bits_stateVec_rfile[24][3 ]),
    .dbg_bits_stateVec_24_rfile_4      (dbg_bits_stateVec_rfile[24][4 ]),
    .dbg_bits_stateVec_24_rfile_5      (dbg_bits_stateVec_rfile[24][5 ]),
    .dbg_bits_stateVec_24_rfile_6      (dbg_bits_stateVec_rfile[24][6 ]),
    .dbg_bits_stateVec_24_rfile_7      (dbg_bits_stateVec_rfile[24][7 ]),
    .dbg_bits_stateVec_24_rfile_8      (dbg_bits_stateVec_rfile[24][8 ]),
    .dbg_bits_stateVec_24_rfile_9      (dbg_bits_stateVec_rfile[24][9 ]),
    .dbg_bits_stateVec_24_rfile_10     (dbg_bits_stateVec_rfile[24][10]),
    .dbg_bits_stateVec_24_rfile_11     (dbg_bits_stateVec_rfile[24][11]),
    .dbg_bits_stateVec_24_rfile_12     (dbg_bits_stateVec_rfile[24][12]),
    .dbg_bits_stateVec_24_rfile_13     (dbg_bits_stateVec_rfile[24][13]),
    .dbg_bits_stateVec_24_rfile_14     (dbg_bits_stateVec_rfile[24][14]),
    .dbg_bits_stateVec_24_rfile_15     (dbg_bits_stateVec_rfile[24][15]),
    .dbg_bits_stateVec_24_rfile_16     (dbg_bits_stateVec_rfile[24][16]),
    .dbg_bits_stateVec_24_rfile_17     (dbg_bits_stateVec_rfile[24][17]),
    .dbg_bits_stateVec_24_rfile_18     (dbg_bits_stateVec_rfile[24][18]),
    .dbg_bits_stateVec_24_rfile_19     (dbg_bits_stateVec_rfile[24][19]),
    .dbg_bits_stateVec_24_rfile_20     (dbg_bits_stateVec_rfile[24][20]),
    .dbg_bits_stateVec_24_rfile_21     (dbg_bits_stateVec_rfile[24][21]),
    .dbg_bits_stateVec_24_rfile_22     (dbg_bits_stateVec_rfile[24][22]),
    .dbg_bits_stateVec_24_rfile_23     (dbg_bits_stateVec_rfile[24][23]),
    .dbg_bits_stateVec_24_rfile_24     (dbg_bits_stateVec_rfile[24][24]),
    .dbg_bits_stateVec_24_rfile_25     (dbg_bits_stateVec_rfile[24][25]),
    .dbg_bits_stateVec_24_rfile_26     (dbg_bits_stateVec_rfile[24][26]),
    .dbg_bits_stateVec_24_rfile_27     (dbg_bits_stateVec_rfile[24][27]),
    .dbg_bits_stateVec_24_rfile_28     (dbg_bits_stateVec_rfile[24][28]),
    .dbg_bits_stateVec_24_rfile_29     (dbg_bits_stateVec_rfile[24][29]),
    .dbg_bits_stateVec_24_rfile_30     (dbg_bits_stateVec_rfile[24][30]),
    .dbg_bits_stateVec_24_rfile_31     (dbg_bits_stateVec_rfile[24][31]),
    .dbg_bits_stateVec_24_regs_PC      (dbg_bits_stateVec_regs_PC  [24]),
    .dbg_bits_stateVec_24_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[24]),
    .dbg_bits_stateVec_25_rfile_0      (dbg_bits_stateVec_rfile[25][0 ]),
    .dbg_bits_stateVec_25_rfile_1      (dbg_bits_stateVec_rfile[25][1 ]),
    .dbg_bits_stateVec_25_rfile_2      (dbg_bits_stateVec_rfile[25][2 ]),
    .dbg_bits_stateVec_25_rfile_3      (dbg_bits_stateVec_rfile[25][3 ]),
    .dbg_bits_stateVec_25_rfile_4      (dbg_bits_stateVec_rfile[25][4 ]),
    .dbg_bits_stateVec_25_rfile_5      (dbg_bits_stateVec_rfile[25][5 ]),
    .dbg_bits_stateVec_25_rfile_6      (dbg_bits_stateVec_rfile[25][6 ]),
    .dbg_bits_stateVec_25_rfile_7      (dbg_bits_stateVec_rfile[25][7 ]),
    .dbg_bits_stateVec_25_rfile_8      (dbg_bits_stateVec_rfile[25][8 ]),
    .dbg_bits_stateVec_25_rfile_9      (dbg_bits_stateVec_rfile[25][9 ]),
    .dbg_bits_stateVec_25_rfile_10     (dbg_bits_stateVec_rfile[25][10]),
    .dbg_bits_stateVec_25_rfile_11     (dbg_bits_stateVec_rfile[25][11]),
    .dbg_bits_stateVec_25_rfile_12     (dbg_bits_stateVec_rfile[25][12]),
    .dbg_bits_stateVec_25_rfile_13     (dbg_bits_stateVec_rfile[25][13]),
    .dbg_bits_stateVec_25_rfile_14     (dbg_bits_stateVec_rfile[25][14]),
    .dbg_bits_stateVec_25_rfile_15     (dbg_bits_stateVec_rfile[25][15]),
    .dbg_bits_stateVec_25_rfile_16     (dbg_bits_stateVec_rfile[25][16]),
    .dbg_bits_stateVec_25_rfile_17     (dbg_bits_stateVec_rfile[25][17]),
    .dbg_bits_stateVec_25_rfile_18     (dbg_bits_stateVec_rfile[25][18]),
    .dbg_bits_stateVec_25_rfile_19     (dbg_bits_stateVec_rfile[25][19]),
    .dbg_bits_stateVec_25_rfile_20     (dbg_bits_stateVec_rfile[25][20]),
    .dbg_bits_stateVec_25_rfile_21     (dbg_bits_stateVec_rfile[25][21]),
    .dbg_bits_stateVec_25_rfile_22     (dbg_bits_stateVec_rfile[25][22]),
    .dbg_bits_stateVec_25_rfile_23     (dbg_bits_stateVec_rfile[25][23]),
    .dbg_bits_stateVec_25_rfile_24     (dbg_bits_stateVec_rfile[25][24]),
    .dbg_bits_stateVec_25_rfile_25     (dbg_bits_stateVec_rfile[25][25]),
    .dbg_bits_stateVec_25_rfile_26     (dbg_bits_stateVec_rfile[25][26]),
    .dbg_bits_stateVec_25_rfile_27     (dbg_bits_stateVec_rfile[25][27]),
    .dbg_bits_stateVec_25_rfile_28     (dbg_bits_stateVec_rfile[25][28]),
    .dbg_bits_stateVec_25_rfile_29     (dbg_bits_stateVec_rfile[25][29]),
    .dbg_bits_stateVec_25_rfile_30     (dbg_bits_stateVec_rfile[25][30]),
    .dbg_bits_stateVec_25_rfile_31     (dbg_bits_stateVec_rfile[25][31]),
    .dbg_bits_stateVec_25_regs_PC      (dbg_bits_stateVec_regs_PC  [25]),
    .dbg_bits_stateVec_25_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[25]),
    .dbg_bits_stateVec_26_rfile_0      (dbg_bits_stateVec_rfile[26][0 ]),
    .dbg_bits_stateVec_26_rfile_1      (dbg_bits_stateVec_rfile[26][1 ]),
    .dbg_bits_stateVec_26_rfile_2      (dbg_bits_stateVec_rfile[26][2 ]),
    .dbg_bits_stateVec_26_rfile_3      (dbg_bits_stateVec_rfile[26][3 ]),
    .dbg_bits_stateVec_26_rfile_4      (dbg_bits_stateVec_rfile[26][4 ]),
    .dbg_bits_stateVec_26_rfile_5      (dbg_bits_stateVec_rfile[26][5 ]),
    .dbg_bits_stateVec_26_rfile_6      (dbg_bits_stateVec_rfile[26][6 ]),
    .dbg_bits_stateVec_26_rfile_7      (dbg_bits_stateVec_rfile[26][7 ]),
    .dbg_bits_stateVec_26_rfile_8      (dbg_bits_stateVec_rfile[26][8 ]),
    .dbg_bits_stateVec_26_rfile_9      (dbg_bits_stateVec_rfile[26][9 ]),
    .dbg_bits_stateVec_26_rfile_10     (dbg_bits_stateVec_rfile[26][10]),
    .dbg_bits_stateVec_26_rfile_11     (dbg_bits_stateVec_rfile[26][11]),
    .dbg_bits_stateVec_26_rfile_12     (dbg_bits_stateVec_rfile[26][12]),
    .dbg_bits_stateVec_26_rfile_13     (dbg_bits_stateVec_rfile[26][13]),
    .dbg_bits_stateVec_26_rfile_14     (dbg_bits_stateVec_rfile[26][14]),
    .dbg_bits_stateVec_26_rfile_15     (dbg_bits_stateVec_rfile[26][15]),
    .dbg_bits_stateVec_26_rfile_16     (dbg_bits_stateVec_rfile[26][16]),
    .dbg_bits_stateVec_26_rfile_17     (dbg_bits_stateVec_rfile[26][17]),
    .dbg_bits_stateVec_26_rfile_18     (dbg_bits_stateVec_rfile[26][18]),
    .dbg_bits_stateVec_26_rfile_19     (dbg_bits_stateVec_rfile[26][19]),
    .dbg_bits_stateVec_26_rfile_20     (dbg_bits_stateVec_rfile[26][20]),
    .dbg_bits_stateVec_26_rfile_21     (dbg_bits_stateVec_rfile[26][21]),
    .dbg_bits_stateVec_26_rfile_22     (dbg_bits_stateVec_rfile[26][22]),
    .dbg_bits_stateVec_26_rfile_23     (dbg_bits_stateVec_rfile[26][23]),
    .dbg_bits_stateVec_26_rfile_24     (dbg_bits_stateVec_rfile[26][24]),
    .dbg_bits_stateVec_26_rfile_25     (dbg_bits_stateVec_rfile[26][25]),
    .dbg_bits_stateVec_26_rfile_26     (dbg_bits_stateVec_rfile[26][26]),
    .dbg_bits_stateVec_26_rfile_27     (dbg_bits_stateVec_rfile[26][27]),
    .dbg_bits_stateVec_26_rfile_28     (dbg_bits_stateVec_rfile[26][28]),
    .dbg_bits_stateVec_26_rfile_29     (dbg_bits_stateVec_rfile[26][29]),
    .dbg_bits_stateVec_26_rfile_30     (dbg_bits_stateVec_rfile[26][30]),
    .dbg_bits_stateVec_26_rfile_31     (dbg_bits_stateVec_rfile[26][31]),
    .dbg_bits_stateVec_26_regs_PC      (dbg_bits_stateVec_regs_PC  [26]),
    .dbg_bits_stateVec_26_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[26]),
    .dbg_bits_stateVec_27_rfile_0      (dbg_bits_stateVec_rfile[27][0 ]),
    .dbg_bits_stateVec_27_rfile_1      (dbg_bits_stateVec_rfile[27][1 ]),
    .dbg_bits_stateVec_27_rfile_2      (dbg_bits_stateVec_rfile[27][2 ]),
    .dbg_bits_stateVec_27_rfile_3      (dbg_bits_stateVec_rfile[27][3 ]),
    .dbg_bits_stateVec_27_rfile_4      (dbg_bits_stateVec_rfile[27][4 ]),
    .dbg_bits_stateVec_27_rfile_5      (dbg_bits_stateVec_rfile[27][5 ]),
    .dbg_bits_stateVec_27_rfile_6      (dbg_bits_stateVec_rfile[27][6 ]),
    .dbg_bits_stateVec_27_rfile_7      (dbg_bits_stateVec_rfile[27][7 ]),
    .dbg_bits_stateVec_27_rfile_8      (dbg_bits_stateVec_rfile[27][8 ]),
    .dbg_bits_stateVec_27_rfile_9      (dbg_bits_stateVec_rfile[27][9 ]),
    .dbg_bits_stateVec_27_rfile_10     (dbg_bits_stateVec_rfile[27][10]),
    .dbg_bits_stateVec_27_rfile_11     (dbg_bits_stateVec_rfile[27][11]),
    .dbg_bits_stateVec_27_rfile_12     (dbg_bits_stateVec_rfile[27][12]),
    .dbg_bits_stateVec_27_rfile_13     (dbg_bits_stateVec_rfile[27][13]),
    .dbg_bits_stateVec_27_rfile_14     (dbg_bits_stateVec_rfile[27][14]),
    .dbg_bits_stateVec_27_rfile_15     (dbg_bits_stateVec_rfile[27][15]),
    .dbg_bits_stateVec_27_rfile_16     (dbg_bits_stateVec_rfile[27][16]),
    .dbg_bits_stateVec_27_rfile_17     (dbg_bits_stateVec_rfile[27][17]),
    .dbg_bits_stateVec_27_rfile_18     (dbg_bits_stateVec_rfile[27][18]),
    .dbg_bits_stateVec_27_rfile_19     (dbg_bits_stateVec_rfile[27][19]),
    .dbg_bits_stateVec_27_rfile_20     (dbg_bits_stateVec_rfile[27][20]),
    .dbg_bits_stateVec_27_rfile_21     (dbg_bits_stateVec_rfile[27][21]),
    .dbg_bits_stateVec_27_rfile_22     (dbg_bits_stateVec_rfile[27][22]),
    .dbg_bits_stateVec_27_rfile_23     (dbg_bits_stateVec_rfile[27][23]),
    .dbg_bits_stateVec_27_rfile_24     (dbg_bits_stateVec_rfile[27][24]),
    .dbg_bits_stateVec_27_rfile_25     (dbg_bits_stateVec_rfile[27][25]),
    .dbg_bits_stateVec_27_rfile_26     (dbg_bits_stateVec_rfile[27][26]),
    .dbg_bits_stateVec_27_rfile_27     (dbg_bits_stateVec_rfile[27][27]),
    .dbg_bits_stateVec_27_rfile_28     (dbg_bits_stateVec_rfile[27][28]),
    .dbg_bits_stateVec_27_rfile_29     (dbg_bits_stateVec_rfile[27][29]),
    .dbg_bits_stateVec_27_rfile_30     (dbg_bits_stateVec_rfile[27][30]),
    .dbg_bits_stateVec_27_rfile_31     (dbg_bits_stateVec_rfile[27][31]),
    .dbg_bits_stateVec_27_regs_PC      (dbg_bits_stateVec_regs_PC  [27]),
    .dbg_bits_stateVec_27_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[27]),
    .dbg_bits_stateVec_28_rfile_0      (dbg_bits_stateVec_rfile[28][0 ]),
    .dbg_bits_stateVec_28_rfile_1      (dbg_bits_stateVec_rfile[28][1 ]),
    .dbg_bits_stateVec_28_rfile_2      (dbg_bits_stateVec_rfile[28][2 ]),
    .dbg_bits_stateVec_28_rfile_3      (dbg_bits_stateVec_rfile[28][3 ]),
    .dbg_bits_stateVec_28_rfile_4      (dbg_bits_stateVec_rfile[28][4 ]),
    .dbg_bits_stateVec_28_rfile_5      (dbg_bits_stateVec_rfile[28][5 ]),
    .dbg_bits_stateVec_28_rfile_6      (dbg_bits_stateVec_rfile[28][6 ]),
    .dbg_bits_stateVec_28_rfile_7      (dbg_bits_stateVec_rfile[28][7 ]),
    .dbg_bits_stateVec_28_rfile_8      (dbg_bits_stateVec_rfile[28][8 ]),
    .dbg_bits_stateVec_28_rfile_9      (dbg_bits_stateVec_rfile[28][9 ]),
    .dbg_bits_stateVec_28_rfile_10     (dbg_bits_stateVec_rfile[28][10]),
    .dbg_bits_stateVec_28_rfile_11     (dbg_bits_stateVec_rfile[28][11]),
    .dbg_bits_stateVec_28_rfile_12     (dbg_bits_stateVec_rfile[28][12]),
    .dbg_bits_stateVec_28_rfile_13     (dbg_bits_stateVec_rfile[28][13]),
    .dbg_bits_stateVec_28_rfile_14     (dbg_bits_stateVec_rfile[28][14]),
    .dbg_bits_stateVec_28_rfile_15     (dbg_bits_stateVec_rfile[28][15]),
    .dbg_bits_stateVec_28_rfile_16     (dbg_bits_stateVec_rfile[28][16]),
    .dbg_bits_stateVec_28_rfile_17     (dbg_bits_stateVec_rfile[28][17]),
    .dbg_bits_stateVec_28_rfile_18     (dbg_bits_stateVec_rfile[28][18]),
    .dbg_bits_stateVec_28_rfile_19     (dbg_bits_stateVec_rfile[28][19]),
    .dbg_bits_stateVec_28_rfile_20     (dbg_bits_stateVec_rfile[28][20]),
    .dbg_bits_stateVec_28_rfile_21     (dbg_bits_stateVec_rfile[28][21]),
    .dbg_bits_stateVec_28_rfile_22     (dbg_bits_stateVec_rfile[28][22]),
    .dbg_bits_stateVec_28_rfile_23     (dbg_bits_stateVec_rfile[28][23]),
    .dbg_bits_stateVec_28_rfile_24     (dbg_bits_stateVec_rfile[28][24]),
    .dbg_bits_stateVec_28_rfile_25     (dbg_bits_stateVec_rfile[28][25]),
    .dbg_bits_stateVec_28_rfile_26     (dbg_bits_stateVec_rfile[28][26]),
    .dbg_bits_stateVec_28_rfile_27     (dbg_bits_stateVec_rfile[28][27]),
    .dbg_bits_stateVec_28_rfile_28     (dbg_bits_stateVec_rfile[28][28]),
    .dbg_bits_stateVec_28_rfile_29     (dbg_bits_stateVec_rfile[28][29]),
    .dbg_bits_stateVec_28_rfile_30     (dbg_bits_stateVec_rfile[28][30]),
    .dbg_bits_stateVec_28_rfile_31     (dbg_bits_stateVec_rfile[28][31]),
    .dbg_bits_stateVec_28_regs_PC      (dbg_bits_stateVec_regs_PC  [28]),
    .dbg_bits_stateVec_28_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[28]),
    .dbg_bits_stateVec_29_rfile_0      (dbg_bits_stateVec_rfile[29][0 ]),
    .dbg_bits_stateVec_29_rfile_1      (dbg_bits_stateVec_rfile[29][1 ]),
    .dbg_bits_stateVec_29_rfile_2      (dbg_bits_stateVec_rfile[29][2 ]),
    .dbg_bits_stateVec_29_rfile_3      (dbg_bits_stateVec_rfile[29][3 ]),
    .dbg_bits_stateVec_29_rfile_4      (dbg_bits_stateVec_rfile[29][4 ]),
    .dbg_bits_stateVec_29_rfile_5      (dbg_bits_stateVec_rfile[29][5 ]),
    .dbg_bits_stateVec_29_rfile_6      (dbg_bits_stateVec_rfile[29][6 ]),
    .dbg_bits_stateVec_29_rfile_7      (dbg_bits_stateVec_rfile[29][7 ]),
    .dbg_bits_stateVec_29_rfile_8      (dbg_bits_stateVec_rfile[29][8 ]),
    .dbg_bits_stateVec_29_rfile_9      (dbg_bits_stateVec_rfile[29][9 ]),
    .dbg_bits_stateVec_29_rfile_10     (dbg_bits_stateVec_rfile[29][10]),
    .dbg_bits_stateVec_29_rfile_11     (dbg_bits_stateVec_rfile[29][11]),
    .dbg_bits_stateVec_29_rfile_12     (dbg_bits_stateVec_rfile[29][12]),
    .dbg_bits_stateVec_29_rfile_13     (dbg_bits_stateVec_rfile[29][13]),
    .dbg_bits_stateVec_29_rfile_14     (dbg_bits_stateVec_rfile[29][14]),
    .dbg_bits_stateVec_29_rfile_15     (dbg_bits_stateVec_rfile[29][15]),
    .dbg_bits_stateVec_29_rfile_16     (dbg_bits_stateVec_rfile[29][16]),
    .dbg_bits_stateVec_29_rfile_17     (dbg_bits_stateVec_rfile[29][17]),
    .dbg_bits_stateVec_29_rfile_18     (dbg_bits_stateVec_rfile[29][18]),
    .dbg_bits_stateVec_29_rfile_19     (dbg_bits_stateVec_rfile[29][19]),
    .dbg_bits_stateVec_29_rfile_20     (dbg_bits_stateVec_rfile[29][20]),
    .dbg_bits_stateVec_29_rfile_21     (dbg_bits_stateVec_rfile[29][21]),
    .dbg_bits_stateVec_29_rfile_22     (dbg_bits_stateVec_rfile[29][22]),
    .dbg_bits_stateVec_29_rfile_23     (dbg_bits_stateVec_rfile[29][23]),
    .dbg_bits_stateVec_29_rfile_24     (dbg_bits_stateVec_rfile[29][24]),
    .dbg_bits_stateVec_29_rfile_25     (dbg_bits_stateVec_rfile[29][25]),
    .dbg_bits_stateVec_29_rfile_26     (dbg_bits_stateVec_rfile[29][26]),
    .dbg_bits_stateVec_29_rfile_27     (dbg_bits_stateVec_rfile[29][27]),
    .dbg_bits_stateVec_29_rfile_28     (dbg_bits_stateVec_rfile[29][28]),
    .dbg_bits_stateVec_29_rfile_29     (dbg_bits_stateVec_rfile[29][29]),
    .dbg_bits_stateVec_29_rfile_30     (dbg_bits_stateVec_rfile[29][30]),
    .dbg_bits_stateVec_29_rfile_31     (dbg_bits_stateVec_rfile[29][31]),
    .dbg_bits_stateVec_29_regs_PC      (dbg_bits_stateVec_regs_PC  [29]),
    .dbg_bits_stateVec_29_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[29]),
    .dbg_bits_stateVec_30_rfile_0      (dbg_bits_stateVec_rfile[30][0 ]),
    .dbg_bits_stateVec_30_rfile_1      (dbg_bits_stateVec_rfile[30][1 ]),
    .dbg_bits_stateVec_30_rfile_2      (dbg_bits_stateVec_rfile[30][2 ]),
    .dbg_bits_stateVec_30_rfile_3      (dbg_bits_stateVec_rfile[30][3 ]),
    .dbg_bits_stateVec_30_rfile_4      (dbg_bits_stateVec_rfile[30][4 ]),
    .dbg_bits_stateVec_30_rfile_5      (dbg_bits_stateVec_rfile[30][5 ]),
    .dbg_bits_stateVec_30_rfile_6      (dbg_bits_stateVec_rfile[30][6 ]),
    .dbg_bits_stateVec_30_rfile_7      (dbg_bits_stateVec_rfile[30][7 ]),
    .dbg_bits_stateVec_30_rfile_8      (dbg_bits_stateVec_rfile[30][8 ]),
    .dbg_bits_stateVec_30_rfile_9      (dbg_bits_stateVec_rfile[30][9 ]),
    .dbg_bits_stateVec_30_rfile_10     (dbg_bits_stateVec_rfile[30][10]),
    .dbg_bits_stateVec_30_rfile_11     (dbg_bits_stateVec_rfile[30][11]),
    .dbg_bits_stateVec_30_rfile_12     (dbg_bits_stateVec_rfile[30][12]),
    .dbg_bits_stateVec_30_rfile_13     (dbg_bits_stateVec_rfile[30][13]),
    .dbg_bits_stateVec_30_rfile_14     (dbg_bits_stateVec_rfile[30][14]),
    .dbg_bits_stateVec_30_rfile_15     (dbg_bits_stateVec_rfile[30][15]),
    .dbg_bits_stateVec_30_rfile_16     (dbg_bits_stateVec_rfile[30][16]),
    .dbg_bits_stateVec_30_rfile_17     (dbg_bits_stateVec_rfile[30][17]),
    .dbg_bits_stateVec_30_rfile_18     (dbg_bits_stateVec_rfile[30][18]),
    .dbg_bits_stateVec_30_rfile_19     (dbg_bits_stateVec_rfile[30][19]),
    .dbg_bits_stateVec_30_rfile_20     (dbg_bits_stateVec_rfile[30][20]),
    .dbg_bits_stateVec_30_rfile_21     (dbg_bits_stateVec_rfile[30][21]),
    .dbg_bits_stateVec_30_rfile_22     (dbg_bits_stateVec_rfile[30][22]),
    .dbg_bits_stateVec_30_rfile_23     (dbg_bits_stateVec_rfile[30][23]),
    .dbg_bits_stateVec_30_rfile_24     (dbg_bits_stateVec_rfile[30][24]),
    .dbg_bits_stateVec_30_rfile_25     (dbg_bits_stateVec_rfile[30][25]),
    .dbg_bits_stateVec_30_rfile_26     (dbg_bits_stateVec_rfile[30][26]),
    .dbg_bits_stateVec_30_rfile_27     (dbg_bits_stateVec_rfile[30][27]),
    .dbg_bits_stateVec_30_rfile_28     (dbg_bits_stateVec_rfile[30][28]),
    .dbg_bits_stateVec_30_rfile_29     (dbg_bits_stateVec_rfile[30][29]),
    .dbg_bits_stateVec_30_rfile_30     (dbg_bits_stateVec_rfile[30][30]),
    .dbg_bits_stateVec_30_rfile_31     (dbg_bits_stateVec_rfile[30][31]),
    .dbg_bits_stateVec_30_regs_PC      (dbg_bits_stateVec_regs_PC  [30]),
    .dbg_bits_stateVec_30_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[30]),
    .dbg_bits_stateVec_31_rfile_0      (dbg_bits_stateVec_rfile[31][0 ]),
    .dbg_bits_stateVec_31_rfile_1      (dbg_bits_stateVec_rfile[31][1 ]),
    .dbg_bits_stateVec_31_rfile_2      (dbg_bits_stateVec_rfile[31][2 ]),
    .dbg_bits_stateVec_31_rfile_3      (dbg_bits_stateVec_rfile[31][3 ]),
    .dbg_bits_stateVec_31_rfile_4      (dbg_bits_stateVec_rfile[31][4 ]),
    .dbg_bits_stateVec_31_rfile_5      (dbg_bits_stateVec_rfile[31][5 ]),
    .dbg_bits_stateVec_31_rfile_6      (dbg_bits_stateVec_rfile[31][6 ]),
    .dbg_bits_stateVec_31_rfile_7      (dbg_bits_stateVec_rfile[31][7 ]),
    .dbg_bits_stateVec_31_rfile_8      (dbg_bits_stateVec_rfile[31][8 ]),
    .dbg_bits_stateVec_31_rfile_9      (dbg_bits_stateVec_rfile[31][9 ]),
    .dbg_bits_stateVec_31_rfile_10     (dbg_bits_stateVec_rfile[31][10]),
    .dbg_bits_stateVec_31_rfile_11     (dbg_bits_stateVec_rfile[31][11]),
    .dbg_bits_stateVec_31_rfile_12     (dbg_bits_stateVec_rfile[31][12]),
    .dbg_bits_stateVec_31_rfile_13     (dbg_bits_stateVec_rfile[31][13]),
    .dbg_bits_stateVec_31_rfile_14     (dbg_bits_stateVec_rfile[31][14]),
    .dbg_bits_stateVec_31_rfile_15     (dbg_bits_stateVec_rfile[31][15]),
    .dbg_bits_stateVec_31_rfile_16     (dbg_bits_stateVec_rfile[31][16]),
    .dbg_bits_stateVec_31_rfile_17     (dbg_bits_stateVec_rfile[31][17]),
    .dbg_bits_stateVec_31_rfile_18     (dbg_bits_stateVec_rfile[31][18]),
    .dbg_bits_stateVec_31_rfile_19     (dbg_bits_stateVec_rfile[31][19]),
    .dbg_bits_stateVec_31_rfile_20     (dbg_bits_stateVec_rfile[31][20]),
    .dbg_bits_stateVec_31_rfile_21     (dbg_bits_stateVec_rfile[31][21]),
    .dbg_bits_stateVec_31_rfile_22     (dbg_bits_stateVec_rfile[31][22]),
    .dbg_bits_stateVec_31_rfile_23     (dbg_bits_stateVec_rfile[31][23]),
    .dbg_bits_stateVec_31_rfile_24     (dbg_bits_stateVec_rfile[31][24]),
    .dbg_bits_stateVec_31_rfile_25     (dbg_bits_stateVec_rfile[31][25]),
    .dbg_bits_stateVec_31_rfile_26     (dbg_bits_stateVec_rfile[31][26]),
    .dbg_bits_stateVec_31_rfile_27     (dbg_bits_stateVec_rfile[31][27]),
    .dbg_bits_stateVec_31_rfile_28     (dbg_bits_stateVec_rfile[31][28]),
    .dbg_bits_stateVec_31_rfile_29     (dbg_bits_stateVec_rfile[31][29]),
    .dbg_bits_stateVec_31_rfile_30     (dbg_bits_stateVec_rfile[31][30]),
    .dbg_bits_stateVec_31_rfile_31     (dbg_bits_stateVec_rfile[31][31]),
    .dbg_bits_stateVec_31_regs_PC      (dbg_bits_stateVec_regs_PC  [31]),
    .dbg_bits_stateVec_31_regs_NZCV    (dbg_bits_stateVec_regs_NZCV[31])
`endif
    );
endmodule
