module ShiftALU( // @[:@1711.2]
  input  [63:0] io_word, // @[:@1714.4]
  input  [5:0]  io_amount, // @[:@1714.4]
  input  [1:0]  io_opcode, // @[:@1714.4]
  output [63:0] io_res // @[:@1714.4]
);
  wire [126:0] _GEN_8192; // @[execute.scala 86:33:@1716.4]
  wire [126:0] _T_15; // @[execute.scala 86:33:@1716.4]
  wire [63:0] _T_16; // @[execute.scala 87:33:@1717.4]
  wire [63:0] _T_17; // @[execute.scala 88:39:@1718.4]
  wire [63:0] _T_18; // @[execute.scala 88:42:@1719.4]
  wire [63:0] _T_19; // @[execute.scala 88:62:@1720.4]
  wire  _T_20; // @[execute.scala 89:52:@1721.4]
  wire  _T_21; // @[execute.scala 89:52:@1722.4]
  wire  _T_22; // @[execute.scala 89:52:@1723.4]
  wire  _T_23; // @[execute.scala 89:52:@1724.4]
  wire  _T_24; // @[execute.scala 89:52:@1725.4]
  wire  _T_25; // @[execute.scala 89:52:@1726.4]
  wire  _T_26; // @[execute.scala 89:52:@1727.4]
  wire  _T_27; // @[execute.scala 89:52:@1728.4]
  wire  _T_28; // @[execute.scala 89:52:@1729.4]
  wire  _T_29; // @[execute.scala 89:52:@1730.4]
  wire  _T_30; // @[execute.scala 89:52:@1731.4]
  wire  _T_31; // @[execute.scala 89:52:@1732.4]
  wire  _T_32; // @[execute.scala 89:52:@1733.4]
  wire  _T_33; // @[execute.scala 89:52:@1734.4]
  wire  _T_34; // @[execute.scala 89:52:@1735.4]
  wire  _T_35; // @[execute.scala 89:52:@1736.4]
  wire  _T_36; // @[execute.scala 89:52:@1737.4]
  wire  _T_37; // @[execute.scala 89:52:@1738.4]
  wire  _T_38; // @[execute.scala 89:52:@1739.4]
  wire  _T_39; // @[execute.scala 89:52:@1740.4]
  wire  _T_40; // @[execute.scala 89:52:@1741.4]
  wire  _T_41; // @[execute.scala 89:52:@1742.4]
  wire  _T_42; // @[execute.scala 89:52:@1743.4]
  wire  _T_43; // @[execute.scala 89:52:@1744.4]
  wire  _T_44; // @[execute.scala 89:52:@1745.4]
  wire  _T_45; // @[execute.scala 89:52:@1746.4]
  wire  _T_46; // @[execute.scala 89:52:@1747.4]
  wire  _T_47; // @[execute.scala 89:52:@1748.4]
  wire  _T_48; // @[execute.scala 89:52:@1749.4]
  wire  _T_49; // @[execute.scala 89:52:@1750.4]
  wire  _T_50; // @[execute.scala 89:52:@1751.4]
  wire  _T_51; // @[execute.scala 89:52:@1752.4]
  wire  _T_52; // @[execute.scala 89:52:@1753.4]
  wire  _T_53; // @[execute.scala 89:52:@1754.4]
  wire  _T_54; // @[execute.scala 89:52:@1755.4]
  wire  _T_55; // @[execute.scala 89:52:@1756.4]
  wire  _T_56; // @[execute.scala 89:52:@1757.4]
  wire  _T_57; // @[execute.scala 89:52:@1758.4]
  wire  _T_58; // @[execute.scala 89:52:@1759.4]
  wire  _T_59; // @[execute.scala 89:52:@1760.4]
  wire  _T_60; // @[execute.scala 89:52:@1761.4]
  wire  _T_61; // @[execute.scala 89:52:@1762.4]
  wire  _T_62; // @[execute.scala 89:52:@1763.4]
  wire  _T_63; // @[execute.scala 89:52:@1764.4]
  wire  _T_64; // @[execute.scala 89:52:@1765.4]
  wire  _T_65; // @[execute.scala 89:52:@1766.4]
  wire  _T_66; // @[execute.scala 89:52:@1767.4]
  wire  _T_67; // @[execute.scala 89:52:@1768.4]
  wire  _T_68; // @[execute.scala 89:52:@1769.4]
  wire  _T_69; // @[execute.scala 89:52:@1770.4]
  wire  _T_70; // @[execute.scala 89:52:@1771.4]
  wire  _T_71; // @[execute.scala 89:52:@1772.4]
  wire  _T_72; // @[execute.scala 89:52:@1773.4]
  wire  _T_73; // @[execute.scala 89:52:@1774.4]
  wire  _T_74; // @[execute.scala 89:52:@1775.4]
  wire  _T_75; // @[execute.scala 89:52:@1776.4]
  wire  _T_76; // @[execute.scala 89:52:@1777.4]
  wire  _T_77; // @[execute.scala 89:52:@1778.4]
  wire  _T_78; // @[execute.scala 89:52:@1779.4]
  wire  _T_79; // @[execute.scala 89:52:@1780.4]
  wire  _T_80; // @[execute.scala 89:52:@1781.4]
  wire  _T_81; // @[execute.scala 89:52:@1782.4]
  wire  _T_82; // @[execute.scala 89:52:@1783.4]
  wire  _T_83; // @[execute.scala 89:52:@1784.4]
  wire [6:0] _GEN_8193; // @[execute.scala 79:37:@1851.4]
  wire [7:0] _T_157; // @[execute.scala 79:37:@1851.4]
  wire [7:0] _T_158; // @[execute.scala 79:37:@1852.4]
  wire [6:0] _T_159; // @[execute.scala 79:37:@1853.4]
  wire [5:0] _T_161; // @[:@1854.4]
  wire  _GEN_1; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_2; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_3; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_4; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_5; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_6; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_7; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_8; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_9; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_10; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_11; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_12; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_13; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_14; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_15; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_16; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_17; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_18; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_19; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_20; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_21; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_22; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_23; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_24; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_25; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_26; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_27; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_28; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_29; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_30; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_31; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_32; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_33; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_34; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_35; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_36; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_37; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_38; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_39; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_40; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_41; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_42; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_43; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_44; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_45; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_46; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_47; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_48; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_49; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_50; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_51; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_52; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_53; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_54; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_55; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_56; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_57; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_58; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_59; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_60; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_61; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_62; // @[execute.scala 79:10:@1857.4]
  wire  _GEN_63; // @[execute.scala 79:10:@1857.4]
  wire  _T_168; // @[execute.scala 79:15:@1858.4]
  wire [6:0] _T_170; // @[execute.scala 79:37:@1859.4]
  wire [6:0] _T_171; // @[execute.scala 79:37:@1860.4]
  wire [5:0] _T_172; // @[execute.scala 79:37:@1861.4]
  wire [6:0] _T_175; // @[execute.scala 79:60:@1862.4]
  wire [5:0] _T_176; // @[execute.scala 79:60:@1863.4]
  wire  _GEN_129; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_130; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_131; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_132; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_133; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_134; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_135; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_136; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_137; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_138; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_139; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_140; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_141; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_142; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_143; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_144; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_145; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_146; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_147; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_148; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_149; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_150; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_151; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_152; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_153; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_154; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_155; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_156; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_157; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_158; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_159; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_160; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_161; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_162; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_163; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_164; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_165; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_166; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_167; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_168; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_169; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_170; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_171; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_172; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_173; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_174; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_175; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_176; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_177; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_178; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_179; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_180; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_181; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_182; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_183; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_184; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_185; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_186; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_187; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_188; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_189; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_190; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_191; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_193; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_194; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_195; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_196; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_197; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_198; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_199; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_200; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_201; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_202; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_203; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_204; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_205; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_206; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_207; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_208; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_209; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_210; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_211; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_212; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_213; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_214; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_215; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_216; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_217; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_218; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_219; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_220; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_221; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_222; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_223; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_224; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_225; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_226; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_227; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_228; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_229; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_230; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_231; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_232; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_233; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_234; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_235; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_236; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_237; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_238; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_239; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_240; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_241; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_242; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_243; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_244; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_245; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_246; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_247; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_248; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_249; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_250; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_251; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_252; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_253; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_254; // @[execute.scala 79:10:@1864.4]
  wire  _GEN_255; // @[execute.scala 79:10:@1864.4]
  wire  _T_178; // @[execute.scala 79:10:@1864.4]
  wire  _T_180; // @[execute.scala 79:15:@1865.4]
  wire [6:0] _T_182; // @[execute.scala 79:37:@1866.4]
  wire [6:0] _T_183; // @[execute.scala 79:37:@1867.4]
  wire [5:0] _T_184; // @[execute.scala 79:37:@1868.4]
  wire [6:0] _T_187; // @[execute.scala 79:60:@1869.4]
  wire [5:0] _T_188; // @[execute.scala 79:60:@1870.4]
  wire  _GEN_257; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_258; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_259; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_260; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_261; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_262; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_263; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_264; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_265; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_266; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_267; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_268; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_269; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_270; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_271; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_272; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_273; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_274; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_275; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_276; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_277; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_278; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_279; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_280; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_281; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_282; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_283; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_284; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_285; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_286; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_287; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_288; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_289; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_290; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_291; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_292; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_293; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_294; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_295; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_296; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_297; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_298; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_299; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_300; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_301; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_302; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_303; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_304; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_305; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_306; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_307; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_308; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_309; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_310; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_311; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_312; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_313; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_314; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_315; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_316; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_317; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_318; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_319; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_321; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_322; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_323; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_324; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_325; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_326; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_327; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_328; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_329; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_330; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_331; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_332; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_333; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_334; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_335; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_336; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_337; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_338; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_339; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_340; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_341; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_342; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_343; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_344; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_345; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_346; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_347; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_348; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_349; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_350; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_351; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_352; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_353; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_354; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_355; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_356; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_357; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_358; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_359; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_360; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_361; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_362; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_363; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_364; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_365; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_366; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_367; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_368; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_369; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_370; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_371; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_372; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_373; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_374; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_375; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_376; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_377; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_378; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_379; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_380; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_381; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_382; // @[execute.scala 79:10:@1871.4]
  wire  _GEN_383; // @[execute.scala 79:10:@1871.4]
  wire  _T_190; // @[execute.scala 79:10:@1871.4]
  wire  _T_192; // @[execute.scala 79:15:@1872.4]
  wire [6:0] _T_194; // @[execute.scala 79:37:@1873.4]
  wire [6:0] _T_195; // @[execute.scala 79:37:@1874.4]
  wire [5:0] _T_196; // @[execute.scala 79:37:@1875.4]
  wire [6:0] _T_199; // @[execute.scala 79:60:@1876.4]
  wire [5:0] _T_200; // @[execute.scala 79:60:@1877.4]
  wire  _GEN_385; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_386; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_387; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_388; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_389; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_390; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_391; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_392; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_393; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_394; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_395; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_396; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_397; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_398; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_399; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_400; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_401; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_402; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_403; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_404; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_405; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_406; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_407; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_408; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_409; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_410; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_411; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_412; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_413; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_414; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_415; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_416; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_417; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_418; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_419; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_420; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_421; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_422; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_423; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_424; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_425; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_426; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_427; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_428; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_429; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_430; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_431; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_432; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_433; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_434; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_435; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_436; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_437; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_438; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_439; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_440; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_441; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_442; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_443; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_444; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_445; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_446; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_447; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_449; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_450; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_451; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_452; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_453; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_454; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_455; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_456; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_457; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_458; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_459; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_460; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_461; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_462; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_463; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_464; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_465; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_466; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_467; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_468; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_469; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_470; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_471; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_472; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_473; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_474; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_475; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_476; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_477; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_478; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_479; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_480; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_481; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_482; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_483; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_484; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_485; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_486; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_487; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_488; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_489; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_490; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_491; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_492; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_493; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_494; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_495; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_496; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_497; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_498; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_499; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_500; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_501; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_502; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_503; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_504; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_505; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_506; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_507; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_508; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_509; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_510; // @[execute.scala 79:10:@1878.4]
  wire  _GEN_511; // @[execute.scala 79:10:@1878.4]
  wire  _T_202; // @[execute.scala 79:10:@1878.4]
  wire  _T_204; // @[execute.scala 79:15:@1879.4]
  wire [6:0] _T_206; // @[execute.scala 79:37:@1880.4]
  wire [6:0] _T_207; // @[execute.scala 79:37:@1881.4]
  wire [5:0] _T_208; // @[execute.scala 79:37:@1882.4]
  wire [6:0] _T_211; // @[execute.scala 79:60:@1883.4]
  wire [5:0] _T_212; // @[execute.scala 79:60:@1884.4]
  wire  _GEN_513; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_514; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_515; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_516; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_517; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_518; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_519; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_520; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_521; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_522; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_523; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_524; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_525; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_526; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_527; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_528; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_529; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_530; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_531; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_532; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_533; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_534; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_535; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_536; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_537; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_538; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_539; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_540; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_541; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_542; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_543; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_544; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_545; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_546; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_547; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_548; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_549; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_550; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_551; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_552; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_553; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_554; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_555; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_556; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_557; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_558; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_559; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_560; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_561; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_562; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_563; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_564; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_565; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_566; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_567; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_568; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_569; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_570; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_571; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_572; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_573; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_574; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_575; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_577; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_578; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_579; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_580; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_581; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_582; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_583; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_584; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_585; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_586; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_587; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_588; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_589; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_590; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_591; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_592; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_593; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_594; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_595; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_596; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_597; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_598; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_599; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_600; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_601; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_602; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_603; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_604; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_605; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_606; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_607; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_608; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_609; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_610; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_611; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_612; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_613; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_614; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_615; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_616; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_617; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_618; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_619; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_620; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_621; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_622; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_623; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_624; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_625; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_626; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_627; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_628; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_629; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_630; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_631; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_632; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_633; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_634; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_635; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_636; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_637; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_638; // @[execute.scala 79:10:@1885.4]
  wire  _GEN_639; // @[execute.scala 79:10:@1885.4]
  wire  _T_214; // @[execute.scala 79:10:@1885.4]
  wire  _T_216; // @[execute.scala 79:15:@1886.4]
  wire [6:0] _T_218; // @[execute.scala 79:37:@1887.4]
  wire [6:0] _T_219; // @[execute.scala 79:37:@1888.4]
  wire [5:0] _T_220; // @[execute.scala 79:37:@1889.4]
  wire [6:0] _T_223; // @[execute.scala 79:60:@1890.4]
  wire [5:0] _T_224; // @[execute.scala 79:60:@1891.4]
  wire  _GEN_641; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_642; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_643; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_644; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_645; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_646; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_647; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_648; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_649; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_650; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_651; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_652; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_653; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_654; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_655; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_656; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_657; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_658; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_659; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_660; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_661; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_662; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_663; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_664; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_665; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_666; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_667; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_668; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_669; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_670; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_671; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_672; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_673; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_674; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_675; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_676; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_677; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_678; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_679; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_680; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_681; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_682; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_683; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_684; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_685; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_686; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_687; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_688; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_689; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_690; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_691; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_692; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_693; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_694; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_695; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_696; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_697; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_698; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_699; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_700; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_701; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_702; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_703; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_705; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_706; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_707; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_708; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_709; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_710; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_711; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_712; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_713; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_714; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_715; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_716; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_717; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_718; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_719; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_720; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_721; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_722; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_723; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_724; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_725; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_726; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_727; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_728; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_729; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_730; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_731; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_732; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_733; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_734; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_735; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_736; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_737; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_738; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_739; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_740; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_741; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_742; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_743; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_744; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_745; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_746; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_747; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_748; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_749; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_750; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_751; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_752; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_753; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_754; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_755; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_756; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_757; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_758; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_759; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_760; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_761; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_762; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_763; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_764; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_765; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_766; // @[execute.scala 79:10:@1892.4]
  wire  _GEN_767; // @[execute.scala 79:10:@1892.4]
  wire  _T_226; // @[execute.scala 79:10:@1892.4]
  wire  _T_228; // @[execute.scala 79:15:@1893.4]
  wire [6:0] _T_230; // @[execute.scala 79:37:@1894.4]
  wire [6:0] _T_231; // @[execute.scala 79:37:@1895.4]
  wire [5:0] _T_232; // @[execute.scala 79:37:@1896.4]
  wire [6:0] _T_235; // @[execute.scala 79:60:@1897.4]
  wire [5:0] _T_236; // @[execute.scala 79:60:@1898.4]
  wire  _GEN_769; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_770; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_771; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_772; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_773; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_774; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_775; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_776; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_777; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_778; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_779; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_780; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_781; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_782; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_783; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_784; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_785; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_786; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_787; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_788; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_789; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_790; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_791; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_792; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_793; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_794; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_795; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_796; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_797; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_798; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_799; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_800; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_801; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_802; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_803; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_804; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_805; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_806; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_807; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_808; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_809; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_810; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_811; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_812; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_813; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_814; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_815; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_816; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_817; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_818; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_819; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_820; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_821; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_822; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_823; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_824; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_825; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_826; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_827; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_828; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_829; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_830; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_831; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_833; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_834; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_835; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_836; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_837; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_838; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_839; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_840; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_841; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_842; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_843; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_844; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_845; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_846; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_847; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_848; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_849; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_850; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_851; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_852; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_853; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_854; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_855; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_856; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_857; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_858; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_859; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_860; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_861; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_862; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_863; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_864; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_865; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_866; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_867; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_868; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_869; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_870; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_871; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_872; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_873; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_874; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_875; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_876; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_877; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_878; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_879; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_880; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_881; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_882; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_883; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_884; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_885; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_886; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_887; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_888; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_889; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_890; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_891; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_892; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_893; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_894; // @[execute.scala 79:10:@1899.4]
  wire  _GEN_895; // @[execute.scala 79:10:@1899.4]
  wire  _T_238; // @[execute.scala 79:10:@1899.4]
  wire  _T_240; // @[execute.scala 79:15:@1900.4]
  wire [6:0] _T_242; // @[execute.scala 79:37:@1901.4]
  wire [6:0] _T_243; // @[execute.scala 79:37:@1902.4]
  wire [5:0] _T_244; // @[execute.scala 79:37:@1903.4]
  wire [6:0] _T_247; // @[execute.scala 79:60:@1904.4]
  wire [5:0] _T_248; // @[execute.scala 79:60:@1905.4]
  wire  _GEN_897; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_898; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_899; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_900; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_901; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_902; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_903; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_904; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_905; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_906; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_907; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_908; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_909; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_910; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_911; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_912; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_913; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_914; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_915; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_916; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_917; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_918; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_919; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_920; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_921; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_922; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_923; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_924; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_925; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_926; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_927; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_928; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_929; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_930; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_931; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_932; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_933; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_934; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_935; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_936; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_937; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_938; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_939; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_940; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_941; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_942; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_943; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_944; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_945; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_946; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_947; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_948; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_949; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_950; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_951; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_952; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_953; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_954; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_955; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_956; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_957; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_958; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_959; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_961; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_962; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_963; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_964; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_965; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_966; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_967; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_968; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_969; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_970; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_971; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_972; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_973; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_974; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_975; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_976; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_977; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_978; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_979; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_980; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_981; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_982; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_983; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_984; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_985; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_986; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_987; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_988; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_989; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_990; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_991; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_992; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_993; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_994; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_995; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_996; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_997; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_998; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_999; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1000; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1001; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1002; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1003; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1004; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1005; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1006; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1007; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1008; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1009; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1010; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1011; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1012; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1013; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1014; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1015; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1016; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1017; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1018; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1019; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1020; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1021; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1022; // @[execute.scala 79:10:@1906.4]
  wire  _GEN_1023; // @[execute.scala 79:10:@1906.4]
  wire  _T_250; // @[execute.scala 79:10:@1906.4]
  wire  _T_252; // @[execute.scala 79:15:@1907.4]
  wire [6:0] _T_254; // @[execute.scala 79:37:@1908.4]
  wire [6:0] _T_255; // @[execute.scala 79:37:@1909.4]
  wire [5:0] _T_256; // @[execute.scala 79:37:@1910.4]
  wire [6:0] _T_259; // @[execute.scala 79:60:@1911.4]
  wire [5:0] _T_260; // @[execute.scala 79:60:@1912.4]
  wire  _GEN_1025; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1026; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1027; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1028; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1029; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1030; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1031; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1032; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1033; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1034; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1035; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1036; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1037; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1038; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1039; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1040; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1041; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1042; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1043; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1044; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1045; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1046; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1047; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1048; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1049; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1050; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1051; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1052; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1053; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1054; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1055; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1056; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1057; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1058; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1059; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1060; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1061; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1062; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1063; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1064; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1065; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1066; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1067; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1068; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1069; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1070; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1071; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1072; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1073; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1074; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1075; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1076; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1077; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1078; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1079; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1080; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1081; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1082; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1083; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1084; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1085; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1086; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1087; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1089; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1090; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1091; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1092; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1093; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1094; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1095; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1096; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1097; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1098; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1099; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1100; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1101; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1102; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1103; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1104; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1105; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1106; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1107; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1108; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1109; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1110; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1111; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1112; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1113; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1114; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1115; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1116; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1117; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1118; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1119; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1120; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1121; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1122; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1123; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1124; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1125; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1126; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1127; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1128; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1129; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1130; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1131; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1132; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1133; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1134; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1135; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1136; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1137; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1138; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1139; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1140; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1141; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1142; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1143; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1144; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1145; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1146; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1147; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1148; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1149; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1150; // @[execute.scala 79:10:@1913.4]
  wire  _GEN_1151; // @[execute.scala 79:10:@1913.4]
  wire  _T_262; // @[execute.scala 79:10:@1913.4]
  wire  _T_264; // @[execute.scala 79:15:@1914.4]
  wire [6:0] _T_266; // @[execute.scala 79:37:@1915.4]
  wire [6:0] _T_267; // @[execute.scala 79:37:@1916.4]
  wire [5:0] _T_268; // @[execute.scala 79:37:@1917.4]
  wire [6:0] _T_271; // @[execute.scala 79:60:@1918.4]
  wire [5:0] _T_272; // @[execute.scala 79:60:@1919.4]
  wire  _GEN_1153; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1154; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1155; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1156; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1157; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1158; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1159; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1160; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1161; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1162; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1163; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1164; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1165; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1166; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1167; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1168; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1169; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1170; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1171; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1172; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1173; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1174; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1175; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1176; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1177; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1178; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1179; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1180; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1181; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1182; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1183; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1184; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1185; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1186; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1187; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1188; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1189; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1190; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1191; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1192; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1193; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1194; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1195; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1196; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1197; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1198; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1199; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1200; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1201; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1202; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1203; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1204; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1205; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1206; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1207; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1208; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1209; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1210; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1211; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1212; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1213; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1214; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1215; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1217; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1218; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1219; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1220; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1221; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1222; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1223; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1224; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1225; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1226; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1227; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1228; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1229; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1230; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1231; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1232; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1233; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1234; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1235; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1236; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1237; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1238; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1239; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1240; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1241; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1242; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1243; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1244; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1245; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1246; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1247; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1248; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1249; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1250; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1251; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1252; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1253; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1254; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1255; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1256; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1257; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1258; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1259; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1260; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1261; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1262; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1263; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1264; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1265; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1266; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1267; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1268; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1269; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1270; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1271; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1272; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1273; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1274; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1275; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1276; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1277; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1278; // @[execute.scala 79:10:@1920.4]
  wire  _GEN_1279; // @[execute.scala 79:10:@1920.4]
  wire  _T_274; // @[execute.scala 79:10:@1920.4]
  wire  _T_276; // @[execute.scala 79:15:@1921.4]
  wire [6:0] _T_278; // @[execute.scala 79:37:@1922.4]
  wire [6:0] _T_279; // @[execute.scala 79:37:@1923.4]
  wire [5:0] _T_280; // @[execute.scala 79:37:@1924.4]
  wire [6:0] _T_283; // @[execute.scala 79:60:@1925.4]
  wire [5:0] _T_284; // @[execute.scala 79:60:@1926.4]
  wire  _GEN_1281; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1282; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1283; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1284; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1285; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1286; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1287; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1288; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1289; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1290; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1291; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1292; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1293; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1294; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1295; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1296; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1297; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1298; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1299; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1300; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1301; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1302; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1303; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1304; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1305; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1306; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1307; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1308; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1309; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1310; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1311; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1312; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1313; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1314; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1315; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1316; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1317; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1318; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1319; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1320; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1321; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1322; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1323; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1324; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1325; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1326; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1327; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1328; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1329; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1330; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1331; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1332; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1333; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1334; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1335; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1336; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1337; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1338; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1339; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1340; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1341; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1342; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1343; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1345; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1346; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1347; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1348; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1349; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1350; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1351; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1352; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1353; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1354; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1355; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1356; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1357; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1358; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1359; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1360; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1361; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1362; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1363; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1364; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1365; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1366; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1367; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1368; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1369; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1370; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1371; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1372; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1373; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1374; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1375; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1376; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1377; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1378; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1379; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1380; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1381; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1382; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1383; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1384; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1385; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1386; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1387; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1388; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1389; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1390; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1391; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1392; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1393; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1394; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1395; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1396; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1397; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1398; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1399; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1400; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1401; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1402; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1403; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1404; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1405; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1406; // @[execute.scala 79:10:@1927.4]
  wire  _GEN_1407; // @[execute.scala 79:10:@1927.4]
  wire  _T_286; // @[execute.scala 79:10:@1927.4]
  wire  _T_288; // @[execute.scala 79:15:@1928.4]
  wire [6:0] _T_290; // @[execute.scala 79:37:@1929.4]
  wire [6:0] _T_291; // @[execute.scala 79:37:@1930.4]
  wire [5:0] _T_292; // @[execute.scala 79:37:@1931.4]
  wire [6:0] _T_295; // @[execute.scala 79:60:@1932.4]
  wire [5:0] _T_296; // @[execute.scala 79:60:@1933.4]
  wire  _GEN_1409; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1410; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1411; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1412; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1413; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1414; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1415; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1416; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1417; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1418; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1419; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1420; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1421; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1422; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1423; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1424; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1425; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1426; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1427; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1428; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1429; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1430; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1431; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1432; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1433; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1434; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1435; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1436; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1437; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1438; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1439; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1440; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1441; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1442; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1443; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1444; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1445; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1446; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1447; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1448; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1449; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1450; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1451; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1452; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1453; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1454; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1455; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1456; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1457; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1458; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1459; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1460; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1461; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1462; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1463; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1464; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1465; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1466; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1467; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1468; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1469; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1470; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1471; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1473; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1474; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1475; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1476; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1477; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1478; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1479; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1480; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1481; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1482; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1483; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1484; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1485; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1486; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1487; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1488; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1489; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1490; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1491; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1492; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1493; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1494; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1495; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1496; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1497; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1498; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1499; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1500; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1501; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1502; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1503; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1504; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1505; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1506; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1507; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1508; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1509; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1510; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1511; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1512; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1513; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1514; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1515; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1516; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1517; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1518; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1519; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1520; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1521; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1522; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1523; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1524; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1525; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1526; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1527; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1528; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1529; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1530; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1531; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1532; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1533; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1534; // @[execute.scala 79:10:@1934.4]
  wire  _GEN_1535; // @[execute.scala 79:10:@1934.4]
  wire  _T_298; // @[execute.scala 79:10:@1934.4]
  wire  _T_300; // @[execute.scala 79:15:@1935.4]
  wire [6:0] _T_302; // @[execute.scala 79:37:@1936.4]
  wire [6:0] _T_303; // @[execute.scala 79:37:@1937.4]
  wire [5:0] _T_304; // @[execute.scala 79:37:@1938.4]
  wire [6:0] _T_307; // @[execute.scala 79:60:@1939.4]
  wire [5:0] _T_308; // @[execute.scala 79:60:@1940.4]
  wire  _GEN_1537; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1538; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1539; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1540; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1541; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1542; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1543; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1544; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1545; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1546; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1547; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1548; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1549; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1550; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1551; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1552; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1553; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1554; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1555; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1556; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1557; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1558; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1559; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1560; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1561; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1562; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1563; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1564; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1565; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1566; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1567; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1568; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1569; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1570; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1571; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1572; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1573; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1574; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1575; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1576; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1577; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1578; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1579; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1580; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1581; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1582; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1583; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1584; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1585; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1586; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1587; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1588; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1589; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1590; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1591; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1592; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1593; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1594; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1595; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1596; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1597; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1598; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1599; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1601; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1602; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1603; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1604; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1605; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1606; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1607; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1608; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1609; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1610; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1611; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1612; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1613; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1614; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1615; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1616; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1617; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1618; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1619; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1620; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1621; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1622; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1623; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1624; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1625; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1626; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1627; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1628; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1629; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1630; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1631; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1632; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1633; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1634; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1635; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1636; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1637; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1638; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1639; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1640; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1641; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1642; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1643; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1644; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1645; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1646; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1647; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1648; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1649; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1650; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1651; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1652; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1653; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1654; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1655; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1656; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1657; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1658; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1659; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1660; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1661; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1662; // @[execute.scala 79:10:@1941.4]
  wire  _GEN_1663; // @[execute.scala 79:10:@1941.4]
  wire  _T_310; // @[execute.scala 79:10:@1941.4]
  wire  _T_312; // @[execute.scala 79:15:@1942.4]
  wire [6:0] _T_314; // @[execute.scala 79:37:@1943.4]
  wire [6:0] _T_315; // @[execute.scala 79:37:@1944.4]
  wire [5:0] _T_316; // @[execute.scala 79:37:@1945.4]
  wire [6:0] _T_319; // @[execute.scala 79:60:@1946.4]
  wire [5:0] _T_320; // @[execute.scala 79:60:@1947.4]
  wire  _GEN_1665; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1666; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1667; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1668; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1669; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1670; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1671; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1672; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1673; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1674; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1675; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1676; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1677; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1678; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1679; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1680; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1681; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1682; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1683; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1684; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1685; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1686; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1687; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1688; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1689; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1690; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1691; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1692; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1693; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1694; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1695; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1696; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1697; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1698; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1699; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1700; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1701; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1702; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1703; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1704; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1705; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1706; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1707; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1708; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1709; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1710; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1711; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1712; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1713; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1714; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1715; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1716; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1717; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1718; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1719; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1720; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1721; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1722; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1723; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1724; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1725; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1726; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1727; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1729; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1730; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1731; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1732; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1733; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1734; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1735; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1736; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1737; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1738; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1739; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1740; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1741; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1742; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1743; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1744; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1745; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1746; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1747; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1748; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1749; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1750; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1751; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1752; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1753; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1754; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1755; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1756; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1757; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1758; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1759; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1760; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1761; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1762; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1763; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1764; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1765; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1766; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1767; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1768; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1769; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1770; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1771; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1772; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1773; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1774; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1775; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1776; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1777; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1778; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1779; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1780; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1781; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1782; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1783; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1784; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1785; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1786; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1787; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1788; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1789; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1790; // @[execute.scala 79:10:@1948.4]
  wire  _GEN_1791; // @[execute.scala 79:10:@1948.4]
  wire  _T_322; // @[execute.scala 79:10:@1948.4]
  wire  _T_324; // @[execute.scala 79:15:@1949.4]
  wire [6:0] _T_326; // @[execute.scala 79:37:@1950.4]
  wire [6:0] _T_327; // @[execute.scala 79:37:@1951.4]
  wire [5:0] _T_328; // @[execute.scala 79:37:@1952.4]
  wire [6:0] _T_331; // @[execute.scala 79:60:@1953.4]
  wire [5:0] _T_332; // @[execute.scala 79:60:@1954.4]
  wire  _GEN_1793; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1794; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1795; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1796; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1797; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1798; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1799; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1800; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1801; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1802; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1803; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1804; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1805; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1806; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1807; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1808; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1809; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1810; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1811; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1812; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1813; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1814; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1815; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1816; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1817; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1818; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1819; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1820; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1821; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1822; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1823; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1824; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1825; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1826; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1827; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1828; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1829; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1830; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1831; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1832; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1833; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1834; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1835; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1836; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1837; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1838; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1839; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1840; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1841; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1842; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1843; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1844; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1845; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1846; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1847; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1848; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1849; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1850; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1851; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1852; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1853; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1854; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1855; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1857; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1858; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1859; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1860; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1861; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1862; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1863; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1864; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1865; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1866; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1867; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1868; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1869; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1870; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1871; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1872; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1873; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1874; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1875; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1876; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1877; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1878; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1879; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1880; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1881; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1882; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1883; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1884; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1885; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1886; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1887; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1888; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1889; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1890; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1891; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1892; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1893; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1894; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1895; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1896; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1897; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1898; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1899; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1900; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1901; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1902; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1903; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1904; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1905; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1906; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1907; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1908; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1909; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1910; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1911; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1912; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1913; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1914; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1915; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1916; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1917; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1918; // @[execute.scala 79:10:@1955.4]
  wire  _GEN_1919; // @[execute.scala 79:10:@1955.4]
  wire  _T_334; // @[execute.scala 79:10:@1955.4]
  wire  _T_336; // @[execute.scala 79:15:@1956.4]
  wire [6:0] _T_338; // @[execute.scala 79:37:@1957.4]
  wire [6:0] _T_339; // @[execute.scala 79:37:@1958.4]
  wire [5:0] _T_340; // @[execute.scala 79:37:@1959.4]
  wire [6:0] _T_343; // @[execute.scala 79:60:@1960.4]
  wire [5:0] _T_344; // @[execute.scala 79:60:@1961.4]
  wire  _GEN_1921; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1922; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1923; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1924; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1925; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1926; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1927; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1928; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1929; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1930; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1931; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1932; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1933; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1934; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1935; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1936; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1937; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1938; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1939; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1940; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1941; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1942; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1943; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1944; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1945; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1946; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1947; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1948; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1949; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1950; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1951; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1952; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1953; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1954; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1955; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1956; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1957; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1958; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1959; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1960; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1961; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1962; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1963; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1964; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1965; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1966; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1967; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1968; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1969; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1970; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1971; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1972; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1973; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1974; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1975; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1976; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1977; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1978; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1979; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1980; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1981; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1982; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1983; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1985; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1986; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1987; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1988; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1989; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1990; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1991; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1992; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1993; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1994; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1995; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1996; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1997; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1998; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_1999; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2000; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2001; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2002; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2003; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2004; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2005; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2006; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2007; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2008; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2009; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2010; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2011; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2012; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2013; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2014; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2015; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2016; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2017; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2018; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2019; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2020; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2021; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2022; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2023; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2024; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2025; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2026; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2027; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2028; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2029; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2030; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2031; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2032; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2033; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2034; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2035; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2036; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2037; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2038; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2039; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2040; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2041; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2042; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2043; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2044; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2045; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2046; // @[execute.scala 79:10:@1962.4]
  wire  _GEN_2047; // @[execute.scala 79:10:@1962.4]
  wire  _T_346; // @[execute.scala 79:10:@1962.4]
  wire  _T_348; // @[execute.scala 79:15:@1963.4]
  wire [6:0] _T_350; // @[execute.scala 79:37:@1964.4]
  wire [6:0] _T_351; // @[execute.scala 79:37:@1965.4]
  wire [5:0] _T_352; // @[execute.scala 79:37:@1966.4]
  wire [6:0] _T_355; // @[execute.scala 79:60:@1967.4]
  wire [5:0] _T_356; // @[execute.scala 79:60:@1968.4]
  wire  _GEN_2049; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2050; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2051; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2052; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2053; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2054; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2055; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2056; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2057; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2058; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2059; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2060; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2061; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2062; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2063; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2064; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2065; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2066; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2067; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2068; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2069; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2070; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2071; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2072; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2073; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2074; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2075; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2076; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2077; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2078; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2079; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2080; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2081; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2082; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2083; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2084; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2085; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2086; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2087; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2088; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2089; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2090; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2091; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2092; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2093; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2094; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2095; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2096; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2097; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2098; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2099; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2100; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2101; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2102; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2103; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2104; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2105; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2106; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2107; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2108; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2109; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2110; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2111; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2113; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2114; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2115; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2116; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2117; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2118; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2119; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2120; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2121; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2122; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2123; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2124; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2125; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2126; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2127; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2128; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2129; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2130; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2131; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2132; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2133; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2134; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2135; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2136; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2137; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2138; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2139; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2140; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2141; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2142; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2143; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2144; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2145; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2146; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2147; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2148; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2149; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2150; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2151; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2152; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2153; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2154; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2155; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2156; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2157; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2158; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2159; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2160; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2161; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2162; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2163; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2164; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2165; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2166; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2167; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2168; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2169; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2170; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2171; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2172; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2173; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2174; // @[execute.scala 79:10:@1969.4]
  wire  _GEN_2175; // @[execute.scala 79:10:@1969.4]
  wire  _T_358; // @[execute.scala 79:10:@1969.4]
  wire  _T_360; // @[execute.scala 79:15:@1970.4]
  wire [6:0] _T_362; // @[execute.scala 79:37:@1971.4]
  wire [6:0] _T_363; // @[execute.scala 79:37:@1972.4]
  wire [5:0] _T_364; // @[execute.scala 79:37:@1973.4]
  wire [6:0] _T_367; // @[execute.scala 79:60:@1974.4]
  wire [5:0] _T_368; // @[execute.scala 79:60:@1975.4]
  wire  _GEN_2177; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2178; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2179; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2180; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2181; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2182; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2183; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2184; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2185; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2186; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2187; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2188; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2189; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2190; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2191; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2192; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2193; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2194; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2195; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2196; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2197; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2198; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2199; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2200; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2201; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2202; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2203; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2204; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2205; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2206; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2207; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2208; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2209; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2210; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2211; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2212; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2213; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2214; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2215; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2216; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2217; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2218; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2219; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2220; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2221; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2222; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2223; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2224; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2225; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2226; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2227; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2228; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2229; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2230; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2231; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2232; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2233; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2234; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2235; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2236; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2237; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2238; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2239; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2241; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2242; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2243; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2244; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2245; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2246; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2247; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2248; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2249; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2250; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2251; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2252; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2253; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2254; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2255; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2256; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2257; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2258; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2259; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2260; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2261; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2262; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2263; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2264; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2265; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2266; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2267; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2268; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2269; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2270; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2271; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2272; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2273; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2274; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2275; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2276; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2277; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2278; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2279; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2280; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2281; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2282; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2283; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2284; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2285; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2286; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2287; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2288; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2289; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2290; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2291; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2292; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2293; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2294; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2295; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2296; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2297; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2298; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2299; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2300; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2301; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2302; // @[execute.scala 79:10:@1976.4]
  wire  _GEN_2303; // @[execute.scala 79:10:@1976.4]
  wire  _T_370; // @[execute.scala 79:10:@1976.4]
  wire  _T_372; // @[execute.scala 79:15:@1977.4]
  wire [6:0] _T_374; // @[execute.scala 79:37:@1978.4]
  wire [6:0] _T_375; // @[execute.scala 79:37:@1979.4]
  wire [5:0] _T_376; // @[execute.scala 79:37:@1980.4]
  wire [6:0] _T_379; // @[execute.scala 79:60:@1981.4]
  wire [5:0] _T_380; // @[execute.scala 79:60:@1982.4]
  wire  _GEN_2305; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2306; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2307; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2308; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2309; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2310; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2311; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2312; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2313; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2314; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2315; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2316; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2317; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2318; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2319; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2320; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2321; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2322; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2323; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2324; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2325; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2326; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2327; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2328; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2329; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2330; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2331; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2332; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2333; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2334; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2335; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2336; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2337; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2338; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2339; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2340; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2341; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2342; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2343; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2344; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2345; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2346; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2347; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2348; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2349; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2350; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2351; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2352; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2353; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2354; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2355; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2356; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2357; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2358; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2359; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2360; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2361; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2362; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2363; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2364; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2365; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2366; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2367; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2369; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2370; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2371; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2372; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2373; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2374; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2375; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2376; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2377; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2378; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2379; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2380; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2381; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2382; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2383; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2384; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2385; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2386; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2387; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2388; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2389; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2390; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2391; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2392; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2393; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2394; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2395; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2396; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2397; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2398; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2399; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2400; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2401; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2402; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2403; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2404; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2405; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2406; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2407; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2408; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2409; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2410; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2411; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2412; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2413; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2414; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2415; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2416; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2417; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2418; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2419; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2420; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2421; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2422; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2423; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2424; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2425; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2426; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2427; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2428; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2429; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2430; // @[execute.scala 79:10:@1983.4]
  wire  _GEN_2431; // @[execute.scala 79:10:@1983.4]
  wire  _T_382; // @[execute.scala 79:10:@1983.4]
  wire  _T_384; // @[execute.scala 79:15:@1984.4]
  wire [6:0] _T_386; // @[execute.scala 79:37:@1985.4]
  wire [6:0] _T_387; // @[execute.scala 79:37:@1986.4]
  wire [5:0] _T_388; // @[execute.scala 79:37:@1987.4]
  wire [6:0] _T_391; // @[execute.scala 79:60:@1988.4]
  wire [5:0] _T_392; // @[execute.scala 79:60:@1989.4]
  wire  _GEN_2433; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2434; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2435; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2436; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2437; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2438; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2439; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2440; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2441; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2442; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2443; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2444; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2445; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2446; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2447; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2448; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2449; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2450; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2451; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2452; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2453; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2454; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2455; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2456; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2457; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2458; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2459; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2460; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2461; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2462; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2463; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2464; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2465; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2466; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2467; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2468; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2469; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2470; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2471; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2472; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2473; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2474; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2475; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2476; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2477; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2478; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2479; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2480; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2481; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2482; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2483; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2484; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2485; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2486; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2487; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2488; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2489; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2490; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2491; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2492; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2493; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2494; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2495; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2497; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2498; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2499; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2500; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2501; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2502; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2503; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2504; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2505; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2506; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2507; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2508; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2509; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2510; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2511; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2512; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2513; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2514; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2515; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2516; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2517; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2518; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2519; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2520; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2521; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2522; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2523; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2524; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2525; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2526; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2527; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2528; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2529; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2530; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2531; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2532; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2533; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2534; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2535; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2536; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2537; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2538; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2539; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2540; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2541; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2542; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2543; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2544; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2545; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2546; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2547; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2548; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2549; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2550; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2551; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2552; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2553; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2554; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2555; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2556; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2557; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2558; // @[execute.scala 79:10:@1990.4]
  wire  _GEN_2559; // @[execute.scala 79:10:@1990.4]
  wire  _T_394; // @[execute.scala 79:10:@1990.4]
  wire  _T_396; // @[execute.scala 79:15:@1991.4]
  wire [6:0] _T_398; // @[execute.scala 79:37:@1992.4]
  wire [6:0] _T_399; // @[execute.scala 79:37:@1993.4]
  wire [5:0] _T_400; // @[execute.scala 79:37:@1994.4]
  wire [6:0] _T_403; // @[execute.scala 79:60:@1995.4]
  wire [5:0] _T_404; // @[execute.scala 79:60:@1996.4]
  wire  _GEN_2561; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2562; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2563; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2564; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2565; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2566; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2567; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2568; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2569; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2570; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2571; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2572; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2573; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2574; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2575; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2576; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2577; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2578; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2579; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2580; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2581; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2582; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2583; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2584; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2585; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2586; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2587; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2588; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2589; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2590; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2591; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2592; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2593; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2594; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2595; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2596; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2597; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2598; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2599; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2600; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2601; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2602; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2603; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2604; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2605; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2606; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2607; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2608; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2609; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2610; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2611; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2612; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2613; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2614; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2615; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2616; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2617; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2618; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2619; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2620; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2621; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2622; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2623; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2625; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2626; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2627; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2628; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2629; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2630; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2631; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2632; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2633; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2634; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2635; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2636; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2637; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2638; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2639; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2640; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2641; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2642; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2643; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2644; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2645; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2646; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2647; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2648; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2649; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2650; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2651; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2652; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2653; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2654; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2655; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2656; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2657; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2658; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2659; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2660; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2661; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2662; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2663; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2664; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2665; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2666; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2667; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2668; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2669; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2670; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2671; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2672; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2673; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2674; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2675; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2676; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2677; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2678; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2679; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2680; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2681; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2682; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2683; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2684; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2685; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2686; // @[execute.scala 79:10:@1997.4]
  wire  _GEN_2687; // @[execute.scala 79:10:@1997.4]
  wire  _T_406; // @[execute.scala 79:10:@1997.4]
  wire  _T_408; // @[execute.scala 79:15:@1998.4]
  wire [6:0] _T_410; // @[execute.scala 79:37:@1999.4]
  wire [6:0] _T_411; // @[execute.scala 79:37:@2000.4]
  wire [5:0] _T_412; // @[execute.scala 79:37:@2001.4]
  wire [6:0] _T_415; // @[execute.scala 79:60:@2002.4]
  wire [5:0] _T_416; // @[execute.scala 79:60:@2003.4]
  wire  _GEN_2689; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2690; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2691; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2692; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2693; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2694; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2695; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2696; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2697; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2698; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2699; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2700; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2701; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2702; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2703; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2704; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2705; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2706; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2707; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2708; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2709; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2710; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2711; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2712; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2713; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2714; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2715; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2716; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2717; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2718; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2719; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2720; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2721; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2722; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2723; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2724; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2725; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2726; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2727; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2728; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2729; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2730; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2731; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2732; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2733; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2734; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2735; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2736; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2737; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2738; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2739; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2740; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2741; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2742; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2743; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2744; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2745; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2746; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2747; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2748; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2749; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2750; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2751; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2753; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2754; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2755; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2756; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2757; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2758; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2759; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2760; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2761; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2762; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2763; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2764; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2765; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2766; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2767; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2768; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2769; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2770; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2771; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2772; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2773; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2774; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2775; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2776; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2777; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2778; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2779; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2780; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2781; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2782; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2783; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2784; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2785; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2786; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2787; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2788; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2789; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2790; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2791; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2792; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2793; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2794; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2795; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2796; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2797; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2798; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2799; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2800; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2801; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2802; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2803; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2804; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2805; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2806; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2807; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2808; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2809; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2810; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2811; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2812; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2813; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2814; // @[execute.scala 79:10:@2004.4]
  wire  _GEN_2815; // @[execute.scala 79:10:@2004.4]
  wire  _T_418; // @[execute.scala 79:10:@2004.4]
  wire  _T_420; // @[execute.scala 79:15:@2005.4]
  wire [6:0] _T_422; // @[execute.scala 79:37:@2006.4]
  wire [6:0] _T_423; // @[execute.scala 79:37:@2007.4]
  wire [5:0] _T_424; // @[execute.scala 79:37:@2008.4]
  wire [6:0] _T_427; // @[execute.scala 79:60:@2009.4]
  wire [5:0] _T_428; // @[execute.scala 79:60:@2010.4]
  wire  _GEN_2817; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2818; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2819; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2820; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2821; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2822; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2823; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2824; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2825; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2826; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2827; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2828; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2829; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2830; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2831; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2832; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2833; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2834; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2835; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2836; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2837; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2838; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2839; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2840; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2841; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2842; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2843; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2844; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2845; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2846; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2847; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2848; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2849; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2850; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2851; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2852; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2853; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2854; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2855; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2856; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2857; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2858; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2859; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2860; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2861; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2862; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2863; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2864; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2865; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2866; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2867; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2868; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2869; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2870; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2871; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2872; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2873; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2874; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2875; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2876; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2877; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2878; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2879; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2881; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2882; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2883; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2884; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2885; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2886; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2887; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2888; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2889; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2890; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2891; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2892; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2893; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2894; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2895; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2896; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2897; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2898; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2899; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2900; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2901; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2902; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2903; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2904; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2905; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2906; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2907; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2908; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2909; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2910; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2911; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2912; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2913; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2914; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2915; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2916; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2917; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2918; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2919; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2920; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2921; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2922; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2923; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2924; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2925; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2926; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2927; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2928; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2929; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2930; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2931; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2932; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2933; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2934; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2935; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2936; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2937; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2938; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2939; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2940; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2941; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2942; // @[execute.scala 79:10:@2011.4]
  wire  _GEN_2943; // @[execute.scala 79:10:@2011.4]
  wire  _T_430; // @[execute.scala 79:10:@2011.4]
  wire  _T_432; // @[execute.scala 79:15:@2012.4]
  wire [6:0] _T_434; // @[execute.scala 79:37:@2013.4]
  wire [6:0] _T_435; // @[execute.scala 79:37:@2014.4]
  wire [5:0] _T_436; // @[execute.scala 79:37:@2015.4]
  wire [6:0] _T_439; // @[execute.scala 79:60:@2016.4]
  wire [5:0] _T_440; // @[execute.scala 79:60:@2017.4]
  wire  _GEN_2945; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2946; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2947; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2948; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2949; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2950; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2951; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2952; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2953; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2954; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2955; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2956; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2957; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2958; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2959; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2960; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2961; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2962; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2963; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2964; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2965; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2966; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2967; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2968; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2969; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2970; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2971; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2972; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2973; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2974; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2975; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2976; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2977; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2978; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2979; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2980; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2981; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2982; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2983; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2984; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2985; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2986; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2987; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2988; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2989; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2990; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2991; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2992; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2993; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2994; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2995; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2996; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2997; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2998; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_2999; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3000; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3001; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3002; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3003; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3004; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3005; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3006; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3007; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3009; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3010; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3011; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3012; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3013; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3014; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3015; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3016; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3017; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3018; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3019; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3020; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3021; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3022; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3023; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3024; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3025; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3026; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3027; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3028; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3029; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3030; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3031; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3032; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3033; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3034; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3035; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3036; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3037; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3038; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3039; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3040; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3041; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3042; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3043; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3044; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3045; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3046; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3047; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3048; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3049; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3050; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3051; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3052; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3053; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3054; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3055; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3056; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3057; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3058; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3059; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3060; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3061; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3062; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3063; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3064; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3065; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3066; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3067; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3068; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3069; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3070; // @[execute.scala 79:10:@2018.4]
  wire  _GEN_3071; // @[execute.scala 79:10:@2018.4]
  wire  _T_442; // @[execute.scala 79:10:@2018.4]
  wire  _T_444; // @[execute.scala 79:15:@2019.4]
  wire [6:0] _T_446; // @[execute.scala 79:37:@2020.4]
  wire [6:0] _T_447; // @[execute.scala 79:37:@2021.4]
  wire [5:0] _T_448; // @[execute.scala 79:37:@2022.4]
  wire [6:0] _T_451; // @[execute.scala 79:60:@2023.4]
  wire [5:0] _T_452; // @[execute.scala 79:60:@2024.4]
  wire  _GEN_3073; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3074; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3075; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3076; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3077; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3078; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3079; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3080; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3081; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3082; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3083; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3084; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3085; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3086; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3087; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3088; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3089; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3090; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3091; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3092; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3093; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3094; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3095; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3096; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3097; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3098; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3099; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3100; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3101; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3102; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3103; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3104; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3105; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3106; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3107; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3108; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3109; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3110; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3111; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3112; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3113; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3114; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3115; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3116; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3117; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3118; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3119; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3120; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3121; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3122; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3123; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3124; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3125; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3126; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3127; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3128; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3129; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3130; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3131; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3132; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3133; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3134; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3135; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3137; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3138; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3139; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3140; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3141; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3142; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3143; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3144; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3145; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3146; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3147; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3148; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3149; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3150; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3151; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3152; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3153; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3154; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3155; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3156; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3157; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3158; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3159; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3160; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3161; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3162; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3163; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3164; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3165; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3166; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3167; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3168; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3169; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3170; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3171; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3172; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3173; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3174; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3175; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3176; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3177; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3178; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3179; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3180; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3181; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3182; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3183; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3184; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3185; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3186; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3187; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3188; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3189; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3190; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3191; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3192; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3193; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3194; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3195; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3196; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3197; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3198; // @[execute.scala 79:10:@2025.4]
  wire  _GEN_3199; // @[execute.scala 79:10:@2025.4]
  wire  _T_454; // @[execute.scala 79:10:@2025.4]
  wire  _T_456; // @[execute.scala 79:15:@2026.4]
  wire [6:0] _T_458; // @[execute.scala 79:37:@2027.4]
  wire [6:0] _T_459; // @[execute.scala 79:37:@2028.4]
  wire [5:0] _T_460; // @[execute.scala 79:37:@2029.4]
  wire [6:0] _T_463; // @[execute.scala 79:60:@2030.4]
  wire [5:0] _T_464; // @[execute.scala 79:60:@2031.4]
  wire  _GEN_3201; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3202; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3203; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3204; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3205; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3206; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3207; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3208; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3209; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3210; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3211; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3212; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3213; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3214; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3215; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3216; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3217; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3218; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3219; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3220; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3221; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3222; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3223; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3224; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3225; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3226; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3227; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3228; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3229; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3230; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3231; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3232; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3233; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3234; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3235; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3236; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3237; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3238; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3239; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3240; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3241; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3242; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3243; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3244; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3245; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3246; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3247; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3248; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3249; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3250; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3251; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3252; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3253; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3254; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3255; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3256; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3257; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3258; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3259; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3260; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3261; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3262; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3263; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3265; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3266; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3267; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3268; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3269; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3270; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3271; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3272; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3273; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3274; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3275; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3276; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3277; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3278; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3279; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3280; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3281; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3282; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3283; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3284; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3285; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3286; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3287; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3288; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3289; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3290; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3291; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3292; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3293; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3294; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3295; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3296; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3297; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3298; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3299; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3300; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3301; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3302; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3303; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3304; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3305; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3306; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3307; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3308; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3309; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3310; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3311; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3312; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3313; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3314; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3315; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3316; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3317; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3318; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3319; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3320; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3321; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3322; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3323; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3324; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3325; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3326; // @[execute.scala 79:10:@2032.4]
  wire  _GEN_3327; // @[execute.scala 79:10:@2032.4]
  wire  _T_466; // @[execute.scala 79:10:@2032.4]
  wire  _T_468; // @[execute.scala 79:15:@2033.4]
  wire [6:0] _T_470; // @[execute.scala 79:37:@2034.4]
  wire [6:0] _T_471; // @[execute.scala 79:37:@2035.4]
  wire [5:0] _T_472; // @[execute.scala 79:37:@2036.4]
  wire [6:0] _T_475; // @[execute.scala 79:60:@2037.4]
  wire [5:0] _T_476; // @[execute.scala 79:60:@2038.4]
  wire  _GEN_3329; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3330; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3331; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3332; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3333; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3334; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3335; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3336; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3337; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3338; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3339; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3340; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3341; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3342; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3343; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3344; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3345; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3346; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3347; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3348; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3349; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3350; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3351; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3352; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3353; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3354; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3355; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3356; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3357; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3358; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3359; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3360; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3361; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3362; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3363; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3364; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3365; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3366; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3367; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3368; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3369; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3370; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3371; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3372; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3373; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3374; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3375; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3376; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3377; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3378; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3379; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3380; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3381; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3382; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3383; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3384; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3385; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3386; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3387; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3388; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3389; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3390; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3391; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3393; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3394; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3395; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3396; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3397; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3398; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3399; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3400; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3401; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3402; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3403; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3404; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3405; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3406; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3407; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3408; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3409; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3410; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3411; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3412; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3413; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3414; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3415; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3416; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3417; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3418; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3419; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3420; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3421; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3422; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3423; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3424; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3425; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3426; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3427; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3428; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3429; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3430; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3431; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3432; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3433; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3434; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3435; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3436; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3437; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3438; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3439; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3440; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3441; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3442; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3443; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3444; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3445; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3446; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3447; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3448; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3449; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3450; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3451; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3452; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3453; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3454; // @[execute.scala 79:10:@2039.4]
  wire  _GEN_3455; // @[execute.scala 79:10:@2039.4]
  wire  _T_478; // @[execute.scala 79:10:@2039.4]
  wire  _T_480; // @[execute.scala 79:15:@2040.4]
  wire [6:0] _T_482; // @[execute.scala 79:37:@2041.4]
  wire [6:0] _T_483; // @[execute.scala 79:37:@2042.4]
  wire [5:0] _T_484; // @[execute.scala 79:37:@2043.4]
  wire [6:0] _T_487; // @[execute.scala 79:60:@2044.4]
  wire [5:0] _T_488; // @[execute.scala 79:60:@2045.4]
  wire  _GEN_3457; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3458; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3459; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3460; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3461; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3462; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3463; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3464; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3465; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3466; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3467; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3468; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3469; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3470; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3471; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3472; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3473; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3474; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3475; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3476; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3477; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3478; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3479; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3480; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3481; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3482; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3483; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3484; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3485; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3486; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3487; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3488; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3489; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3490; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3491; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3492; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3493; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3494; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3495; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3496; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3497; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3498; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3499; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3500; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3501; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3502; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3503; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3504; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3505; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3506; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3507; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3508; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3509; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3510; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3511; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3512; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3513; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3514; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3515; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3516; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3517; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3518; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3519; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3521; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3522; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3523; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3524; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3525; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3526; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3527; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3528; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3529; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3530; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3531; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3532; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3533; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3534; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3535; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3536; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3537; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3538; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3539; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3540; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3541; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3542; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3543; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3544; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3545; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3546; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3547; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3548; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3549; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3550; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3551; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3552; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3553; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3554; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3555; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3556; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3557; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3558; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3559; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3560; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3561; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3562; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3563; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3564; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3565; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3566; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3567; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3568; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3569; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3570; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3571; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3572; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3573; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3574; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3575; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3576; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3577; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3578; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3579; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3580; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3581; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3582; // @[execute.scala 79:10:@2046.4]
  wire  _GEN_3583; // @[execute.scala 79:10:@2046.4]
  wire  _T_490; // @[execute.scala 79:10:@2046.4]
  wire  _T_492; // @[execute.scala 79:15:@2047.4]
  wire [6:0] _T_494; // @[execute.scala 79:37:@2048.4]
  wire [6:0] _T_495; // @[execute.scala 79:37:@2049.4]
  wire [5:0] _T_496; // @[execute.scala 79:37:@2050.4]
  wire [6:0] _T_499; // @[execute.scala 79:60:@2051.4]
  wire [5:0] _T_500; // @[execute.scala 79:60:@2052.4]
  wire  _GEN_3585; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3586; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3587; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3588; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3589; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3590; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3591; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3592; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3593; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3594; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3595; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3596; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3597; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3598; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3599; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3600; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3601; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3602; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3603; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3604; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3605; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3606; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3607; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3608; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3609; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3610; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3611; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3612; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3613; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3614; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3615; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3616; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3617; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3618; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3619; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3620; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3621; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3622; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3623; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3624; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3625; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3626; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3627; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3628; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3629; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3630; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3631; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3632; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3633; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3634; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3635; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3636; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3637; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3638; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3639; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3640; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3641; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3642; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3643; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3644; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3645; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3646; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3647; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3649; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3650; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3651; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3652; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3653; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3654; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3655; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3656; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3657; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3658; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3659; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3660; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3661; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3662; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3663; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3664; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3665; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3666; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3667; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3668; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3669; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3670; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3671; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3672; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3673; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3674; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3675; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3676; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3677; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3678; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3679; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3680; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3681; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3682; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3683; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3684; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3685; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3686; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3687; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3688; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3689; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3690; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3691; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3692; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3693; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3694; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3695; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3696; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3697; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3698; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3699; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3700; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3701; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3702; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3703; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3704; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3705; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3706; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3707; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3708; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3709; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3710; // @[execute.scala 79:10:@2053.4]
  wire  _GEN_3711; // @[execute.scala 79:10:@2053.4]
  wire  _T_502; // @[execute.scala 79:10:@2053.4]
  wire  _T_504; // @[execute.scala 79:15:@2054.4]
  wire [6:0] _T_506; // @[execute.scala 79:37:@2055.4]
  wire [6:0] _T_507; // @[execute.scala 79:37:@2056.4]
  wire [5:0] _T_508; // @[execute.scala 79:37:@2057.4]
  wire [6:0] _T_511; // @[execute.scala 79:60:@2058.4]
  wire [5:0] _T_512; // @[execute.scala 79:60:@2059.4]
  wire  _GEN_3713; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3714; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3715; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3716; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3717; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3718; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3719; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3720; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3721; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3722; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3723; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3724; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3725; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3726; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3727; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3728; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3729; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3730; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3731; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3732; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3733; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3734; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3735; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3736; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3737; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3738; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3739; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3740; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3741; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3742; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3743; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3744; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3745; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3746; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3747; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3748; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3749; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3750; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3751; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3752; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3753; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3754; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3755; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3756; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3757; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3758; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3759; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3760; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3761; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3762; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3763; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3764; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3765; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3766; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3767; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3768; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3769; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3770; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3771; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3772; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3773; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3774; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3775; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3777; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3778; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3779; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3780; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3781; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3782; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3783; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3784; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3785; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3786; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3787; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3788; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3789; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3790; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3791; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3792; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3793; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3794; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3795; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3796; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3797; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3798; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3799; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3800; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3801; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3802; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3803; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3804; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3805; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3806; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3807; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3808; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3809; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3810; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3811; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3812; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3813; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3814; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3815; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3816; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3817; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3818; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3819; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3820; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3821; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3822; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3823; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3824; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3825; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3826; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3827; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3828; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3829; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3830; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3831; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3832; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3833; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3834; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3835; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3836; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3837; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3838; // @[execute.scala 79:10:@2060.4]
  wire  _GEN_3839; // @[execute.scala 79:10:@2060.4]
  wire  _T_514; // @[execute.scala 79:10:@2060.4]
  wire  _T_516; // @[execute.scala 79:15:@2061.4]
  wire [6:0] _T_518; // @[execute.scala 79:37:@2062.4]
  wire [6:0] _T_519; // @[execute.scala 79:37:@2063.4]
  wire [5:0] _T_520; // @[execute.scala 79:37:@2064.4]
  wire [6:0] _T_523; // @[execute.scala 79:60:@2065.4]
  wire [5:0] _T_524; // @[execute.scala 79:60:@2066.4]
  wire  _GEN_3841; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3842; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3843; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3844; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3845; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3846; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3847; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3848; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3849; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3850; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3851; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3852; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3853; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3854; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3855; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3856; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3857; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3858; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3859; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3860; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3861; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3862; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3863; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3864; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3865; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3866; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3867; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3868; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3869; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3870; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3871; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3872; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3873; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3874; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3875; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3876; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3877; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3878; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3879; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3880; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3881; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3882; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3883; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3884; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3885; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3886; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3887; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3888; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3889; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3890; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3891; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3892; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3893; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3894; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3895; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3896; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3897; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3898; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3899; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3900; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3901; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3902; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3903; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3905; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3906; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3907; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3908; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3909; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3910; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3911; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3912; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3913; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3914; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3915; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3916; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3917; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3918; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3919; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3920; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3921; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3922; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3923; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3924; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3925; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3926; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3927; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3928; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3929; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3930; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3931; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3932; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3933; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3934; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3935; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3936; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3937; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3938; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3939; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3940; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3941; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3942; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3943; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3944; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3945; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3946; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3947; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3948; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3949; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3950; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3951; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3952; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3953; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3954; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3955; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3956; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3957; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3958; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3959; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3960; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3961; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3962; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3963; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3964; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3965; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3966; // @[execute.scala 79:10:@2067.4]
  wire  _GEN_3967; // @[execute.scala 79:10:@2067.4]
  wire  _T_526; // @[execute.scala 79:10:@2067.4]
  wire  _T_528; // @[execute.scala 79:15:@2068.4]
  wire [6:0] _T_530; // @[execute.scala 79:37:@2069.4]
  wire [6:0] _T_531; // @[execute.scala 79:37:@2070.4]
  wire [5:0] _T_532; // @[execute.scala 79:37:@2071.4]
  wire [6:0] _T_535; // @[execute.scala 79:60:@2072.4]
  wire [5:0] _T_536; // @[execute.scala 79:60:@2073.4]
  wire  _GEN_3969; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3970; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3971; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3972; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3973; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3974; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3975; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3976; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3977; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3978; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3979; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3980; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3981; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3982; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3983; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3984; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3985; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3986; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3987; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3988; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3989; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3990; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3991; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3992; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3993; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3994; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3995; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3996; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3997; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3998; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_3999; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4000; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4001; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4002; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4003; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4004; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4005; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4006; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4007; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4008; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4009; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4010; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4011; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4012; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4013; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4014; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4015; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4016; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4017; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4018; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4019; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4020; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4021; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4022; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4023; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4024; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4025; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4026; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4027; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4028; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4029; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4030; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4031; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4033; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4034; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4035; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4036; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4037; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4038; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4039; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4040; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4041; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4042; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4043; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4044; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4045; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4046; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4047; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4048; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4049; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4050; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4051; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4052; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4053; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4054; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4055; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4056; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4057; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4058; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4059; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4060; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4061; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4062; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4063; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4064; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4065; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4066; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4067; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4068; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4069; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4070; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4071; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4072; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4073; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4074; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4075; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4076; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4077; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4078; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4079; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4080; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4081; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4082; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4083; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4084; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4085; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4086; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4087; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4088; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4089; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4090; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4091; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4092; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4093; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4094; // @[execute.scala 79:10:@2074.4]
  wire  _GEN_4095; // @[execute.scala 79:10:@2074.4]
  wire  _T_538; // @[execute.scala 79:10:@2074.4]
  wire  _T_540; // @[execute.scala 79:15:@2075.4]
  wire [6:0] _T_542; // @[execute.scala 79:37:@2076.4]
  wire [6:0] _T_543; // @[execute.scala 79:37:@2077.4]
  wire [5:0] _T_544; // @[execute.scala 79:37:@2078.4]
  wire [6:0] _T_547; // @[execute.scala 79:60:@2079.4]
  wire [5:0] _T_548; // @[execute.scala 79:60:@2080.4]
  wire  _GEN_4097; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4098; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4099; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4100; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4101; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4102; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4103; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4104; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4105; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4106; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4107; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4108; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4109; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4110; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4111; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4112; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4113; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4114; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4115; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4116; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4117; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4118; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4119; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4120; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4121; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4122; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4123; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4124; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4125; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4126; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4127; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4128; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4129; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4130; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4131; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4132; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4133; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4134; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4135; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4136; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4137; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4138; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4139; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4140; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4141; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4142; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4143; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4144; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4145; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4146; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4147; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4148; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4149; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4150; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4151; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4152; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4153; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4154; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4155; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4156; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4157; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4158; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4159; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4161; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4162; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4163; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4164; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4165; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4166; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4167; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4168; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4169; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4170; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4171; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4172; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4173; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4174; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4175; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4176; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4177; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4178; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4179; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4180; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4181; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4182; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4183; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4184; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4185; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4186; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4187; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4188; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4189; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4190; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4191; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4192; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4193; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4194; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4195; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4196; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4197; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4198; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4199; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4200; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4201; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4202; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4203; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4204; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4205; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4206; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4207; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4208; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4209; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4210; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4211; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4212; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4213; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4214; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4215; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4216; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4217; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4218; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4219; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4220; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4221; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4222; // @[execute.scala 79:10:@2081.4]
  wire  _GEN_4223; // @[execute.scala 79:10:@2081.4]
  wire  _T_550; // @[execute.scala 79:10:@2081.4]
  wire  _T_552; // @[execute.scala 79:15:@2082.4]
  wire [6:0] _T_554; // @[execute.scala 79:37:@2083.4]
  wire [6:0] _T_555; // @[execute.scala 79:37:@2084.4]
  wire [5:0] _T_556; // @[execute.scala 79:37:@2085.4]
  wire [6:0] _T_559; // @[execute.scala 79:60:@2086.4]
  wire [5:0] _T_560; // @[execute.scala 79:60:@2087.4]
  wire  _GEN_4225; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4226; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4227; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4228; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4229; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4230; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4231; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4232; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4233; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4234; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4235; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4236; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4237; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4238; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4239; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4240; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4241; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4242; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4243; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4244; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4245; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4246; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4247; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4248; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4249; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4250; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4251; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4252; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4253; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4254; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4255; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4256; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4257; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4258; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4259; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4260; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4261; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4262; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4263; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4264; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4265; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4266; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4267; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4268; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4269; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4270; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4271; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4272; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4273; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4274; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4275; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4276; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4277; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4278; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4279; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4280; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4281; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4282; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4283; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4284; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4285; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4286; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4287; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4289; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4290; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4291; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4292; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4293; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4294; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4295; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4296; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4297; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4298; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4299; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4300; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4301; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4302; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4303; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4304; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4305; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4306; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4307; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4308; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4309; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4310; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4311; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4312; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4313; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4314; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4315; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4316; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4317; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4318; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4319; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4320; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4321; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4322; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4323; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4324; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4325; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4326; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4327; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4328; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4329; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4330; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4331; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4332; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4333; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4334; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4335; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4336; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4337; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4338; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4339; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4340; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4341; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4342; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4343; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4344; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4345; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4346; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4347; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4348; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4349; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4350; // @[execute.scala 79:10:@2088.4]
  wire  _GEN_4351; // @[execute.scala 79:10:@2088.4]
  wire  _T_562; // @[execute.scala 79:10:@2088.4]
  wire  _T_564; // @[execute.scala 79:15:@2089.4]
  wire [6:0] _T_566; // @[execute.scala 79:37:@2090.4]
  wire [6:0] _T_567; // @[execute.scala 79:37:@2091.4]
  wire [5:0] _T_568; // @[execute.scala 79:37:@2092.4]
  wire [6:0] _T_571; // @[execute.scala 79:60:@2093.4]
  wire [5:0] _T_572; // @[execute.scala 79:60:@2094.4]
  wire  _GEN_4353; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4354; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4355; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4356; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4357; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4358; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4359; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4360; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4361; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4362; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4363; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4364; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4365; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4366; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4367; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4368; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4369; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4370; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4371; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4372; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4373; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4374; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4375; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4376; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4377; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4378; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4379; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4380; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4381; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4382; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4383; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4384; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4385; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4386; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4387; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4388; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4389; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4390; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4391; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4392; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4393; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4394; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4395; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4396; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4397; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4398; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4399; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4400; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4401; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4402; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4403; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4404; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4405; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4406; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4407; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4408; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4409; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4410; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4411; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4412; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4413; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4414; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4415; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4417; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4418; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4419; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4420; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4421; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4422; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4423; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4424; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4425; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4426; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4427; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4428; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4429; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4430; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4431; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4432; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4433; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4434; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4435; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4436; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4437; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4438; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4439; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4440; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4441; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4442; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4443; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4444; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4445; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4446; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4447; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4448; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4449; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4450; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4451; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4452; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4453; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4454; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4455; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4456; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4457; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4458; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4459; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4460; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4461; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4462; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4463; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4464; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4465; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4466; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4467; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4468; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4469; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4470; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4471; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4472; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4473; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4474; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4475; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4476; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4477; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4478; // @[execute.scala 79:10:@2095.4]
  wire  _GEN_4479; // @[execute.scala 79:10:@2095.4]
  wire  _T_574; // @[execute.scala 79:10:@2095.4]
  wire  _T_576; // @[execute.scala 79:15:@2096.4]
  wire [6:0] _T_578; // @[execute.scala 79:37:@2097.4]
  wire [6:0] _T_579; // @[execute.scala 79:37:@2098.4]
  wire [5:0] _T_580; // @[execute.scala 79:37:@2099.4]
  wire [6:0] _T_583; // @[execute.scala 79:60:@2100.4]
  wire [5:0] _T_584; // @[execute.scala 79:60:@2101.4]
  wire  _GEN_4481; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4482; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4483; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4484; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4485; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4486; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4487; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4488; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4489; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4490; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4491; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4492; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4493; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4494; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4495; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4496; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4497; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4498; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4499; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4500; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4501; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4502; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4503; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4504; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4505; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4506; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4507; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4508; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4509; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4510; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4511; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4512; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4513; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4514; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4515; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4516; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4517; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4518; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4519; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4520; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4521; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4522; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4523; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4524; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4525; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4526; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4527; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4528; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4529; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4530; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4531; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4532; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4533; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4534; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4535; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4536; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4537; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4538; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4539; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4540; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4541; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4542; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4543; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4545; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4546; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4547; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4548; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4549; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4550; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4551; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4552; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4553; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4554; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4555; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4556; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4557; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4558; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4559; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4560; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4561; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4562; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4563; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4564; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4565; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4566; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4567; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4568; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4569; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4570; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4571; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4572; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4573; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4574; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4575; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4576; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4577; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4578; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4579; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4580; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4581; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4582; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4583; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4584; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4585; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4586; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4587; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4588; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4589; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4590; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4591; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4592; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4593; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4594; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4595; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4596; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4597; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4598; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4599; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4600; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4601; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4602; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4603; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4604; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4605; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4606; // @[execute.scala 79:10:@2102.4]
  wire  _GEN_4607; // @[execute.scala 79:10:@2102.4]
  wire  _T_586; // @[execute.scala 79:10:@2102.4]
  wire  _T_588; // @[execute.scala 79:15:@2103.4]
  wire [6:0] _T_590; // @[execute.scala 79:37:@2104.4]
  wire [6:0] _T_591; // @[execute.scala 79:37:@2105.4]
  wire [5:0] _T_592; // @[execute.scala 79:37:@2106.4]
  wire [6:0] _T_595; // @[execute.scala 79:60:@2107.4]
  wire [5:0] _T_596; // @[execute.scala 79:60:@2108.4]
  wire  _GEN_4609; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4610; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4611; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4612; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4613; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4614; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4615; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4616; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4617; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4618; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4619; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4620; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4621; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4622; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4623; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4624; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4625; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4626; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4627; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4628; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4629; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4630; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4631; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4632; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4633; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4634; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4635; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4636; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4637; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4638; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4639; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4640; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4641; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4642; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4643; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4644; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4645; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4646; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4647; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4648; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4649; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4650; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4651; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4652; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4653; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4654; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4655; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4656; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4657; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4658; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4659; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4660; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4661; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4662; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4663; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4664; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4665; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4666; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4667; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4668; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4669; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4670; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4671; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4673; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4674; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4675; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4676; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4677; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4678; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4679; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4680; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4681; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4682; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4683; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4684; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4685; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4686; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4687; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4688; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4689; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4690; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4691; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4692; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4693; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4694; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4695; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4696; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4697; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4698; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4699; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4700; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4701; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4702; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4703; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4704; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4705; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4706; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4707; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4708; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4709; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4710; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4711; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4712; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4713; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4714; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4715; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4716; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4717; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4718; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4719; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4720; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4721; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4722; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4723; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4724; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4725; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4726; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4727; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4728; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4729; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4730; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4731; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4732; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4733; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4734; // @[execute.scala 79:10:@2109.4]
  wire  _GEN_4735; // @[execute.scala 79:10:@2109.4]
  wire  _T_598; // @[execute.scala 79:10:@2109.4]
  wire  _T_600; // @[execute.scala 79:15:@2110.4]
  wire [6:0] _T_602; // @[execute.scala 79:37:@2111.4]
  wire [6:0] _T_603; // @[execute.scala 79:37:@2112.4]
  wire [5:0] _T_604; // @[execute.scala 79:37:@2113.4]
  wire [6:0] _T_607; // @[execute.scala 79:60:@2114.4]
  wire [5:0] _T_608; // @[execute.scala 79:60:@2115.4]
  wire  _GEN_4737; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4738; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4739; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4740; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4741; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4742; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4743; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4744; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4745; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4746; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4747; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4748; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4749; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4750; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4751; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4752; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4753; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4754; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4755; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4756; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4757; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4758; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4759; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4760; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4761; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4762; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4763; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4764; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4765; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4766; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4767; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4768; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4769; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4770; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4771; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4772; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4773; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4774; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4775; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4776; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4777; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4778; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4779; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4780; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4781; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4782; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4783; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4784; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4785; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4786; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4787; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4788; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4789; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4790; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4791; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4792; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4793; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4794; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4795; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4796; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4797; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4798; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4799; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4801; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4802; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4803; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4804; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4805; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4806; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4807; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4808; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4809; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4810; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4811; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4812; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4813; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4814; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4815; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4816; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4817; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4818; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4819; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4820; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4821; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4822; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4823; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4824; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4825; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4826; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4827; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4828; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4829; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4830; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4831; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4832; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4833; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4834; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4835; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4836; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4837; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4838; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4839; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4840; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4841; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4842; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4843; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4844; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4845; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4846; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4847; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4848; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4849; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4850; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4851; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4852; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4853; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4854; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4855; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4856; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4857; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4858; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4859; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4860; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4861; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4862; // @[execute.scala 79:10:@2116.4]
  wire  _GEN_4863; // @[execute.scala 79:10:@2116.4]
  wire  _T_610; // @[execute.scala 79:10:@2116.4]
  wire  _T_612; // @[execute.scala 79:15:@2117.4]
  wire [6:0] _T_614; // @[execute.scala 79:37:@2118.4]
  wire [6:0] _T_615; // @[execute.scala 79:37:@2119.4]
  wire [5:0] _T_616; // @[execute.scala 79:37:@2120.4]
  wire [6:0] _T_619; // @[execute.scala 79:60:@2121.4]
  wire [5:0] _T_620; // @[execute.scala 79:60:@2122.4]
  wire  _GEN_4865; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4866; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4867; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4868; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4869; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4870; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4871; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4872; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4873; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4874; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4875; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4876; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4877; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4878; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4879; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4880; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4881; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4882; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4883; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4884; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4885; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4886; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4887; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4888; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4889; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4890; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4891; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4892; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4893; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4894; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4895; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4896; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4897; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4898; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4899; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4900; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4901; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4902; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4903; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4904; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4905; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4906; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4907; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4908; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4909; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4910; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4911; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4912; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4913; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4914; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4915; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4916; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4917; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4918; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4919; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4920; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4921; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4922; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4923; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4924; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4925; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4926; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4927; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4929; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4930; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4931; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4932; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4933; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4934; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4935; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4936; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4937; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4938; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4939; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4940; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4941; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4942; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4943; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4944; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4945; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4946; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4947; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4948; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4949; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4950; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4951; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4952; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4953; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4954; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4955; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4956; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4957; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4958; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4959; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4960; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4961; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4962; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4963; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4964; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4965; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4966; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4967; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4968; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4969; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4970; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4971; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4972; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4973; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4974; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4975; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4976; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4977; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4978; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4979; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4980; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4981; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4982; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4983; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4984; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4985; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4986; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4987; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4988; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4989; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4990; // @[execute.scala 79:10:@2123.4]
  wire  _GEN_4991; // @[execute.scala 79:10:@2123.4]
  wire  _T_622; // @[execute.scala 79:10:@2123.4]
  wire  _T_624; // @[execute.scala 79:15:@2124.4]
  wire [6:0] _T_626; // @[execute.scala 79:37:@2125.4]
  wire [6:0] _T_627; // @[execute.scala 79:37:@2126.4]
  wire [5:0] _T_628; // @[execute.scala 79:37:@2127.4]
  wire [6:0] _T_631; // @[execute.scala 79:60:@2128.4]
  wire [5:0] _T_632; // @[execute.scala 79:60:@2129.4]
  wire  _GEN_4993; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_4994; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_4995; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_4996; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_4997; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_4998; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_4999; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5000; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5001; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5002; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5003; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5004; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5005; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5006; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5007; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5008; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5009; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5010; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5011; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5012; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5013; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5014; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5015; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5016; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5017; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5018; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5019; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5020; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5021; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5022; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5023; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5024; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5025; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5026; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5027; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5028; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5029; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5030; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5031; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5032; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5033; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5034; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5035; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5036; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5037; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5038; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5039; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5040; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5041; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5042; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5043; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5044; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5045; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5046; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5047; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5048; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5049; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5050; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5051; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5052; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5053; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5054; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5055; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5057; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5058; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5059; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5060; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5061; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5062; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5063; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5064; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5065; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5066; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5067; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5068; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5069; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5070; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5071; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5072; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5073; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5074; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5075; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5076; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5077; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5078; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5079; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5080; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5081; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5082; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5083; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5084; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5085; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5086; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5087; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5088; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5089; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5090; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5091; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5092; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5093; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5094; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5095; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5096; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5097; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5098; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5099; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5100; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5101; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5102; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5103; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5104; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5105; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5106; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5107; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5108; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5109; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5110; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5111; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5112; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5113; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5114; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5115; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5116; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5117; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5118; // @[execute.scala 79:10:@2130.4]
  wire  _GEN_5119; // @[execute.scala 79:10:@2130.4]
  wire  _T_634; // @[execute.scala 79:10:@2130.4]
  wire  _T_636; // @[execute.scala 79:15:@2131.4]
  wire [6:0] _T_638; // @[execute.scala 79:37:@2132.4]
  wire [6:0] _T_639; // @[execute.scala 79:37:@2133.4]
  wire [5:0] _T_640; // @[execute.scala 79:37:@2134.4]
  wire [6:0] _T_643; // @[execute.scala 79:60:@2135.4]
  wire [5:0] _T_644; // @[execute.scala 79:60:@2136.4]
  wire  _GEN_5121; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5122; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5123; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5124; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5125; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5126; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5127; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5128; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5129; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5130; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5131; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5132; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5133; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5134; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5135; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5136; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5137; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5138; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5139; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5140; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5141; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5142; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5143; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5144; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5145; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5146; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5147; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5148; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5149; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5150; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5151; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5152; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5153; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5154; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5155; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5156; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5157; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5158; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5159; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5160; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5161; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5162; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5163; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5164; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5165; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5166; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5167; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5168; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5169; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5170; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5171; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5172; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5173; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5174; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5175; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5176; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5177; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5178; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5179; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5180; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5181; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5182; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5183; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5185; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5186; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5187; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5188; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5189; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5190; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5191; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5192; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5193; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5194; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5195; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5196; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5197; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5198; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5199; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5200; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5201; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5202; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5203; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5204; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5205; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5206; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5207; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5208; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5209; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5210; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5211; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5212; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5213; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5214; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5215; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5216; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5217; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5218; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5219; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5220; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5221; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5222; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5223; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5224; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5225; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5226; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5227; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5228; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5229; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5230; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5231; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5232; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5233; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5234; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5235; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5236; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5237; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5238; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5239; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5240; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5241; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5242; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5243; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5244; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5245; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5246; // @[execute.scala 79:10:@2137.4]
  wire  _GEN_5247; // @[execute.scala 79:10:@2137.4]
  wire  _T_646; // @[execute.scala 79:10:@2137.4]
  wire  _T_648; // @[execute.scala 79:15:@2138.4]
  wire [6:0] _T_650; // @[execute.scala 79:37:@2139.4]
  wire [6:0] _T_651; // @[execute.scala 79:37:@2140.4]
  wire [5:0] _T_652; // @[execute.scala 79:37:@2141.4]
  wire [6:0] _T_655; // @[execute.scala 79:60:@2142.4]
  wire [5:0] _T_656; // @[execute.scala 79:60:@2143.4]
  wire  _GEN_5249; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5250; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5251; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5252; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5253; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5254; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5255; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5256; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5257; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5258; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5259; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5260; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5261; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5262; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5263; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5264; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5265; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5266; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5267; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5268; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5269; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5270; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5271; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5272; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5273; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5274; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5275; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5276; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5277; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5278; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5279; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5280; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5281; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5282; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5283; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5284; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5285; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5286; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5287; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5288; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5289; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5290; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5291; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5292; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5293; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5294; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5295; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5296; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5297; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5298; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5299; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5300; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5301; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5302; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5303; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5304; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5305; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5306; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5307; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5308; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5309; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5310; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5311; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5313; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5314; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5315; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5316; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5317; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5318; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5319; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5320; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5321; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5322; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5323; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5324; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5325; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5326; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5327; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5328; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5329; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5330; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5331; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5332; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5333; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5334; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5335; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5336; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5337; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5338; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5339; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5340; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5341; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5342; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5343; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5344; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5345; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5346; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5347; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5348; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5349; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5350; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5351; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5352; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5353; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5354; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5355; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5356; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5357; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5358; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5359; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5360; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5361; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5362; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5363; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5364; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5365; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5366; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5367; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5368; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5369; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5370; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5371; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5372; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5373; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5374; // @[execute.scala 79:10:@2144.4]
  wire  _GEN_5375; // @[execute.scala 79:10:@2144.4]
  wire  _T_658; // @[execute.scala 79:10:@2144.4]
  wire  _T_660; // @[execute.scala 79:15:@2145.4]
  wire [6:0] _T_662; // @[execute.scala 79:37:@2146.4]
  wire [6:0] _T_663; // @[execute.scala 79:37:@2147.4]
  wire [5:0] _T_664; // @[execute.scala 79:37:@2148.4]
  wire [6:0] _T_667; // @[execute.scala 79:60:@2149.4]
  wire [5:0] _T_668; // @[execute.scala 79:60:@2150.4]
  wire  _GEN_5377; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5378; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5379; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5380; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5381; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5382; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5383; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5384; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5385; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5386; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5387; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5388; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5389; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5390; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5391; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5392; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5393; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5394; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5395; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5396; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5397; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5398; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5399; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5400; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5401; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5402; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5403; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5404; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5405; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5406; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5407; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5408; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5409; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5410; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5411; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5412; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5413; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5414; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5415; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5416; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5417; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5418; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5419; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5420; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5421; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5422; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5423; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5424; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5425; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5426; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5427; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5428; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5429; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5430; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5431; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5432; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5433; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5434; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5435; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5436; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5437; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5438; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5439; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5441; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5442; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5443; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5444; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5445; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5446; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5447; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5448; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5449; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5450; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5451; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5452; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5453; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5454; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5455; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5456; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5457; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5458; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5459; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5460; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5461; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5462; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5463; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5464; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5465; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5466; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5467; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5468; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5469; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5470; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5471; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5472; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5473; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5474; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5475; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5476; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5477; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5478; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5479; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5480; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5481; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5482; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5483; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5484; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5485; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5486; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5487; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5488; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5489; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5490; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5491; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5492; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5493; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5494; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5495; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5496; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5497; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5498; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5499; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5500; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5501; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5502; // @[execute.scala 79:10:@2151.4]
  wire  _GEN_5503; // @[execute.scala 79:10:@2151.4]
  wire  _T_670; // @[execute.scala 79:10:@2151.4]
  wire  _T_672; // @[execute.scala 79:15:@2152.4]
  wire [6:0] _T_674; // @[execute.scala 79:37:@2153.4]
  wire [6:0] _T_675; // @[execute.scala 79:37:@2154.4]
  wire [5:0] _T_676; // @[execute.scala 79:37:@2155.4]
  wire [6:0] _T_679; // @[execute.scala 79:60:@2156.4]
  wire [5:0] _T_680; // @[execute.scala 79:60:@2157.4]
  wire  _GEN_5505; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5506; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5507; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5508; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5509; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5510; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5511; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5512; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5513; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5514; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5515; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5516; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5517; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5518; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5519; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5520; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5521; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5522; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5523; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5524; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5525; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5526; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5527; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5528; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5529; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5530; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5531; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5532; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5533; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5534; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5535; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5536; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5537; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5538; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5539; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5540; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5541; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5542; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5543; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5544; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5545; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5546; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5547; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5548; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5549; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5550; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5551; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5552; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5553; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5554; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5555; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5556; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5557; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5558; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5559; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5560; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5561; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5562; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5563; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5564; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5565; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5566; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5567; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5569; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5570; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5571; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5572; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5573; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5574; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5575; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5576; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5577; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5578; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5579; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5580; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5581; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5582; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5583; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5584; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5585; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5586; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5587; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5588; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5589; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5590; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5591; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5592; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5593; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5594; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5595; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5596; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5597; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5598; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5599; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5600; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5601; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5602; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5603; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5604; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5605; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5606; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5607; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5608; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5609; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5610; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5611; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5612; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5613; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5614; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5615; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5616; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5617; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5618; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5619; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5620; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5621; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5622; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5623; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5624; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5625; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5626; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5627; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5628; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5629; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5630; // @[execute.scala 79:10:@2158.4]
  wire  _GEN_5631; // @[execute.scala 79:10:@2158.4]
  wire  _T_682; // @[execute.scala 79:10:@2158.4]
  wire  _T_684; // @[execute.scala 79:15:@2159.4]
  wire [6:0] _T_686; // @[execute.scala 79:37:@2160.4]
  wire [6:0] _T_687; // @[execute.scala 79:37:@2161.4]
  wire [5:0] _T_688; // @[execute.scala 79:37:@2162.4]
  wire [6:0] _T_691; // @[execute.scala 79:60:@2163.4]
  wire [5:0] _T_692; // @[execute.scala 79:60:@2164.4]
  wire  _GEN_5633; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5634; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5635; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5636; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5637; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5638; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5639; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5640; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5641; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5642; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5643; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5644; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5645; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5646; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5647; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5648; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5649; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5650; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5651; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5652; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5653; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5654; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5655; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5656; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5657; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5658; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5659; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5660; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5661; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5662; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5663; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5664; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5665; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5666; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5667; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5668; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5669; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5670; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5671; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5672; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5673; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5674; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5675; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5676; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5677; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5678; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5679; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5680; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5681; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5682; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5683; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5684; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5685; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5686; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5687; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5688; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5689; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5690; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5691; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5692; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5693; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5694; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5695; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5697; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5698; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5699; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5700; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5701; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5702; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5703; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5704; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5705; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5706; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5707; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5708; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5709; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5710; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5711; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5712; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5713; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5714; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5715; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5716; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5717; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5718; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5719; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5720; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5721; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5722; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5723; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5724; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5725; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5726; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5727; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5728; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5729; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5730; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5731; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5732; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5733; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5734; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5735; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5736; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5737; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5738; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5739; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5740; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5741; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5742; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5743; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5744; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5745; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5746; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5747; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5748; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5749; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5750; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5751; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5752; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5753; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5754; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5755; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5756; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5757; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5758; // @[execute.scala 79:10:@2165.4]
  wire  _GEN_5759; // @[execute.scala 79:10:@2165.4]
  wire  _T_694; // @[execute.scala 79:10:@2165.4]
  wire  _T_696; // @[execute.scala 79:15:@2166.4]
  wire [6:0] _T_698; // @[execute.scala 79:37:@2167.4]
  wire [6:0] _T_699; // @[execute.scala 79:37:@2168.4]
  wire [5:0] _T_700; // @[execute.scala 79:37:@2169.4]
  wire [6:0] _T_703; // @[execute.scala 79:60:@2170.4]
  wire [5:0] _T_704; // @[execute.scala 79:60:@2171.4]
  wire  _GEN_5761; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5762; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5763; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5764; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5765; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5766; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5767; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5768; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5769; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5770; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5771; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5772; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5773; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5774; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5775; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5776; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5777; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5778; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5779; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5780; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5781; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5782; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5783; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5784; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5785; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5786; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5787; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5788; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5789; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5790; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5791; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5792; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5793; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5794; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5795; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5796; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5797; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5798; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5799; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5800; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5801; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5802; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5803; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5804; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5805; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5806; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5807; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5808; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5809; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5810; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5811; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5812; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5813; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5814; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5815; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5816; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5817; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5818; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5819; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5820; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5821; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5822; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5823; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5825; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5826; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5827; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5828; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5829; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5830; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5831; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5832; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5833; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5834; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5835; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5836; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5837; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5838; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5839; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5840; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5841; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5842; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5843; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5844; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5845; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5846; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5847; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5848; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5849; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5850; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5851; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5852; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5853; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5854; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5855; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5856; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5857; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5858; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5859; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5860; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5861; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5862; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5863; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5864; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5865; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5866; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5867; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5868; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5869; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5870; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5871; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5872; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5873; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5874; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5875; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5876; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5877; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5878; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5879; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5880; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5881; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5882; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5883; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5884; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5885; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5886; // @[execute.scala 79:10:@2172.4]
  wire  _GEN_5887; // @[execute.scala 79:10:@2172.4]
  wire  _T_706; // @[execute.scala 79:10:@2172.4]
  wire  _T_708; // @[execute.scala 79:15:@2173.4]
  wire [6:0] _T_710; // @[execute.scala 79:37:@2174.4]
  wire [6:0] _T_711; // @[execute.scala 79:37:@2175.4]
  wire [5:0] _T_712; // @[execute.scala 79:37:@2176.4]
  wire [6:0] _T_715; // @[execute.scala 79:60:@2177.4]
  wire [5:0] _T_716; // @[execute.scala 79:60:@2178.4]
  wire  _GEN_5889; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5890; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5891; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5892; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5893; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5894; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5895; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5896; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5897; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5898; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5899; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5900; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5901; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5902; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5903; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5904; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5905; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5906; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5907; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5908; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5909; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5910; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5911; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5912; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5913; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5914; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5915; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5916; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5917; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5918; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5919; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5920; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5921; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5922; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5923; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5924; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5925; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5926; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5927; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5928; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5929; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5930; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5931; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5932; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5933; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5934; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5935; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5936; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5937; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5938; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5939; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5940; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5941; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5942; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5943; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5944; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5945; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5946; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5947; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5948; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5949; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5950; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5951; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5953; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5954; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5955; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5956; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5957; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5958; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5959; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5960; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5961; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5962; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5963; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5964; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5965; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5966; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5967; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5968; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5969; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5970; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5971; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5972; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5973; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5974; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5975; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5976; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5977; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5978; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5979; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5980; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5981; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5982; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5983; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5984; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5985; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5986; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5987; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5988; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5989; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5990; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5991; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5992; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5993; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5994; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5995; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5996; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5997; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5998; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_5999; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6000; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6001; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6002; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6003; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6004; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6005; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6006; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6007; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6008; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6009; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6010; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6011; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6012; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6013; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6014; // @[execute.scala 79:10:@2179.4]
  wire  _GEN_6015; // @[execute.scala 79:10:@2179.4]
  wire  _T_718; // @[execute.scala 79:10:@2179.4]
  wire  _T_720; // @[execute.scala 79:15:@2180.4]
  wire [6:0] _T_722; // @[execute.scala 79:37:@2181.4]
  wire [6:0] _T_723; // @[execute.scala 79:37:@2182.4]
  wire [5:0] _T_724; // @[execute.scala 79:37:@2183.4]
  wire [6:0] _T_727; // @[execute.scala 79:60:@2184.4]
  wire [5:0] _T_728; // @[execute.scala 79:60:@2185.4]
  wire  _GEN_6017; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6018; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6019; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6020; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6021; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6022; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6023; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6024; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6025; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6026; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6027; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6028; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6029; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6030; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6031; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6032; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6033; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6034; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6035; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6036; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6037; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6038; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6039; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6040; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6041; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6042; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6043; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6044; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6045; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6046; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6047; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6048; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6049; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6050; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6051; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6052; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6053; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6054; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6055; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6056; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6057; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6058; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6059; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6060; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6061; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6062; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6063; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6064; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6065; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6066; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6067; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6068; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6069; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6070; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6071; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6072; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6073; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6074; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6075; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6076; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6077; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6078; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6079; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6081; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6082; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6083; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6084; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6085; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6086; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6087; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6088; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6089; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6090; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6091; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6092; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6093; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6094; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6095; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6096; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6097; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6098; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6099; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6100; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6101; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6102; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6103; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6104; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6105; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6106; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6107; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6108; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6109; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6110; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6111; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6112; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6113; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6114; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6115; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6116; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6117; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6118; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6119; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6120; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6121; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6122; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6123; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6124; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6125; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6126; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6127; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6128; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6129; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6130; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6131; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6132; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6133; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6134; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6135; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6136; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6137; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6138; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6139; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6140; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6141; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6142; // @[execute.scala 79:10:@2186.4]
  wire  _GEN_6143; // @[execute.scala 79:10:@2186.4]
  wire  _T_730; // @[execute.scala 79:10:@2186.4]
  wire  _T_732; // @[execute.scala 79:15:@2187.4]
  wire [6:0] _T_734; // @[execute.scala 79:37:@2188.4]
  wire [6:0] _T_735; // @[execute.scala 79:37:@2189.4]
  wire [5:0] _T_736; // @[execute.scala 79:37:@2190.4]
  wire [6:0] _T_739; // @[execute.scala 79:60:@2191.4]
  wire [5:0] _T_740; // @[execute.scala 79:60:@2192.4]
  wire  _GEN_6145; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6146; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6147; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6148; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6149; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6150; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6151; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6152; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6153; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6154; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6155; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6156; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6157; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6158; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6159; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6160; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6161; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6162; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6163; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6164; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6165; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6166; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6167; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6168; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6169; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6170; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6171; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6172; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6173; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6174; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6175; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6176; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6177; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6178; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6179; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6180; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6181; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6182; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6183; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6184; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6185; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6186; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6187; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6188; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6189; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6190; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6191; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6192; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6193; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6194; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6195; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6196; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6197; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6198; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6199; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6200; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6201; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6202; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6203; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6204; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6205; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6206; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6207; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6209; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6210; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6211; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6212; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6213; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6214; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6215; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6216; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6217; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6218; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6219; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6220; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6221; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6222; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6223; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6224; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6225; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6226; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6227; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6228; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6229; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6230; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6231; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6232; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6233; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6234; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6235; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6236; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6237; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6238; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6239; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6240; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6241; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6242; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6243; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6244; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6245; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6246; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6247; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6248; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6249; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6250; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6251; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6252; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6253; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6254; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6255; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6256; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6257; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6258; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6259; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6260; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6261; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6262; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6263; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6264; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6265; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6266; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6267; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6268; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6269; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6270; // @[execute.scala 79:10:@2193.4]
  wire  _GEN_6271; // @[execute.scala 79:10:@2193.4]
  wire  _T_742; // @[execute.scala 79:10:@2193.4]
  wire  _T_744; // @[execute.scala 79:15:@2194.4]
  wire [6:0] _T_746; // @[execute.scala 79:37:@2195.4]
  wire [6:0] _T_747; // @[execute.scala 79:37:@2196.4]
  wire [5:0] _T_748; // @[execute.scala 79:37:@2197.4]
  wire [6:0] _T_751; // @[execute.scala 79:60:@2198.4]
  wire [5:0] _T_752; // @[execute.scala 79:60:@2199.4]
  wire  _GEN_6273; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6274; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6275; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6276; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6277; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6278; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6279; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6280; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6281; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6282; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6283; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6284; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6285; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6286; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6287; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6288; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6289; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6290; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6291; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6292; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6293; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6294; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6295; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6296; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6297; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6298; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6299; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6300; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6301; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6302; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6303; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6304; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6305; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6306; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6307; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6308; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6309; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6310; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6311; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6312; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6313; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6314; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6315; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6316; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6317; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6318; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6319; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6320; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6321; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6322; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6323; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6324; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6325; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6326; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6327; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6328; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6329; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6330; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6331; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6332; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6333; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6334; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6335; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6337; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6338; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6339; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6340; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6341; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6342; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6343; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6344; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6345; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6346; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6347; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6348; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6349; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6350; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6351; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6352; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6353; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6354; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6355; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6356; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6357; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6358; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6359; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6360; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6361; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6362; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6363; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6364; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6365; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6366; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6367; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6368; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6369; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6370; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6371; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6372; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6373; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6374; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6375; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6376; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6377; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6378; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6379; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6380; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6381; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6382; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6383; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6384; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6385; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6386; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6387; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6388; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6389; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6390; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6391; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6392; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6393; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6394; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6395; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6396; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6397; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6398; // @[execute.scala 79:10:@2200.4]
  wire  _GEN_6399; // @[execute.scala 79:10:@2200.4]
  wire  _T_754; // @[execute.scala 79:10:@2200.4]
  wire  _T_756; // @[execute.scala 79:15:@2201.4]
  wire [6:0] _T_758; // @[execute.scala 79:37:@2202.4]
  wire [6:0] _T_759; // @[execute.scala 79:37:@2203.4]
  wire [5:0] _T_760; // @[execute.scala 79:37:@2204.4]
  wire [6:0] _T_763; // @[execute.scala 79:60:@2205.4]
  wire [5:0] _T_764; // @[execute.scala 79:60:@2206.4]
  wire  _GEN_6401; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6402; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6403; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6404; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6405; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6406; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6407; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6408; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6409; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6410; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6411; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6412; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6413; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6414; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6415; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6416; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6417; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6418; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6419; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6420; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6421; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6422; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6423; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6424; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6425; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6426; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6427; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6428; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6429; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6430; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6431; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6432; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6433; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6434; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6435; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6436; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6437; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6438; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6439; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6440; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6441; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6442; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6443; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6444; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6445; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6446; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6447; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6448; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6449; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6450; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6451; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6452; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6453; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6454; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6455; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6456; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6457; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6458; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6459; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6460; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6461; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6462; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6463; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6465; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6466; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6467; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6468; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6469; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6470; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6471; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6472; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6473; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6474; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6475; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6476; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6477; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6478; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6479; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6480; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6481; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6482; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6483; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6484; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6485; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6486; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6487; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6488; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6489; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6490; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6491; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6492; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6493; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6494; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6495; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6496; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6497; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6498; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6499; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6500; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6501; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6502; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6503; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6504; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6505; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6506; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6507; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6508; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6509; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6510; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6511; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6512; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6513; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6514; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6515; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6516; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6517; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6518; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6519; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6520; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6521; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6522; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6523; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6524; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6525; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6526; // @[execute.scala 79:10:@2207.4]
  wire  _GEN_6527; // @[execute.scala 79:10:@2207.4]
  wire  _T_766; // @[execute.scala 79:10:@2207.4]
  wire  _T_768; // @[execute.scala 79:15:@2208.4]
  wire [6:0] _T_770; // @[execute.scala 79:37:@2209.4]
  wire [6:0] _T_771; // @[execute.scala 79:37:@2210.4]
  wire [5:0] _T_772; // @[execute.scala 79:37:@2211.4]
  wire [6:0] _T_775; // @[execute.scala 79:60:@2212.4]
  wire [5:0] _T_776; // @[execute.scala 79:60:@2213.4]
  wire  _GEN_6529; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6530; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6531; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6532; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6533; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6534; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6535; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6536; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6537; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6538; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6539; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6540; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6541; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6542; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6543; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6544; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6545; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6546; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6547; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6548; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6549; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6550; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6551; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6552; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6553; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6554; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6555; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6556; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6557; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6558; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6559; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6560; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6561; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6562; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6563; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6564; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6565; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6566; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6567; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6568; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6569; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6570; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6571; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6572; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6573; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6574; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6575; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6576; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6577; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6578; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6579; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6580; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6581; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6582; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6583; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6584; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6585; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6586; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6587; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6588; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6589; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6590; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6591; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6593; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6594; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6595; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6596; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6597; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6598; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6599; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6600; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6601; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6602; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6603; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6604; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6605; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6606; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6607; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6608; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6609; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6610; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6611; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6612; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6613; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6614; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6615; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6616; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6617; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6618; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6619; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6620; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6621; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6622; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6623; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6624; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6625; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6626; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6627; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6628; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6629; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6630; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6631; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6632; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6633; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6634; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6635; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6636; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6637; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6638; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6639; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6640; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6641; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6642; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6643; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6644; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6645; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6646; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6647; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6648; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6649; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6650; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6651; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6652; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6653; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6654; // @[execute.scala 79:10:@2214.4]
  wire  _GEN_6655; // @[execute.scala 79:10:@2214.4]
  wire  _T_778; // @[execute.scala 79:10:@2214.4]
  wire  _T_780; // @[execute.scala 79:15:@2215.4]
  wire [6:0] _T_782; // @[execute.scala 79:37:@2216.4]
  wire [6:0] _T_783; // @[execute.scala 79:37:@2217.4]
  wire [5:0] _T_784; // @[execute.scala 79:37:@2218.4]
  wire [6:0] _T_787; // @[execute.scala 79:60:@2219.4]
  wire [5:0] _T_788; // @[execute.scala 79:60:@2220.4]
  wire  _GEN_6657; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6658; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6659; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6660; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6661; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6662; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6663; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6664; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6665; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6666; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6667; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6668; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6669; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6670; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6671; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6672; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6673; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6674; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6675; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6676; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6677; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6678; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6679; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6680; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6681; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6682; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6683; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6684; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6685; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6686; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6687; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6688; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6689; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6690; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6691; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6692; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6693; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6694; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6695; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6696; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6697; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6698; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6699; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6700; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6701; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6702; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6703; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6704; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6705; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6706; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6707; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6708; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6709; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6710; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6711; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6712; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6713; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6714; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6715; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6716; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6717; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6718; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6719; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6721; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6722; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6723; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6724; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6725; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6726; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6727; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6728; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6729; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6730; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6731; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6732; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6733; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6734; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6735; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6736; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6737; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6738; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6739; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6740; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6741; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6742; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6743; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6744; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6745; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6746; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6747; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6748; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6749; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6750; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6751; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6752; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6753; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6754; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6755; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6756; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6757; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6758; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6759; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6760; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6761; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6762; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6763; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6764; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6765; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6766; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6767; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6768; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6769; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6770; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6771; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6772; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6773; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6774; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6775; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6776; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6777; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6778; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6779; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6780; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6781; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6782; // @[execute.scala 79:10:@2221.4]
  wire  _GEN_6783; // @[execute.scala 79:10:@2221.4]
  wire  _T_790; // @[execute.scala 79:10:@2221.4]
  wire  _T_792; // @[execute.scala 79:15:@2222.4]
  wire [6:0] _T_794; // @[execute.scala 79:37:@2223.4]
  wire [6:0] _T_795; // @[execute.scala 79:37:@2224.4]
  wire [5:0] _T_796; // @[execute.scala 79:37:@2225.4]
  wire [6:0] _T_799; // @[execute.scala 79:60:@2226.4]
  wire [5:0] _T_800; // @[execute.scala 79:60:@2227.4]
  wire  _GEN_6785; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6786; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6787; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6788; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6789; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6790; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6791; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6792; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6793; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6794; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6795; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6796; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6797; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6798; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6799; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6800; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6801; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6802; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6803; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6804; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6805; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6806; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6807; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6808; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6809; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6810; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6811; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6812; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6813; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6814; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6815; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6816; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6817; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6818; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6819; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6820; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6821; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6822; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6823; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6824; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6825; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6826; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6827; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6828; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6829; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6830; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6831; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6832; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6833; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6834; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6835; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6836; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6837; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6838; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6839; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6840; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6841; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6842; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6843; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6844; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6845; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6846; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6847; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6849; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6850; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6851; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6852; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6853; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6854; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6855; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6856; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6857; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6858; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6859; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6860; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6861; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6862; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6863; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6864; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6865; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6866; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6867; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6868; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6869; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6870; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6871; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6872; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6873; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6874; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6875; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6876; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6877; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6878; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6879; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6880; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6881; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6882; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6883; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6884; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6885; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6886; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6887; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6888; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6889; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6890; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6891; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6892; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6893; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6894; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6895; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6896; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6897; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6898; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6899; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6900; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6901; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6902; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6903; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6904; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6905; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6906; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6907; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6908; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6909; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6910; // @[execute.scala 79:10:@2228.4]
  wire  _GEN_6911; // @[execute.scala 79:10:@2228.4]
  wire  _T_802; // @[execute.scala 79:10:@2228.4]
  wire  _T_804; // @[execute.scala 79:15:@2229.4]
  wire [6:0] _T_806; // @[execute.scala 79:37:@2230.4]
  wire [6:0] _T_807; // @[execute.scala 79:37:@2231.4]
  wire [5:0] _T_808; // @[execute.scala 79:37:@2232.4]
  wire [6:0] _T_811; // @[execute.scala 79:60:@2233.4]
  wire [5:0] _T_812; // @[execute.scala 79:60:@2234.4]
  wire  _GEN_6913; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6914; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6915; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6916; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6917; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6918; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6919; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6920; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6921; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6922; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6923; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6924; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6925; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6926; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6927; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6928; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6929; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6930; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6931; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6932; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6933; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6934; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6935; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6936; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6937; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6938; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6939; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6940; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6941; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6942; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6943; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6944; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6945; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6946; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6947; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6948; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6949; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6950; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6951; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6952; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6953; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6954; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6955; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6956; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6957; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6958; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6959; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6960; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6961; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6962; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6963; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6964; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6965; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6966; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6967; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6968; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6969; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6970; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6971; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6972; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6973; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6974; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6975; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6977; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6978; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6979; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6980; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6981; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6982; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6983; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6984; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6985; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6986; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6987; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6988; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6989; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6990; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6991; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6992; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6993; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6994; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6995; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6996; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6997; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6998; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_6999; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7000; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7001; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7002; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7003; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7004; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7005; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7006; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7007; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7008; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7009; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7010; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7011; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7012; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7013; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7014; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7015; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7016; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7017; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7018; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7019; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7020; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7021; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7022; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7023; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7024; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7025; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7026; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7027; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7028; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7029; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7030; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7031; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7032; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7033; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7034; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7035; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7036; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7037; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7038; // @[execute.scala 79:10:@2235.4]
  wire  _GEN_7039; // @[execute.scala 79:10:@2235.4]
  wire  _T_814; // @[execute.scala 79:10:@2235.4]
  wire  _T_816; // @[execute.scala 79:15:@2236.4]
  wire [6:0] _T_818; // @[execute.scala 79:37:@2237.4]
  wire [6:0] _T_819; // @[execute.scala 79:37:@2238.4]
  wire [5:0] _T_820; // @[execute.scala 79:37:@2239.4]
  wire [6:0] _T_823; // @[execute.scala 79:60:@2240.4]
  wire [5:0] _T_824; // @[execute.scala 79:60:@2241.4]
  wire  _GEN_7041; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7042; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7043; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7044; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7045; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7046; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7047; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7048; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7049; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7050; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7051; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7052; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7053; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7054; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7055; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7056; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7057; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7058; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7059; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7060; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7061; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7062; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7063; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7064; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7065; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7066; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7067; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7068; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7069; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7070; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7071; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7072; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7073; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7074; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7075; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7076; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7077; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7078; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7079; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7080; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7081; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7082; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7083; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7084; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7085; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7086; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7087; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7088; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7089; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7090; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7091; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7092; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7093; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7094; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7095; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7096; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7097; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7098; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7099; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7100; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7101; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7102; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7103; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7105; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7106; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7107; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7108; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7109; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7110; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7111; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7112; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7113; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7114; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7115; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7116; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7117; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7118; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7119; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7120; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7121; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7122; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7123; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7124; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7125; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7126; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7127; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7128; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7129; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7130; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7131; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7132; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7133; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7134; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7135; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7136; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7137; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7138; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7139; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7140; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7141; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7142; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7143; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7144; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7145; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7146; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7147; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7148; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7149; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7150; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7151; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7152; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7153; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7154; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7155; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7156; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7157; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7158; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7159; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7160; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7161; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7162; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7163; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7164; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7165; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7166; // @[execute.scala 79:10:@2242.4]
  wire  _GEN_7167; // @[execute.scala 79:10:@2242.4]
  wire  _T_826; // @[execute.scala 79:10:@2242.4]
  wire  _T_828; // @[execute.scala 79:15:@2243.4]
  wire [6:0] _T_830; // @[execute.scala 79:37:@2244.4]
  wire [6:0] _T_831; // @[execute.scala 79:37:@2245.4]
  wire [5:0] _T_832; // @[execute.scala 79:37:@2246.4]
  wire [6:0] _T_835; // @[execute.scala 79:60:@2247.4]
  wire [5:0] _T_836; // @[execute.scala 79:60:@2248.4]
  wire  _GEN_7169; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7170; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7171; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7172; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7173; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7174; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7175; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7176; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7177; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7178; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7179; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7180; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7181; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7182; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7183; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7184; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7185; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7186; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7187; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7188; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7189; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7190; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7191; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7192; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7193; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7194; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7195; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7196; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7197; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7198; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7199; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7200; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7201; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7202; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7203; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7204; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7205; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7206; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7207; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7208; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7209; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7210; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7211; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7212; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7213; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7214; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7215; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7216; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7217; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7218; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7219; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7220; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7221; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7222; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7223; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7224; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7225; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7226; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7227; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7228; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7229; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7230; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7231; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7233; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7234; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7235; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7236; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7237; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7238; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7239; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7240; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7241; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7242; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7243; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7244; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7245; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7246; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7247; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7248; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7249; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7250; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7251; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7252; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7253; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7254; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7255; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7256; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7257; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7258; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7259; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7260; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7261; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7262; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7263; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7264; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7265; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7266; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7267; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7268; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7269; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7270; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7271; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7272; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7273; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7274; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7275; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7276; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7277; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7278; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7279; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7280; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7281; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7282; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7283; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7284; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7285; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7286; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7287; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7288; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7289; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7290; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7291; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7292; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7293; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7294; // @[execute.scala 79:10:@2249.4]
  wire  _GEN_7295; // @[execute.scala 79:10:@2249.4]
  wire  _T_838; // @[execute.scala 79:10:@2249.4]
  wire  _T_840; // @[execute.scala 79:15:@2250.4]
  wire [6:0] _T_842; // @[execute.scala 79:37:@2251.4]
  wire [6:0] _T_843; // @[execute.scala 79:37:@2252.4]
  wire [5:0] _T_844; // @[execute.scala 79:37:@2253.4]
  wire [6:0] _T_847; // @[execute.scala 79:60:@2254.4]
  wire [5:0] _T_848; // @[execute.scala 79:60:@2255.4]
  wire  _GEN_7297; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7298; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7299; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7300; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7301; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7302; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7303; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7304; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7305; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7306; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7307; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7308; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7309; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7310; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7311; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7312; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7313; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7314; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7315; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7316; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7317; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7318; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7319; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7320; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7321; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7322; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7323; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7324; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7325; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7326; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7327; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7328; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7329; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7330; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7331; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7332; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7333; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7334; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7335; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7336; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7337; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7338; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7339; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7340; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7341; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7342; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7343; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7344; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7345; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7346; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7347; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7348; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7349; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7350; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7351; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7352; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7353; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7354; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7355; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7356; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7357; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7358; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7359; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7361; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7362; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7363; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7364; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7365; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7366; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7367; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7368; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7369; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7370; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7371; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7372; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7373; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7374; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7375; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7376; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7377; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7378; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7379; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7380; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7381; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7382; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7383; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7384; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7385; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7386; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7387; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7388; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7389; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7390; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7391; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7392; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7393; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7394; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7395; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7396; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7397; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7398; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7399; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7400; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7401; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7402; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7403; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7404; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7405; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7406; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7407; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7408; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7409; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7410; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7411; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7412; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7413; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7414; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7415; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7416; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7417; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7418; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7419; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7420; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7421; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7422; // @[execute.scala 79:10:@2256.4]
  wire  _GEN_7423; // @[execute.scala 79:10:@2256.4]
  wire  _T_850; // @[execute.scala 79:10:@2256.4]
  wire  _T_852; // @[execute.scala 79:15:@2257.4]
  wire [6:0] _T_854; // @[execute.scala 79:37:@2258.4]
  wire [6:0] _T_855; // @[execute.scala 79:37:@2259.4]
  wire [5:0] _T_856; // @[execute.scala 79:37:@2260.4]
  wire [6:0] _T_859; // @[execute.scala 79:60:@2261.4]
  wire [5:0] _T_860; // @[execute.scala 79:60:@2262.4]
  wire  _GEN_7425; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7426; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7427; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7428; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7429; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7430; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7431; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7432; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7433; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7434; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7435; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7436; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7437; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7438; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7439; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7440; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7441; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7442; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7443; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7444; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7445; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7446; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7447; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7448; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7449; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7450; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7451; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7452; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7453; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7454; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7455; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7456; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7457; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7458; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7459; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7460; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7461; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7462; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7463; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7464; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7465; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7466; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7467; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7468; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7469; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7470; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7471; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7472; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7473; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7474; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7475; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7476; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7477; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7478; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7479; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7480; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7481; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7482; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7483; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7484; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7485; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7486; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7487; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7489; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7490; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7491; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7492; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7493; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7494; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7495; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7496; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7497; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7498; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7499; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7500; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7501; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7502; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7503; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7504; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7505; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7506; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7507; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7508; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7509; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7510; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7511; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7512; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7513; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7514; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7515; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7516; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7517; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7518; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7519; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7520; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7521; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7522; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7523; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7524; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7525; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7526; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7527; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7528; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7529; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7530; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7531; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7532; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7533; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7534; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7535; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7536; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7537; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7538; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7539; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7540; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7541; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7542; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7543; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7544; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7545; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7546; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7547; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7548; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7549; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7550; // @[execute.scala 79:10:@2263.4]
  wire  _GEN_7551; // @[execute.scala 79:10:@2263.4]
  wire  _T_862; // @[execute.scala 79:10:@2263.4]
  wire  _T_864; // @[execute.scala 79:15:@2264.4]
  wire [6:0] _T_866; // @[execute.scala 79:37:@2265.4]
  wire [6:0] _T_867; // @[execute.scala 79:37:@2266.4]
  wire [5:0] _T_868; // @[execute.scala 79:37:@2267.4]
  wire [6:0] _T_871; // @[execute.scala 79:60:@2268.4]
  wire [5:0] _T_872; // @[execute.scala 79:60:@2269.4]
  wire  _GEN_7553; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7554; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7555; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7556; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7557; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7558; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7559; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7560; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7561; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7562; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7563; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7564; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7565; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7566; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7567; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7568; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7569; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7570; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7571; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7572; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7573; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7574; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7575; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7576; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7577; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7578; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7579; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7580; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7581; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7582; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7583; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7584; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7585; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7586; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7587; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7588; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7589; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7590; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7591; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7592; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7593; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7594; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7595; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7596; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7597; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7598; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7599; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7600; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7601; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7602; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7603; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7604; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7605; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7606; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7607; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7608; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7609; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7610; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7611; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7612; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7613; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7614; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7615; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7617; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7618; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7619; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7620; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7621; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7622; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7623; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7624; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7625; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7626; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7627; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7628; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7629; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7630; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7631; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7632; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7633; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7634; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7635; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7636; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7637; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7638; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7639; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7640; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7641; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7642; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7643; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7644; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7645; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7646; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7647; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7648; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7649; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7650; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7651; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7652; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7653; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7654; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7655; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7656; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7657; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7658; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7659; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7660; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7661; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7662; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7663; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7664; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7665; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7666; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7667; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7668; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7669; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7670; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7671; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7672; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7673; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7674; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7675; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7676; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7677; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7678; // @[execute.scala 79:10:@2270.4]
  wire  _GEN_7679; // @[execute.scala 79:10:@2270.4]
  wire  _T_874; // @[execute.scala 79:10:@2270.4]
  wire  _T_876; // @[execute.scala 79:15:@2271.4]
  wire [6:0] _T_878; // @[execute.scala 79:37:@2272.4]
  wire [6:0] _T_879; // @[execute.scala 79:37:@2273.4]
  wire [5:0] _T_880; // @[execute.scala 79:37:@2274.4]
  wire [6:0] _T_883; // @[execute.scala 79:60:@2275.4]
  wire [5:0] _T_884; // @[execute.scala 79:60:@2276.4]
  wire  _GEN_7681; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7682; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7683; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7684; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7685; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7686; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7687; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7688; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7689; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7690; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7691; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7692; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7693; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7694; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7695; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7696; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7697; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7698; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7699; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7700; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7701; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7702; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7703; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7704; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7705; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7706; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7707; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7708; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7709; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7710; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7711; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7712; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7713; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7714; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7715; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7716; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7717; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7718; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7719; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7720; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7721; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7722; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7723; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7724; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7725; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7726; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7727; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7728; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7729; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7730; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7731; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7732; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7733; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7734; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7735; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7736; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7737; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7738; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7739; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7740; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7741; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7742; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7743; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7745; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7746; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7747; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7748; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7749; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7750; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7751; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7752; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7753; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7754; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7755; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7756; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7757; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7758; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7759; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7760; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7761; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7762; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7763; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7764; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7765; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7766; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7767; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7768; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7769; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7770; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7771; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7772; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7773; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7774; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7775; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7776; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7777; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7778; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7779; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7780; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7781; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7782; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7783; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7784; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7785; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7786; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7787; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7788; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7789; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7790; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7791; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7792; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7793; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7794; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7795; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7796; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7797; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7798; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7799; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7800; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7801; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7802; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7803; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7804; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7805; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7806; // @[execute.scala 79:10:@2277.4]
  wire  _GEN_7807; // @[execute.scala 79:10:@2277.4]
  wire  _T_886; // @[execute.scala 79:10:@2277.4]
  wire  _T_888; // @[execute.scala 79:15:@2278.4]
  wire [6:0] _T_890; // @[execute.scala 79:37:@2279.4]
  wire [6:0] _T_891; // @[execute.scala 79:37:@2280.4]
  wire [5:0] _T_892; // @[execute.scala 79:37:@2281.4]
  wire [6:0] _T_895; // @[execute.scala 79:60:@2282.4]
  wire [5:0] _T_896; // @[execute.scala 79:60:@2283.4]
  wire  _GEN_7809; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7810; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7811; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7812; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7813; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7814; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7815; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7816; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7817; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7818; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7819; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7820; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7821; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7822; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7823; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7824; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7825; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7826; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7827; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7828; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7829; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7830; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7831; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7832; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7833; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7834; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7835; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7836; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7837; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7838; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7839; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7840; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7841; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7842; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7843; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7844; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7845; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7846; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7847; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7848; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7849; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7850; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7851; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7852; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7853; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7854; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7855; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7856; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7857; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7858; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7859; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7860; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7861; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7862; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7863; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7864; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7865; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7866; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7867; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7868; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7869; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7870; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7871; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7873; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7874; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7875; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7876; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7877; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7878; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7879; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7880; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7881; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7882; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7883; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7884; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7885; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7886; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7887; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7888; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7889; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7890; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7891; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7892; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7893; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7894; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7895; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7896; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7897; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7898; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7899; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7900; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7901; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7902; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7903; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7904; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7905; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7906; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7907; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7908; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7909; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7910; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7911; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7912; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7913; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7914; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7915; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7916; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7917; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7918; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7919; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7920; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7921; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7922; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7923; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7924; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7925; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7926; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7927; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7928; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7929; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7930; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7931; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7932; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7933; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7934; // @[execute.scala 79:10:@2284.4]
  wire  _GEN_7935; // @[execute.scala 79:10:@2284.4]
  wire  _T_898; // @[execute.scala 79:10:@2284.4]
  wire  _T_900; // @[execute.scala 79:15:@2285.4]
  wire [6:0] _T_902; // @[execute.scala 79:37:@2286.4]
  wire [6:0] _T_903; // @[execute.scala 79:37:@2287.4]
  wire [5:0] _T_904; // @[execute.scala 79:37:@2288.4]
  wire [6:0] _T_907; // @[execute.scala 79:60:@2289.4]
  wire [5:0] _T_908; // @[execute.scala 79:60:@2290.4]
  wire  _GEN_7937; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7938; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7939; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7940; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7941; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7942; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7943; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7944; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7945; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7946; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7947; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7948; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7949; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7950; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7951; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7952; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7953; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7954; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7955; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7956; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7957; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7958; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7959; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7960; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7961; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7962; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7963; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7964; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7965; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7966; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7967; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7968; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7969; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7970; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7971; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7972; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7973; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7974; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7975; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7976; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7977; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7978; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7979; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7980; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7981; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7982; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7983; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7984; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7985; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7986; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7987; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7988; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7989; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7990; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7991; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7992; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7993; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7994; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7995; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7996; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7997; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7998; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_7999; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8001; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8002; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8003; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8004; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8005; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8006; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8007; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8008; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8009; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8010; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8011; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8012; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8013; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8014; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8015; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8016; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8017; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8018; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8019; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8020; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8021; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8022; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8023; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8024; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8025; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8026; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8027; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8028; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8029; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8030; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8031; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8032; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8033; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8034; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8035; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8036; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8037; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8038; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8039; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8040; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8041; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8042; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8043; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8044; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8045; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8046; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8047; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8048; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8049; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8050; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8051; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8052; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8053; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8054; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8055; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8056; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8057; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8058; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8059; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8060; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8061; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8062; // @[execute.scala 79:10:@2291.4]
  wire  _GEN_8063; // @[execute.scala 79:10:@2291.4]
  wire  _T_910; // @[execute.scala 79:10:@2291.4]
  wire  _T_912; // @[execute.scala 79:15:@2292.4]
  wire [6:0] _T_914; // @[execute.scala 79:37:@2293.4]
  wire [6:0] _T_915; // @[execute.scala 79:37:@2294.4]
  wire [5:0] _T_916; // @[execute.scala 79:37:@2295.4]
  wire [6:0] _T_919; // @[execute.scala 79:60:@2296.4]
  wire [5:0] _T_920; // @[execute.scala 79:60:@2297.4]
  wire  _GEN_8065; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8066; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8067; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8068; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8069; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8070; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8071; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8072; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8073; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8074; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8075; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8076; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8077; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8078; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8079; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8080; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8081; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8082; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8083; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8084; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8085; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8086; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8087; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8088; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8089; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8090; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8091; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8092; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8093; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8094; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8095; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8096; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8097; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8098; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8099; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8100; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8101; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8102; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8103; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8104; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8105; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8106; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8107; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8108; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8109; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8110; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8111; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8112; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8113; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8114; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8115; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8116; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8117; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8118; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8119; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8120; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8121; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8122; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8123; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8124; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8125; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8126; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8127; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8129; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8130; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8131; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8132; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8133; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8134; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8135; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8136; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8137; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8138; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8139; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8140; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8141; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8142; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8143; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8144; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8145; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8146; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8147; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8148; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8149; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8150; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8151; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8152; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8153; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8154; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8155; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8156; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8157; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8158; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8159; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8160; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8161; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8162; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8163; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8164; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8165; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8166; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8167; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8168; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8169; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8170; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8171; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8172; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8173; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8174; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8175; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8176; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8177; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8178; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8179; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8180; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8181; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8182; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8183; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8184; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8185; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8186; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8187; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8188; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8189; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8190; // @[execute.scala 79:10:@2298.4]
  wire  _GEN_8191; // @[execute.scala 79:10:@2298.4]
  wire  _T_922; // @[execute.scala 79:10:@2298.4]
  wire [7:0] _T_999; // @[execute.scala 89:73:@2370.4]
  wire [15:0] _T_1007; // @[execute.scala 89:73:@2378.4]
  wire [7:0] _T_1014; // @[execute.scala 89:73:@2385.4]
  wire [31:0] _T_1023; // @[execute.scala 89:73:@2394.4]
  wire [7:0] _T_1030; // @[execute.scala 89:73:@2401.4]
  wire [15:0] _T_1038; // @[execute.scala 89:73:@2409.4]
  wire [7:0] _T_1045; // @[execute.scala 89:73:@2416.4]
  wire [31:0] _T_1054; // @[execute.scala 89:73:@2425.4]
  wire [63:0] _T_1055; // @[execute.scala 89:73:@2426.4]
  wire  _T_1056; // @[Mux.scala 46:19:@2427.4]
  wire [63:0] _T_1057; // @[Mux.scala 46:16:@2428.4]
  wire  _T_1058; // @[Mux.scala 46:19:@2429.4]
  wire [63:0] _T_1059; // @[Mux.scala 46:16:@2430.4]
  wire  _T_1060; // @[Mux.scala 46:19:@2431.4]
  wire [63:0] _T_1061; // @[Mux.scala 46:16:@2432.4]
  wire  _T_1062; // @[Mux.scala 46:19:@2433.4]
  wire [126:0] res; // @[Mux.scala 46:16:@2434.4]
  assign _GEN_8192 = {{63'd0}, io_word}; // @[execute.scala 86:33:@1716.4]
  assign _T_15 = _GEN_8192 << io_amount; // @[execute.scala 86:33:@1716.4]
  assign _T_16 = io_word >> io_amount; // @[execute.scala 87:33:@1717.4]
  assign _T_17 = $signed(io_word); // @[execute.scala 88:39:@1718.4]
  assign _T_18 = $signed(_T_17) >>> io_amount; // @[execute.scala 88:42:@1719.4]
  assign _T_19 = $unsigned(_T_18); // @[execute.scala 88:62:@1720.4]
  assign _T_20 = io_word[0]; // @[execute.scala 89:52:@1721.4]
  assign _T_21 = io_word[1]; // @[execute.scala 89:52:@1722.4]
  assign _T_22 = io_word[2]; // @[execute.scala 89:52:@1723.4]
  assign _T_23 = io_word[3]; // @[execute.scala 89:52:@1724.4]
  assign _T_24 = io_word[4]; // @[execute.scala 89:52:@1725.4]
  assign _T_25 = io_word[5]; // @[execute.scala 89:52:@1726.4]
  assign _T_26 = io_word[6]; // @[execute.scala 89:52:@1727.4]
  assign _T_27 = io_word[7]; // @[execute.scala 89:52:@1728.4]
  assign _T_28 = io_word[8]; // @[execute.scala 89:52:@1729.4]
  assign _T_29 = io_word[9]; // @[execute.scala 89:52:@1730.4]
  assign _T_30 = io_word[10]; // @[execute.scala 89:52:@1731.4]
  assign _T_31 = io_word[11]; // @[execute.scala 89:52:@1732.4]
  assign _T_32 = io_word[12]; // @[execute.scala 89:52:@1733.4]
  assign _T_33 = io_word[13]; // @[execute.scala 89:52:@1734.4]
  assign _T_34 = io_word[14]; // @[execute.scala 89:52:@1735.4]
  assign _T_35 = io_word[15]; // @[execute.scala 89:52:@1736.4]
  assign _T_36 = io_word[16]; // @[execute.scala 89:52:@1737.4]
  assign _T_37 = io_word[17]; // @[execute.scala 89:52:@1738.4]
  assign _T_38 = io_word[18]; // @[execute.scala 89:52:@1739.4]
  assign _T_39 = io_word[19]; // @[execute.scala 89:52:@1740.4]
  assign _T_40 = io_word[20]; // @[execute.scala 89:52:@1741.4]
  assign _T_41 = io_word[21]; // @[execute.scala 89:52:@1742.4]
  assign _T_42 = io_word[22]; // @[execute.scala 89:52:@1743.4]
  assign _T_43 = io_word[23]; // @[execute.scala 89:52:@1744.4]
  assign _T_44 = io_word[24]; // @[execute.scala 89:52:@1745.4]
  assign _T_45 = io_word[25]; // @[execute.scala 89:52:@1746.4]
  assign _T_46 = io_word[26]; // @[execute.scala 89:52:@1747.4]
  assign _T_47 = io_word[27]; // @[execute.scala 89:52:@1748.4]
  assign _T_48 = io_word[28]; // @[execute.scala 89:52:@1749.4]
  assign _T_49 = io_word[29]; // @[execute.scala 89:52:@1750.4]
  assign _T_50 = io_word[30]; // @[execute.scala 89:52:@1751.4]
  assign _T_51 = io_word[31]; // @[execute.scala 89:52:@1752.4]
  assign _T_52 = io_word[32]; // @[execute.scala 89:52:@1753.4]
  assign _T_53 = io_word[33]; // @[execute.scala 89:52:@1754.4]
  assign _T_54 = io_word[34]; // @[execute.scala 89:52:@1755.4]
  assign _T_55 = io_word[35]; // @[execute.scala 89:52:@1756.4]
  assign _T_56 = io_word[36]; // @[execute.scala 89:52:@1757.4]
  assign _T_57 = io_word[37]; // @[execute.scala 89:52:@1758.4]
  assign _T_58 = io_word[38]; // @[execute.scala 89:52:@1759.4]
  assign _T_59 = io_word[39]; // @[execute.scala 89:52:@1760.4]
  assign _T_60 = io_word[40]; // @[execute.scala 89:52:@1761.4]
  assign _T_61 = io_word[41]; // @[execute.scala 89:52:@1762.4]
  assign _T_62 = io_word[42]; // @[execute.scala 89:52:@1763.4]
  assign _T_63 = io_word[43]; // @[execute.scala 89:52:@1764.4]
  assign _T_64 = io_word[44]; // @[execute.scala 89:52:@1765.4]
  assign _T_65 = io_word[45]; // @[execute.scala 89:52:@1766.4]
  assign _T_66 = io_word[46]; // @[execute.scala 89:52:@1767.4]
  assign _T_67 = io_word[47]; // @[execute.scala 89:52:@1768.4]
  assign _T_68 = io_word[48]; // @[execute.scala 89:52:@1769.4]
  assign _T_69 = io_word[49]; // @[execute.scala 89:52:@1770.4]
  assign _T_70 = io_word[50]; // @[execute.scala 89:52:@1771.4]
  assign _T_71 = io_word[51]; // @[execute.scala 89:52:@1772.4]
  assign _T_72 = io_word[52]; // @[execute.scala 89:52:@1773.4]
  assign _T_73 = io_word[53]; // @[execute.scala 89:52:@1774.4]
  assign _T_74 = io_word[54]; // @[execute.scala 89:52:@1775.4]
  assign _T_75 = io_word[55]; // @[execute.scala 89:52:@1776.4]
  assign _T_76 = io_word[56]; // @[execute.scala 89:52:@1777.4]
  assign _T_77 = io_word[57]; // @[execute.scala 89:52:@1778.4]
  assign _T_78 = io_word[58]; // @[execute.scala 89:52:@1779.4]
  assign _T_79 = io_word[59]; // @[execute.scala 89:52:@1780.4]
  assign _T_80 = io_word[60]; // @[execute.scala 89:52:@1781.4]
  assign _T_81 = io_word[61]; // @[execute.scala 89:52:@1782.4]
  assign _T_82 = io_word[62]; // @[execute.scala 89:52:@1783.4]
  assign _T_83 = io_word[63]; // @[execute.scala 89:52:@1784.4]
  assign _GEN_8193 = {{1'd0}, io_amount}; // @[execute.scala 79:37:@1851.4]
  assign _T_157 = _GEN_8193 - 7'h40; // @[execute.scala 79:37:@1851.4]
  assign _T_158 = $unsigned(_T_157); // @[execute.scala 79:37:@1852.4]
  assign _T_159 = _T_158[6:0]; // @[execute.scala 79:37:@1853.4]
  assign _T_161 = _T_159[5:0]; // @[:@1854.4]
  assign _GEN_1 = 6'h1 == _T_161 ? _T_21 : _T_20; // @[execute.scala 79:10:@1857.4]
  assign _GEN_2 = 6'h2 == _T_161 ? _T_22 : _GEN_1; // @[execute.scala 79:10:@1857.4]
  assign _GEN_3 = 6'h3 == _T_161 ? _T_23 : _GEN_2; // @[execute.scala 79:10:@1857.4]
  assign _GEN_4 = 6'h4 == _T_161 ? _T_24 : _GEN_3; // @[execute.scala 79:10:@1857.4]
  assign _GEN_5 = 6'h5 == _T_161 ? _T_25 : _GEN_4; // @[execute.scala 79:10:@1857.4]
  assign _GEN_6 = 6'h6 == _T_161 ? _T_26 : _GEN_5; // @[execute.scala 79:10:@1857.4]
  assign _GEN_7 = 6'h7 == _T_161 ? _T_27 : _GEN_6; // @[execute.scala 79:10:@1857.4]
  assign _GEN_8 = 6'h8 == _T_161 ? _T_28 : _GEN_7; // @[execute.scala 79:10:@1857.4]
  assign _GEN_9 = 6'h9 == _T_161 ? _T_29 : _GEN_8; // @[execute.scala 79:10:@1857.4]
  assign _GEN_10 = 6'ha == _T_161 ? _T_30 : _GEN_9; // @[execute.scala 79:10:@1857.4]
  assign _GEN_11 = 6'hb == _T_161 ? _T_31 : _GEN_10; // @[execute.scala 79:10:@1857.4]
  assign _GEN_12 = 6'hc == _T_161 ? _T_32 : _GEN_11; // @[execute.scala 79:10:@1857.4]
  assign _GEN_13 = 6'hd == _T_161 ? _T_33 : _GEN_12; // @[execute.scala 79:10:@1857.4]
  assign _GEN_14 = 6'he == _T_161 ? _T_34 : _GEN_13; // @[execute.scala 79:10:@1857.4]
  assign _GEN_15 = 6'hf == _T_161 ? _T_35 : _GEN_14; // @[execute.scala 79:10:@1857.4]
  assign _GEN_16 = 6'h10 == _T_161 ? _T_36 : _GEN_15; // @[execute.scala 79:10:@1857.4]
  assign _GEN_17 = 6'h11 == _T_161 ? _T_37 : _GEN_16; // @[execute.scala 79:10:@1857.4]
  assign _GEN_18 = 6'h12 == _T_161 ? _T_38 : _GEN_17; // @[execute.scala 79:10:@1857.4]
  assign _GEN_19 = 6'h13 == _T_161 ? _T_39 : _GEN_18; // @[execute.scala 79:10:@1857.4]
  assign _GEN_20 = 6'h14 == _T_161 ? _T_40 : _GEN_19; // @[execute.scala 79:10:@1857.4]
  assign _GEN_21 = 6'h15 == _T_161 ? _T_41 : _GEN_20; // @[execute.scala 79:10:@1857.4]
  assign _GEN_22 = 6'h16 == _T_161 ? _T_42 : _GEN_21; // @[execute.scala 79:10:@1857.4]
  assign _GEN_23 = 6'h17 == _T_161 ? _T_43 : _GEN_22; // @[execute.scala 79:10:@1857.4]
  assign _GEN_24 = 6'h18 == _T_161 ? _T_44 : _GEN_23; // @[execute.scala 79:10:@1857.4]
  assign _GEN_25 = 6'h19 == _T_161 ? _T_45 : _GEN_24; // @[execute.scala 79:10:@1857.4]
  assign _GEN_26 = 6'h1a == _T_161 ? _T_46 : _GEN_25; // @[execute.scala 79:10:@1857.4]
  assign _GEN_27 = 6'h1b == _T_161 ? _T_47 : _GEN_26; // @[execute.scala 79:10:@1857.4]
  assign _GEN_28 = 6'h1c == _T_161 ? _T_48 : _GEN_27; // @[execute.scala 79:10:@1857.4]
  assign _GEN_29 = 6'h1d == _T_161 ? _T_49 : _GEN_28; // @[execute.scala 79:10:@1857.4]
  assign _GEN_30 = 6'h1e == _T_161 ? _T_50 : _GEN_29; // @[execute.scala 79:10:@1857.4]
  assign _GEN_31 = 6'h1f == _T_161 ? _T_51 : _GEN_30; // @[execute.scala 79:10:@1857.4]
  assign _GEN_32 = 6'h20 == _T_161 ? _T_52 : _GEN_31; // @[execute.scala 79:10:@1857.4]
  assign _GEN_33 = 6'h21 == _T_161 ? _T_53 : _GEN_32; // @[execute.scala 79:10:@1857.4]
  assign _GEN_34 = 6'h22 == _T_161 ? _T_54 : _GEN_33; // @[execute.scala 79:10:@1857.4]
  assign _GEN_35 = 6'h23 == _T_161 ? _T_55 : _GEN_34; // @[execute.scala 79:10:@1857.4]
  assign _GEN_36 = 6'h24 == _T_161 ? _T_56 : _GEN_35; // @[execute.scala 79:10:@1857.4]
  assign _GEN_37 = 6'h25 == _T_161 ? _T_57 : _GEN_36; // @[execute.scala 79:10:@1857.4]
  assign _GEN_38 = 6'h26 == _T_161 ? _T_58 : _GEN_37; // @[execute.scala 79:10:@1857.4]
  assign _GEN_39 = 6'h27 == _T_161 ? _T_59 : _GEN_38; // @[execute.scala 79:10:@1857.4]
  assign _GEN_40 = 6'h28 == _T_161 ? _T_60 : _GEN_39; // @[execute.scala 79:10:@1857.4]
  assign _GEN_41 = 6'h29 == _T_161 ? _T_61 : _GEN_40; // @[execute.scala 79:10:@1857.4]
  assign _GEN_42 = 6'h2a == _T_161 ? _T_62 : _GEN_41; // @[execute.scala 79:10:@1857.4]
  assign _GEN_43 = 6'h2b == _T_161 ? _T_63 : _GEN_42; // @[execute.scala 79:10:@1857.4]
  assign _GEN_44 = 6'h2c == _T_161 ? _T_64 : _GEN_43; // @[execute.scala 79:10:@1857.4]
  assign _GEN_45 = 6'h2d == _T_161 ? _T_65 : _GEN_44; // @[execute.scala 79:10:@1857.4]
  assign _GEN_46 = 6'h2e == _T_161 ? _T_66 : _GEN_45; // @[execute.scala 79:10:@1857.4]
  assign _GEN_47 = 6'h2f == _T_161 ? _T_67 : _GEN_46; // @[execute.scala 79:10:@1857.4]
  assign _GEN_48 = 6'h30 == _T_161 ? _T_68 : _GEN_47; // @[execute.scala 79:10:@1857.4]
  assign _GEN_49 = 6'h31 == _T_161 ? _T_69 : _GEN_48; // @[execute.scala 79:10:@1857.4]
  assign _GEN_50 = 6'h32 == _T_161 ? _T_70 : _GEN_49; // @[execute.scala 79:10:@1857.4]
  assign _GEN_51 = 6'h33 == _T_161 ? _T_71 : _GEN_50; // @[execute.scala 79:10:@1857.4]
  assign _GEN_52 = 6'h34 == _T_161 ? _T_72 : _GEN_51; // @[execute.scala 79:10:@1857.4]
  assign _GEN_53 = 6'h35 == _T_161 ? _T_73 : _GEN_52; // @[execute.scala 79:10:@1857.4]
  assign _GEN_54 = 6'h36 == _T_161 ? _T_74 : _GEN_53; // @[execute.scala 79:10:@1857.4]
  assign _GEN_55 = 6'h37 == _T_161 ? _T_75 : _GEN_54; // @[execute.scala 79:10:@1857.4]
  assign _GEN_56 = 6'h38 == _T_161 ? _T_76 : _GEN_55; // @[execute.scala 79:10:@1857.4]
  assign _GEN_57 = 6'h39 == _T_161 ? _T_77 : _GEN_56; // @[execute.scala 79:10:@1857.4]
  assign _GEN_58 = 6'h3a == _T_161 ? _T_78 : _GEN_57; // @[execute.scala 79:10:@1857.4]
  assign _GEN_59 = 6'h3b == _T_161 ? _T_79 : _GEN_58; // @[execute.scala 79:10:@1857.4]
  assign _GEN_60 = 6'h3c == _T_161 ? _T_80 : _GEN_59; // @[execute.scala 79:10:@1857.4]
  assign _GEN_61 = 6'h3d == _T_161 ? _T_81 : _GEN_60; // @[execute.scala 79:10:@1857.4]
  assign _GEN_62 = 6'h3e == _T_161 ? _T_82 : _GEN_61; // @[execute.scala 79:10:@1857.4]
  assign _GEN_63 = 6'h3f == _T_161 ? _T_83 : _GEN_62; // @[execute.scala 79:10:@1857.4]
  assign _T_168 = io_amount < 6'h3f; // @[execute.scala 79:15:@1858.4]
  assign _T_170 = io_amount - 6'h3f; // @[execute.scala 79:37:@1859.4]
  assign _T_171 = $unsigned(_T_170); // @[execute.scala 79:37:@1860.4]
  assign _T_172 = _T_171[5:0]; // @[execute.scala 79:37:@1861.4]
  assign _T_175 = 6'h1 + io_amount; // @[execute.scala 79:60:@1862.4]
  assign _T_176 = 6'h1 + io_amount; // @[execute.scala 79:60:@1863.4]
  assign _GEN_129 = 6'h1 == _T_172 ? _T_21 : _T_20; // @[execute.scala 79:10:@1864.4]
  assign _GEN_130 = 6'h2 == _T_172 ? _T_22 : _GEN_129; // @[execute.scala 79:10:@1864.4]
  assign _GEN_131 = 6'h3 == _T_172 ? _T_23 : _GEN_130; // @[execute.scala 79:10:@1864.4]
  assign _GEN_132 = 6'h4 == _T_172 ? _T_24 : _GEN_131; // @[execute.scala 79:10:@1864.4]
  assign _GEN_133 = 6'h5 == _T_172 ? _T_25 : _GEN_132; // @[execute.scala 79:10:@1864.4]
  assign _GEN_134 = 6'h6 == _T_172 ? _T_26 : _GEN_133; // @[execute.scala 79:10:@1864.4]
  assign _GEN_135 = 6'h7 == _T_172 ? _T_27 : _GEN_134; // @[execute.scala 79:10:@1864.4]
  assign _GEN_136 = 6'h8 == _T_172 ? _T_28 : _GEN_135; // @[execute.scala 79:10:@1864.4]
  assign _GEN_137 = 6'h9 == _T_172 ? _T_29 : _GEN_136; // @[execute.scala 79:10:@1864.4]
  assign _GEN_138 = 6'ha == _T_172 ? _T_30 : _GEN_137; // @[execute.scala 79:10:@1864.4]
  assign _GEN_139 = 6'hb == _T_172 ? _T_31 : _GEN_138; // @[execute.scala 79:10:@1864.4]
  assign _GEN_140 = 6'hc == _T_172 ? _T_32 : _GEN_139; // @[execute.scala 79:10:@1864.4]
  assign _GEN_141 = 6'hd == _T_172 ? _T_33 : _GEN_140; // @[execute.scala 79:10:@1864.4]
  assign _GEN_142 = 6'he == _T_172 ? _T_34 : _GEN_141; // @[execute.scala 79:10:@1864.4]
  assign _GEN_143 = 6'hf == _T_172 ? _T_35 : _GEN_142; // @[execute.scala 79:10:@1864.4]
  assign _GEN_144 = 6'h10 == _T_172 ? _T_36 : _GEN_143; // @[execute.scala 79:10:@1864.4]
  assign _GEN_145 = 6'h11 == _T_172 ? _T_37 : _GEN_144; // @[execute.scala 79:10:@1864.4]
  assign _GEN_146 = 6'h12 == _T_172 ? _T_38 : _GEN_145; // @[execute.scala 79:10:@1864.4]
  assign _GEN_147 = 6'h13 == _T_172 ? _T_39 : _GEN_146; // @[execute.scala 79:10:@1864.4]
  assign _GEN_148 = 6'h14 == _T_172 ? _T_40 : _GEN_147; // @[execute.scala 79:10:@1864.4]
  assign _GEN_149 = 6'h15 == _T_172 ? _T_41 : _GEN_148; // @[execute.scala 79:10:@1864.4]
  assign _GEN_150 = 6'h16 == _T_172 ? _T_42 : _GEN_149; // @[execute.scala 79:10:@1864.4]
  assign _GEN_151 = 6'h17 == _T_172 ? _T_43 : _GEN_150; // @[execute.scala 79:10:@1864.4]
  assign _GEN_152 = 6'h18 == _T_172 ? _T_44 : _GEN_151; // @[execute.scala 79:10:@1864.4]
  assign _GEN_153 = 6'h19 == _T_172 ? _T_45 : _GEN_152; // @[execute.scala 79:10:@1864.4]
  assign _GEN_154 = 6'h1a == _T_172 ? _T_46 : _GEN_153; // @[execute.scala 79:10:@1864.4]
  assign _GEN_155 = 6'h1b == _T_172 ? _T_47 : _GEN_154; // @[execute.scala 79:10:@1864.4]
  assign _GEN_156 = 6'h1c == _T_172 ? _T_48 : _GEN_155; // @[execute.scala 79:10:@1864.4]
  assign _GEN_157 = 6'h1d == _T_172 ? _T_49 : _GEN_156; // @[execute.scala 79:10:@1864.4]
  assign _GEN_158 = 6'h1e == _T_172 ? _T_50 : _GEN_157; // @[execute.scala 79:10:@1864.4]
  assign _GEN_159 = 6'h1f == _T_172 ? _T_51 : _GEN_158; // @[execute.scala 79:10:@1864.4]
  assign _GEN_160 = 6'h20 == _T_172 ? _T_52 : _GEN_159; // @[execute.scala 79:10:@1864.4]
  assign _GEN_161 = 6'h21 == _T_172 ? _T_53 : _GEN_160; // @[execute.scala 79:10:@1864.4]
  assign _GEN_162 = 6'h22 == _T_172 ? _T_54 : _GEN_161; // @[execute.scala 79:10:@1864.4]
  assign _GEN_163 = 6'h23 == _T_172 ? _T_55 : _GEN_162; // @[execute.scala 79:10:@1864.4]
  assign _GEN_164 = 6'h24 == _T_172 ? _T_56 : _GEN_163; // @[execute.scala 79:10:@1864.4]
  assign _GEN_165 = 6'h25 == _T_172 ? _T_57 : _GEN_164; // @[execute.scala 79:10:@1864.4]
  assign _GEN_166 = 6'h26 == _T_172 ? _T_58 : _GEN_165; // @[execute.scala 79:10:@1864.4]
  assign _GEN_167 = 6'h27 == _T_172 ? _T_59 : _GEN_166; // @[execute.scala 79:10:@1864.4]
  assign _GEN_168 = 6'h28 == _T_172 ? _T_60 : _GEN_167; // @[execute.scala 79:10:@1864.4]
  assign _GEN_169 = 6'h29 == _T_172 ? _T_61 : _GEN_168; // @[execute.scala 79:10:@1864.4]
  assign _GEN_170 = 6'h2a == _T_172 ? _T_62 : _GEN_169; // @[execute.scala 79:10:@1864.4]
  assign _GEN_171 = 6'h2b == _T_172 ? _T_63 : _GEN_170; // @[execute.scala 79:10:@1864.4]
  assign _GEN_172 = 6'h2c == _T_172 ? _T_64 : _GEN_171; // @[execute.scala 79:10:@1864.4]
  assign _GEN_173 = 6'h2d == _T_172 ? _T_65 : _GEN_172; // @[execute.scala 79:10:@1864.4]
  assign _GEN_174 = 6'h2e == _T_172 ? _T_66 : _GEN_173; // @[execute.scala 79:10:@1864.4]
  assign _GEN_175 = 6'h2f == _T_172 ? _T_67 : _GEN_174; // @[execute.scala 79:10:@1864.4]
  assign _GEN_176 = 6'h30 == _T_172 ? _T_68 : _GEN_175; // @[execute.scala 79:10:@1864.4]
  assign _GEN_177 = 6'h31 == _T_172 ? _T_69 : _GEN_176; // @[execute.scala 79:10:@1864.4]
  assign _GEN_178 = 6'h32 == _T_172 ? _T_70 : _GEN_177; // @[execute.scala 79:10:@1864.4]
  assign _GEN_179 = 6'h33 == _T_172 ? _T_71 : _GEN_178; // @[execute.scala 79:10:@1864.4]
  assign _GEN_180 = 6'h34 == _T_172 ? _T_72 : _GEN_179; // @[execute.scala 79:10:@1864.4]
  assign _GEN_181 = 6'h35 == _T_172 ? _T_73 : _GEN_180; // @[execute.scala 79:10:@1864.4]
  assign _GEN_182 = 6'h36 == _T_172 ? _T_74 : _GEN_181; // @[execute.scala 79:10:@1864.4]
  assign _GEN_183 = 6'h37 == _T_172 ? _T_75 : _GEN_182; // @[execute.scala 79:10:@1864.4]
  assign _GEN_184 = 6'h38 == _T_172 ? _T_76 : _GEN_183; // @[execute.scala 79:10:@1864.4]
  assign _GEN_185 = 6'h39 == _T_172 ? _T_77 : _GEN_184; // @[execute.scala 79:10:@1864.4]
  assign _GEN_186 = 6'h3a == _T_172 ? _T_78 : _GEN_185; // @[execute.scala 79:10:@1864.4]
  assign _GEN_187 = 6'h3b == _T_172 ? _T_79 : _GEN_186; // @[execute.scala 79:10:@1864.4]
  assign _GEN_188 = 6'h3c == _T_172 ? _T_80 : _GEN_187; // @[execute.scala 79:10:@1864.4]
  assign _GEN_189 = 6'h3d == _T_172 ? _T_81 : _GEN_188; // @[execute.scala 79:10:@1864.4]
  assign _GEN_190 = 6'h3e == _T_172 ? _T_82 : _GEN_189; // @[execute.scala 79:10:@1864.4]
  assign _GEN_191 = 6'h3f == _T_172 ? _T_83 : _GEN_190; // @[execute.scala 79:10:@1864.4]
  assign _GEN_193 = 6'h1 == _T_176 ? _T_21 : _T_20; // @[execute.scala 79:10:@1864.4]
  assign _GEN_194 = 6'h2 == _T_176 ? _T_22 : _GEN_193; // @[execute.scala 79:10:@1864.4]
  assign _GEN_195 = 6'h3 == _T_176 ? _T_23 : _GEN_194; // @[execute.scala 79:10:@1864.4]
  assign _GEN_196 = 6'h4 == _T_176 ? _T_24 : _GEN_195; // @[execute.scala 79:10:@1864.4]
  assign _GEN_197 = 6'h5 == _T_176 ? _T_25 : _GEN_196; // @[execute.scala 79:10:@1864.4]
  assign _GEN_198 = 6'h6 == _T_176 ? _T_26 : _GEN_197; // @[execute.scala 79:10:@1864.4]
  assign _GEN_199 = 6'h7 == _T_176 ? _T_27 : _GEN_198; // @[execute.scala 79:10:@1864.4]
  assign _GEN_200 = 6'h8 == _T_176 ? _T_28 : _GEN_199; // @[execute.scala 79:10:@1864.4]
  assign _GEN_201 = 6'h9 == _T_176 ? _T_29 : _GEN_200; // @[execute.scala 79:10:@1864.4]
  assign _GEN_202 = 6'ha == _T_176 ? _T_30 : _GEN_201; // @[execute.scala 79:10:@1864.4]
  assign _GEN_203 = 6'hb == _T_176 ? _T_31 : _GEN_202; // @[execute.scala 79:10:@1864.4]
  assign _GEN_204 = 6'hc == _T_176 ? _T_32 : _GEN_203; // @[execute.scala 79:10:@1864.4]
  assign _GEN_205 = 6'hd == _T_176 ? _T_33 : _GEN_204; // @[execute.scala 79:10:@1864.4]
  assign _GEN_206 = 6'he == _T_176 ? _T_34 : _GEN_205; // @[execute.scala 79:10:@1864.4]
  assign _GEN_207 = 6'hf == _T_176 ? _T_35 : _GEN_206; // @[execute.scala 79:10:@1864.4]
  assign _GEN_208 = 6'h10 == _T_176 ? _T_36 : _GEN_207; // @[execute.scala 79:10:@1864.4]
  assign _GEN_209 = 6'h11 == _T_176 ? _T_37 : _GEN_208; // @[execute.scala 79:10:@1864.4]
  assign _GEN_210 = 6'h12 == _T_176 ? _T_38 : _GEN_209; // @[execute.scala 79:10:@1864.4]
  assign _GEN_211 = 6'h13 == _T_176 ? _T_39 : _GEN_210; // @[execute.scala 79:10:@1864.4]
  assign _GEN_212 = 6'h14 == _T_176 ? _T_40 : _GEN_211; // @[execute.scala 79:10:@1864.4]
  assign _GEN_213 = 6'h15 == _T_176 ? _T_41 : _GEN_212; // @[execute.scala 79:10:@1864.4]
  assign _GEN_214 = 6'h16 == _T_176 ? _T_42 : _GEN_213; // @[execute.scala 79:10:@1864.4]
  assign _GEN_215 = 6'h17 == _T_176 ? _T_43 : _GEN_214; // @[execute.scala 79:10:@1864.4]
  assign _GEN_216 = 6'h18 == _T_176 ? _T_44 : _GEN_215; // @[execute.scala 79:10:@1864.4]
  assign _GEN_217 = 6'h19 == _T_176 ? _T_45 : _GEN_216; // @[execute.scala 79:10:@1864.4]
  assign _GEN_218 = 6'h1a == _T_176 ? _T_46 : _GEN_217; // @[execute.scala 79:10:@1864.4]
  assign _GEN_219 = 6'h1b == _T_176 ? _T_47 : _GEN_218; // @[execute.scala 79:10:@1864.4]
  assign _GEN_220 = 6'h1c == _T_176 ? _T_48 : _GEN_219; // @[execute.scala 79:10:@1864.4]
  assign _GEN_221 = 6'h1d == _T_176 ? _T_49 : _GEN_220; // @[execute.scala 79:10:@1864.4]
  assign _GEN_222 = 6'h1e == _T_176 ? _T_50 : _GEN_221; // @[execute.scala 79:10:@1864.4]
  assign _GEN_223 = 6'h1f == _T_176 ? _T_51 : _GEN_222; // @[execute.scala 79:10:@1864.4]
  assign _GEN_224 = 6'h20 == _T_176 ? _T_52 : _GEN_223; // @[execute.scala 79:10:@1864.4]
  assign _GEN_225 = 6'h21 == _T_176 ? _T_53 : _GEN_224; // @[execute.scala 79:10:@1864.4]
  assign _GEN_226 = 6'h22 == _T_176 ? _T_54 : _GEN_225; // @[execute.scala 79:10:@1864.4]
  assign _GEN_227 = 6'h23 == _T_176 ? _T_55 : _GEN_226; // @[execute.scala 79:10:@1864.4]
  assign _GEN_228 = 6'h24 == _T_176 ? _T_56 : _GEN_227; // @[execute.scala 79:10:@1864.4]
  assign _GEN_229 = 6'h25 == _T_176 ? _T_57 : _GEN_228; // @[execute.scala 79:10:@1864.4]
  assign _GEN_230 = 6'h26 == _T_176 ? _T_58 : _GEN_229; // @[execute.scala 79:10:@1864.4]
  assign _GEN_231 = 6'h27 == _T_176 ? _T_59 : _GEN_230; // @[execute.scala 79:10:@1864.4]
  assign _GEN_232 = 6'h28 == _T_176 ? _T_60 : _GEN_231; // @[execute.scala 79:10:@1864.4]
  assign _GEN_233 = 6'h29 == _T_176 ? _T_61 : _GEN_232; // @[execute.scala 79:10:@1864.4]
  assign _GEN_234 = 6'h2a == _T_176 ? _T_62 : _GEN_233; // @[execute.scala 79:10:@1864.4]
  assign _GEN_235 = 6'h2b == _T_176 ? _T_63 : _GEN_234; // @[execute.scala 79:10:@1864.4]
  assign _GEN_236 = 6'h2c == _T_176 ? _T_64 : _GEN_235; // @[execute.scala 79:10:@1864.4]
  assign _GEN_237 = 6'h2d == _T_176 ? _T_65 : _GEN_236; // @[execute.scala 79:10:@1864.4]
  assign _GEN_238 = 6'h2e == _T_176 ? _T_66 : _GEN_237; // @[execute.scala 79:10:@1864.4]
  assign _GEN_239 = 6'h2f == _T_176 ? _T_67 : _GEN_238; // @[execute.scala 79:10:@1864.4]
  assign _GEN_240 = 6'h30 == _T_176 ? _T_68 : _GEN_239; // @[execute.scala 79:10:@1864.4]
  assign _GEN_241 = 6'h31 == _T_176 ? _T_69 : _GEN_240; // @[execute.scala 79:10:@1864.4]
  assign _GEN_242 = 6'h32 == _T_176 ? _T_70 : _GEN_241; // @[execute.scala 79:10:@1864.4]
  assign _GEN_243 = 6'h33 == _T_176 ? _T_71 : _GEN_242; // @[execute.scala 79:10:@1864.4]
  assign _GEN_244 = 6'h34 == _T_176 ? _T_72 : _GEN_243; // @[execute.scala 79:10:@1864.4]
  assign _GEN_245 = 6'h35 == _T_176 ? _T_73 : _GEN_244; // @[execute.scala 79:10:@1864.4]
  assign _GEN_246 = 6'h36 == _T_176 ? _T_74 : _GEN_245; // @[execute.scala 79:10:@1864.4]
  assign _GEN_247 = 6'h37 == _T_176 ? _T_75 : _GEN_246; // @[execute.scala 79:10:@1864.4]
  assign _GEN_248 = 6'h38 == _T_176 ? _T_76 : _GEN_247; // @[execute.scala 79:10:@1864.4]
  assign _GEN_249 = 6'h39 == _T_176 ? _T_77 : _GEN_248; // @[execute.scala 79:10:@1864.4]
  assign _GEN_250 = 6'h3a == _T_176 ? _T_78 : _GEN_249; // @[execute.scala 79:10:@1864.4]
  assign _GEN_251 = 6'h3b == _T_176 ? _T_79 : _GEN_250; // @[execute.scala 79:10:@1864.4]
  assign _GEN_252 = 6'h3c == _T_176 ? _T_80 : _GEN_251; // @[execute.scala 79:10:@1864.4]
  assign _GEN_253 = 6'h3d == _T_176 ? _T_81 : _GEN_252; // @[execute.scala 79:10:@1864.4]
  assign _GEN_254 = 6'h3e == _T_176 ? _T_82 : _GEN_253; // @[execute.scala 79:10:@1864.4]
  assign _GEN_255 = 6'h3f == _T_176 ? _T_83 : _GEN_254; // @[execute.scala 79:10:@1864.4]
  assign _T_178 = _T_168 ? _GEN_191 : _GEN_255; // @[execute.scala 79:10:@1864.4]
  assign _T_180 = io_amount < 6'h3e; // @[execute.scala 79:15:@1865.4]
  assign _T_182 = io_amount - 6'h3e; // @[execute.scala 79:37:@1866.4]
  assign _T_183 = $unsigned(_T_182); // @[execute.scala 79:37:@1867.4]
  assign _T_184 = _T_183[5:0]; // @[execute.scala 79:37:@1868.4]
  assign _T_187 = 6'h2 + io_amount; // @[execute.scala 79:60:@1869.4]
  assign _T_188 = 6'h2 + io_amount; // @[execute.scala 79:60:@1870.4]
  assign _GEN_257 = 6'h1 == _T_184 ? _T_21 : _T_20; // @[execute.scala 79:10:@1871.4]
  assign _GEN_258 = 6'h2 == _T_184 ? _T_22 : _GEN_257; // @[execute.scala 79:10:@1871.4]
  assign _GEN_259 = 6'h3 == _T_184 ? _T_23 : _GEN_258; // @[execute.scala 79:10:@1871.4]
  assign _GEN_260 = 6'h4 == _T_184 ? _T_24 : _GEN_259; // @[execute.scala 79:10:@1871.4]
  assign _GEN_261 = 6'h5 == _T_184 ? _T_25 : _GEN_260; // @[execute.scala 79:10:@1871.4]
  assign _GEN_262 = 6'h6 == _T_184 ? _T_26 : _GEN_261; // @[execute.scala 79:10:@1871.4]
  assign _GEN_263 = 6'h7 == _T_184 ? _T_27 : _GEN_262; // @[execute.scala 79:10:@1871.4]
  assign _GEN_264 = 6'h8 == _T_184 ? _T_28 : _GEN_263; // @[execute.scala 79:10:@1871.4]
  assign _GEN_265 = 6'h9 == _T_184 ? _T_29 : _GEN_264; // @[execute.scala 79:10:@1871.4]
  assign _GEN_266 = 6'ha == _T_184 ? _T_30 : _GEN_265; // @[execute.scala 79:10:@1871.4]
  assign _GEN_267 = 6'hb == _T_184 ? _T_31 : _GEN_266; // @[execute.scala 79:10:@1871.4]
  assign _GEN_268 = 6'hc == _T_184 ? _T_32 : _GEN_267; // @[execute.scala 79:10:@1871.4]
  assign _GEN_269 = 6'hd == _T_184 ? _T_33 : _GEN_268; // @[execute.scala 79:10:@1871.4]
  assign _GEN_270 = 6'he == _T_184 ? _T_34 : _GEN_269; // @[execute.scala 79:10:@1871.4]
  assign _GEN_271 = 6'hf == _T_184 ? _T_35 : _GEN_270; // @[execute.scala 79:10:@1871.4]
  assign _GEN_272 = 6'h10 == _T_184 ? _T_36 : _GEN_271; // @[execute.scala 79:10:@1871.4]
  assign _GEN_273 = 6'h11 == _T_184 ? _T_37 : _GEN_272; // @[execute.scala 79:10:@1871.4]
  assign _GEN_274 = 6'h12 == _T_184 ? _T_38 : _GEN_273; // @[execute.scala 79:10:@1871.4]
  assign _GEN_275 = 6'h13 == _T_184 ? _T_39 : _GEN_274; // @[execute.scala 79:10:@1871.4]
  assign _GEN_276 = 6'h14 == _T_184 ? _T_40 : _GEN_275; // @[execute.scala 79:10:@1871.4]
  assign _GEN_277 = 6'h15 == _T_184 ? _T_41 : _GEN_276; // @[execute.scala 79:10:@1871.4]
  assign _GEN_278 = 6'h16 == _T_184 ? _T_42 : _GEN_277; // @[execute.scala 79:10:@1871.4]
  assign _GEN_279 = 6'h17 == _T_184 ? _T_43 : _GEN_278; // @[execute.scala 79:10:@1871.4]
  assign _GEN_280 = 6'h18 == _T_184 ? _T_44 : _GEN_279; // @[execute.scala 79:10:@1871.4]
  assign _GEN_281 = 6'h19 == _T_184 ? _T_45 : _GEN_280; // @[execute.scala 79:10:@1871.4]
  assign _GEN_282 = 6'h1a == _T_184 ? _T_46 : _GEN_281; // @[execute.scala 79:10:@1871.4]
  assign _GEN_283 = 6'h1b == _T_184 ? _T_47 : _GEN_282; // @[execute.scala 79:10:@1871.4]
  assign _GEN_284 = 6'h1c == _T_184 ? _T_48 : _GEN_283; // @[execute.scala 79:10:@1871.4]
  assign _GEN_285 = 6'h1d == _T_184 ? _T_49 : _GEN_284; // @[execute.scala 79:10:@1871.4]
  assign _GEN_286 = 6'h1e == _T_184 ? _T_50 : _GEN_285; // @[execute.scala 79:10:@1871.4]
  assign _GEN_287 = 6'h1f == _T_184 ? _T_51 : _GEN_286; // @[execute.scala 79:10:@1871.4]
  assign _GEN_288 = 6'h20 == _T_184 ? _T_52 : _GEN_287; // @[execute.scala 79:10:@1871.4]
  assign _GEN_289 = 6'h21 == _T_184 ? _T_53 : _GEN_288; // @[execute.scala 79:10:@1871.4]
  assign _GEN_290 = 6'h22 == _T_184 ? _T_54 : _GEN_289; // @[execute.scala 79:10:@1871.4]
  assign _GEN_291 = 6'h23 == _T_184 ? _T_55 : _GEN_290; // @[execute.scala 79:10:@1871.4]
  assign _GEN_292 = 6'h24 == _T_184 ? _T_56 : _GEN_291; // @[execute.scala 79:10:@1871.4]
  assign _GEN_293 = 6'h25 == _T_184 ? _T_57 : _GEN_292; // @[execute.scala 79:10:@1871.4]
  assign _GEN_294 = 6'h26 == _T_184 ? _T_58 : _GEN_293; // @[execute.scala 79:10:@1871.4]
  assign _GEN_295 = 6'h27 == _T_184 ? _T_59 : _GEN_294; // @[execute.scala 79:10:@1871.4]
  assign _GEN_296 = 6'h28 == _T_184 ? _T_60 : _GEN_295; // @[execute.scala 79:10:@1871.4]
  assign _GEN_297 = 6'h29 == _T_184 ? _T_61 : _GEN_296; // @[execute.scala 79:10:@1871.4]
  assign _GEN_298 = 6'h2a == _T_184 ? _T_62 : _GEN_297; // @[execute.scala 79:10:@1871.4]
  assign _GEN_299 = 6'h2b == _T_184 ? _T_63 : _GEN_298; // @[execute.scala 79:10:@1871.4]
  assign _GEN_300 = 6'h2c == _T_184 ? _T_64 : _GEN_299; // @[execute.scala 79:10:@1871.4]
  assign _GEN_301 = 6'h2d == _T_184 ? _T_65 : _GEN_300; // @[execute.scala 79:10:@1871.4]
  assign _GEN_302 = 6'h2e == _T_184 ? _T_66 : _GEN_301; // @[execute.scala 79:10:@1871.4]
  assign _GEN_303 = 6'h2f == _T_184 ? _T_67 : _GEN_302; // @[execute.scala 79:10:@1871.4]
  assign _GEN_304 = 6'h30 == _T_184 ? _T_68 : _GEN_303; // @[execute.scala 79:10:@1871.4]
  assign _GEN_305 = 6'h31 == _T_184 ? _T_69 : _GEN_304; // @[execute.scala 79:10:@1871.4]
  assign _GEN_306 = 6'h32 == _T_184 ? _T_70 : _GEN_305; // @[execute.scala 79:10:@1871.4]
  assign _GEN_307 = 6'h33 == _T_184 ? _T_71 : _GEN_306; // @[execute.scala 79:10:@1871.4]
  assign _GEN_308 = 6'h34 == _T_184 ? _T_72 : _GEN_307; // @[execute.scala 79:10:@1871.4]
  assign _GEN_309 = 6'h35 == _T_184 ? _T_73 : _GEN_308; // @[execute.scala 79:10:@1871.4]
  assign _GEN_310 = 6'h36 == _T_184 ? _T_74 : _GEN_309; // @[execute.scala 79:10:@1871.4]
  assign _GEN_311 = 6'h37 == _T_184 ? _T_75 : _GEN_310; // @[execute.scala 79:10:@1871.4]
  assign _GEN_312 = 6'h38 == _T_184 ? _T_76 : _GEN_311; // @[execute.scala 79:10:@1871.4]
  assign _GEN_313 = 6'h39 == _T_184 ? _T_77 : _GEN_312; // @[execute.scala 79:10:@1871.4]
  assign _GEN_314 = 6'h3a == _T_184 ? _T_78 : _GEN_313; // @[execute.scala 79:10:@1871.4]
  assign _GEN_315 = 6'h3b == _T_184 ? _T_79 : _GEN_314; // @[execute.scala 79:10:@1871.4]
  assign _GEN_316 = 6'h3c == _T_184 ? _T_80 : _GEN_315; // @[execute.scala 79:10:@1871.4]
  assign _GEN_317 = 6'h3d == _T_184 ? _T_81 : _GEN_316; // @[execute.scala 79:10:@1871.4]
  assign _GEN_318 = 6'h3e == _T_184 ? _T_82 : _GEN_317; // @[execute.scala 79:10:@1871.4]
  assign _GEN_319 = 6'h3f == _T_184 ? _T_83 : _GEN_318; // @[execute.scala 79:10:@1871.4]
  assign _GEN_321 = 6'h1 == _T_188 ? _T_21 : _T_20; // @[execute.scala 79:10:@1871.4]
  assign _GEN_322 = 6'h2 == _T_188 ? _T_22 : _GEN_321; // @[execute.scala 79:10:@1871.4]
  assign _GEN_323 = 6'h3 == _T_188 ? _T_23 : _GEN_322; // @[execute.scala 79:10:@1871.4]
  assign _GEN_324 = 6'h4 == _T_188 ? _T_24 : _GEN_323; // @[execute.scala 79:10:@1871.4]
  assign _GEN_325 = 6'h5 == _T_188 ? _T_25 : _GEN_324; // @[execute.scala 79:10:@1871.4]
  assign _GEN_326 = 6'h6 == _T_188 ? _T_26 : _GEN_325; // @[execute.scala 79:10:@1871.4]
  assign _GEN_327 = 6'h7 == _T_188 ? _T_27 : _GEN_326; // @[execute.scala 79:10:@1871.4]
  assign _GEN_328 = 6'h8 == _T_188 ? _T_28 : _GEN_327; // @[execute.scala 79:10:@1871.4]
  assign _GEN_329 = 6'h9 == _T_188 ? _T_29 : _GEN_328; // @[execute.scala 79:10:@1871.4]
  assign _GEN_330 = 6'ha == _T_188 ? _T_30 : _GEN_329; // @[execute.scala 79:10:@1871.4]
  assign _GEN_331 = 6'hb == _T_188 ? _T_31 : _GEN_330; // @[execute.scala 79:10:@1871.4]
  assign _GEN_332 = 6'hc == _T_188 ? _T_32 : _GEN_331; // @[execute.scala 79:10:@1871.4]
  assign _GEN_333 = 6'hd == _T_188 ? _T_33 : _GEN_332; // @[execute.scala 79:10:@1871.4]
  assign _GEN_334 = 6'he == _T_188 ? _T_34 : _GEN_333; // @[execute.scala 79:10:@1871.4]
  assign _GEN_335 = 6'hf == _T_188 ? _T_35 : _GEN_334; // @[execute.scala 79:10:@1871.4]
  assign _GEN_336 = 6'h10 == _T_188 ? _T_36 : _GEN_335; // @[execute.scala 79:10:@1871.4]
  assign _GEN_337 = 6'h11 == _T_188 ? _T_37 : _GEN_336; // @[execute.scala 79:10:@1871.4]
  assign _GEN_338 = 6'h12 == _T_188 ? _T_38 : _GEN_337; // @[execute.scala 79:10:@1871.4]
  assign _GEN_339 = 6'h13 == _T_188 ? _T_39 : _GEN_338; // @[execute.scala 79:10:@1871.4]
  assign _GEN_340 = 6'h14 == _T_188 ? _T_40 : _GEN_339; // @[execute.scala 79:10:@1871.4]
  assign _GEN_341 = 6'h15 == _T_188 ? _T_41 : _GEN_340; // @[execute.scala 79:10:@1871.4]
  assign _GEN_342 = 6'h16 == _T_188 ? _T_42 : _GEN_341; // @[execute.scala 79:10:@1871.4]
  assign _GEN_343 = 6'h17 == _T_188 ? _T_43 : _GEN_342; // @[execute.scala 79:10:@1871.4]
  assign _GEN_344 = 6'h18 == _T_188 ? _T_44 : _GEN_343; // @[execute.scala 79:10:@1871.4]
  assign _GEN_345 = 6'h19 == _T_188 ? _T_45 : _GEN_344; // @[execute.scala 79:10:@1871.4]
  assign _GEN_346 = 6'h1a == _T_188 ? _T_46 : _GEN_345; // @[execute.scala 79:10:@1871.4]
  assign _GEN_347 = 6'h1b == _T_188 ? _T_47 : _GEN_346; // @[execute.scala 79:10:@1871.4]
  assign _GEN_348 = 6'h1c == _T_188 ? _T_48 : _GEN_347; // @[execute.scala 79:10:@1871.4]
  assign _GEN_349 = 6'h1d == _T_188 ? _T_49 : _GEN_348; // @[execute.scala 79:10:@1871.4]
  assign _GEN_350 = 6'h1e == _T_188 ? _T_50 : _GEN_349; // @[execute.scala 79:10:@1871.4]
  assign _GEN_351 = 6'h1f == _T_188 ? _T_51 : _GEN_350; // @[execute.scala 79:10:@1871.4]
  assign _GEN_352 = 6'h20 == _T_188 ? _T_52 : _GEN_351; // @[execute.scala 79:10:@1871.4]
  assign _GEN_353 = 6'h21 == _T_188 ? _T_53 : _GEN_352; // @[execute.scala 79:10:@1871.4]
  assign _GEN_354 = 6'h22 == _T_188 ? _T_54 : _GEN_353; // @[execute.scala 79:10:@1871.4]
  assign _GEN_355 = 6'h23 == _T_188 ? _T_55 : _GEN_354; // @[execute.scala 79:10:@1871.4]
  assign _GEN_356 = 6'h24 == _T_188 ? _T_56 : _GEN_355; // @[execute.scala 79:10:@1871.4]
  assign _GEN_357 = 6'h25 == _T_188 ? _T_57 : _GEN_356; // @[execute.scala 79:10:@1871.4]
  assign _GEN_358 = 6'h26 == _T_188 ? _T_58 : _GEN_357; // @[execute.scala 79:10:@1871.4]
  assign _GEN_359 = 6'h27 == _T_188 ? _T_59 : _GEN_358; // @[execute.scala 79:10:@1871.4]
  assign _GEN_360 = 6'h28 == _T_188 ? _T_60 : _GEN_359; // @[execute.scala 79:10:@1871.4]
  assign _GEN_361 = 6'h29 == _T_188 ? _T_61 : _GEN_360; // @[execute.scala 79:10:@1871.4]
  assign _GEN_362 = 6'h2a == _T_188 ? _T_62 : _GEN_361; // @[execute.scala 79:10:@1871.4]
  assign _GEN_363 = 6'h2b == _T_188 ? _T_63 : _GEN_362; // @[execute.scala 79:10:@1871.4]
  assign _GEN_364 = 6'h2c == _T_188 ? _T_64 : _GEN_363; // @[execute.scala 79:10:@1871.4]
  assign _GEN_365 = 6'h2d == _T_188 ? _T_65 : _GEN_364; // @[execute.scala 79:10:@1871.4]
  assign _GEN_366 = 6'h2e == _T_188 ? _T_66 : _GEN_365; // @[execute.scala 79:10:@1871.4]
  assign _GEN_367 = 6'h2f == _T_188 ? _T_67 : _GEN_366; // @[execute.scala 79:10:@1871.4]
  assign _GEN_368 = 6'h30 == _T_188 ? _T_68 : _GEN_367; // @[execute.scala 79:10:@1871.4]
  assign _GEN_369 = 6'h31 == _T_188 ? _T_69 : _GEN_368; // @[execute.scala 79:10:@1871.4]
  assign _GEN_370 = 6'h32 == _T_188 ? _T_70 : _GEN_369; // @[execute.scala 79:10:@1871.4]
  assign _GEN_371 = 6'h33 == _T_188 ? _T_71 : _GEN_370; // @[execute.scala 79:10:@1871.4]
  assign _GEN_372 = 6'h34 == _T_188 ? _T_72 : _GEN_371; // @[execute.scala 79:10:@1871.4]
  assign _GEN_373 = 6'h35 == _T_188 ? _T_73 : _GEN_372; // @[execute.scala 79:10:@1871.4]
  assign _GEN_374 = 6'h36 == _T_188 ? _T_74 : _GEN_373; // @[execute.scala 79:10:@1871.4]
  assign _GEN_375 = 6'h37 == _T_188 ? _T_75 : _GEN_374; // @[execute.scala 79:10:@1871.4]
  assign _GEN_376 = 6'h38 == _T_188 ? _T_76 : _GEN_375; // @[execute.scala 79:10:@1871.4]
  assign _GEN_377 = 6'h39 == _T_188 ? _T_77 : _GEN_376; // @[execute.scala 79:10:@1871.4]
  assign _GEN_378 = 6'h3a == _T_188 ? _T_78 : _GEN_377; // @[execute.scala 79:10:@1871.4]
  assign _GEN_379 = 6'h3b == _T_188 ? _T_79 : _GEN_378; // @[execute.scala 79:10:@1871.4]
  assign _GEN_380 = 6'h3c == _T_188 ? _T_80 : _GEN_379; // @[execute.scala 79:10:@1871.4]
  assign _GEN_381 = 6'h3d == _T_188 ? _T_81 : _GEN_380; // @[execute.scala 79:10:@1871.4]
  assign _GEN_382 = 6'h3e == _T_188 ? _T_82 : _GEN_381; // @[execute.scala 79:10:@1871.4]
  assign _GEN_383 = 6'h3f == _T_188 ? _T_83 : _GEN_382; // @[execute.scala 79:10:@1871.4]
  assign _T_190 = _T_180 ? _GEN_319 : _GEN_383; // @[execute.scala 79:10:@1871.4]
  assign _T_192 = io_amount < 6'h3d; // @[execute.scala 79:15:@1872.4]
  assign _T_194 = io_amount - 6'h3d; // @[execute.scala 79:37:@1873.4]
  assign _T_195 = $unsigned(_T_194); // @[execute.scala 79:37:@1874.4]
  assign _T_196 = _T_195[5:0]; // @[execute.scala 79:37:@1875.4]
  assign _T_199 = 6'h3 + io_amount; // @[execute.scala 79:60:@1876.4]
  assign _T_200 = 6'h3 + io_amount; // @[execute.scala 79:60:@1877.4]
  assign _GEN_385 = 6'h1 == _T_196 ? _T_21 : _T_20; // @[execute.scala 79:10:@1878.4]
  assign _GEN_386 = 6'h2 == _T_196 ? _T_22 : _GEN_385; // @[execute.scala 79:10:@1878.4]
  assign _GEN_387 = 6'h3 == _T_196 ? _T_23 : _GEN_386; // @[execute.scala 79:10:@1878.4]
  assign _GEN_388 = 6'h4 == _T_196 ? _T_24 : _GEN_387; // @[execute.scala 79:10:@1878.4]
  assign _GEN_389 = 6'h5 == _T_196 ? _T_25 : _GEN_388; // @[execute.scala 79:10:@1878.4]
  assign _GEN_390 = 6'h6 == _T_196 ? _T_26 : _GEN_389; // @[execute.scala 79:10:@1878.4]
  assign _GEN_391 = 6'h7 == _T_196 ? _T_27 : _GEN_390; // @[execute.scala 79:10:@1878.4]
  assign _GEN_392 = 6'h8 == _T_196 ? _T_28 : _GEN_391; // @[execute.scala 79:10:@1878.4]
  assign _GEN_393 = 6'h9 == _T_196 ? _T_29 : _GEN_392; // @[execute.scala 79:10:@1878.4]
  assign _GEN_394 = 6'ha == _T_196 ? _T_30 : _GEN_393; // @[execute.scala 79:10:@1878.4]
  assign _GEN_395 = 6'hb == _T_196 ? _T_31 : _GEN_394; // @[execute.scala 79:10:@1878.4]
  assign _GEN_396 = 6'hc == _T_196 ? _T_32 : _GEN_395; // @[execute.scala 79:10:@1878.4]
  assign _GEN_397 = 6'hd == _T_196 ? _T_33 : _GEN_396; // @[execute.scala 79:10:@1878.4]
  assign _GEN_398 = 6'he == _T_196 ? _T_34 : _GEN_397; // @[execute.scala 79:10:@1878.4]
  assign _GEN_399 = 6'hf == _T_196 ? _T_35 : _GEN_398; // @[execute.scala 79:10:@1878.4]
  assign _GEN_400 = 6'h10 == _T_196 ? _T_36 : _GEN_399; // @[execute.scala 79:10:@1878.4]
  assign _GEN_401 = 6'h11 == _T_196 ? _T_37 : _GEN_400; // @[execute.scala 79:10:@1878.4]
  assign _GEN_402 = 6'h12 == _T_196 ? _T_38 : _GEN_401; // @[execute.scala 79:10:@1878.4]
  assign _GEN_403 = 6'h13 == _T_196 ? _T_39 : _GEN_402; // @[execute.scala 79:10:@1878.4]
  assign _GEN_404 = 6'h14 == _T_196 ? _T_40 : _GEN_403; // @[execute.scala 79:10:@1878.4]
  assign _GEN_405 = 6'h15 == _T_196 ? _T_41 : _GEN_404; // @[execute.scala 79:10:@1878.4]
  assign _GEN_406 = 6'h16 == _T_196 ? _T_42 : _GEN_405; // @[execute.scala 79:10:@1878.4]
  assign _GEN_407 = 6'h17 == _T_196 ? _T_43 : _GEN_406; // @[execute.scala 79:10:@1878.4]
  assign _GEN_408 = 6'h18 == _T_196 ? _T_44 : _GEN_407; // @[execute.scala 79:10:@1878.4]
  assign _GEN_409 = 6'h19 == _T_196 ? _T_45 : _GEN_408; // @[execute.scala 79:10:@1878.4]
  assign _GEN_410 = 6'h1a == _T_196 ? _T_46 : _GEN_409; // @[execute.scala 79:10:@1878.4]
  assign _GEN_411 = 6'h1b == _T_196 ? _T_47 : _GEN_410; // @[execute.scala 79:10:@1878.4]
  assign _GEN_412 = 6'h1c == _T_196 ? _T_48 : _GEN_411; // @[execute.scala 79:10:@1878.4]
  assign _GEN_413 = 6'h1d == _T_196 ? _T_49 : _GEN_412; // @[execute.scala 79:10:@1878.4]
  assign _GEN_414 = 6'h1e == _T_196 ? _T_50 : _GEN_413; // @[execute.scala 79:10:@1878.4]
  assign _GEN_415 = 6'h1f == _T_196 ? _T_51 : _GEN_414; // @[execute.scala 79:10:@1878.4]
  assign _GEN_416 = 6'h20 == _T_196 ? _T_52 : _GEN_415; // @[execute.scala 79:10:@1878.4]
  assign _GEN_417 = 6'h21 == _T_196 ? _T_53 : _GEN_416; // @[execute.scala 79:10:@1878.4]
  assign _GEN_418 = 6'h22 == _T_196 ? _T_54 : _GEN_417; // @[execute.scala 79:10:@1878.4]
  assign _GEN_419 = 6'h23 == _T_196 ? _T_55 : _GEN_418; // @[execute.scala 79:10:@1878.4]
  assign _GEN_420 = 6'h24 == _T_196 ? _T_56 : _GEN_419; // @[execute.scala 79:10:@1878.4]
  assign _GEN_421 = 6'h25 == _T_196 ? _T_57 : _GEN_420; // @[execute.scala 79:10:@1878.4]
  assign _GEN_422 = 6'h26 == _T_196 ? _T_58 : _GEN_421; // @[execute.scala 79:10:@1878.4]
  assign _GEN_423 = 6'h27 == _T_196 ? _T_59 : _GEN_422; // @[execute.scala 79:10:@1878.4]
  assign _GEN_424 = 6'h28 == _T_196 ? _T_60 : _GEN_423; // @[execute.scala 79:10:@1878.4]
  assign _GEN_425 = 6'h29 == _T_196 ? _T_61 : _GEN_424; // @[execute.scala 79:10:@1878.4]
  assign _GEN_426 = 6'h2a == _T_196 ? _T_62 : _GEN_425; // @[execute.scala 79:10:@1878.4]
  assign _GEN_427 = 6'h2b == _T_196 ? _T_63 : _GEN_426; // @[execute.scala 79:10:@1878.4]
  assign _GEN_428 = 6'h2c == _T_196 ? _T_64 : _GEN_427; // @[execute.scala 79:10:@1878.4]
  assign _GEN_429 = 6'h2d == _T_196 ? _T_65 : _GEN_428; // @[execute.scala 79:10:@1878.4]
  assign _GEN_430 = 6'h2e == _T_196 ? _T_66 : _GEN_429; // @[execute.scala 79:10:@1878.4]
  assign _GEN_431 = 6'h2f == _T_196 ? _T_67 : _GEN_430; // @[execute.scala 79:10:@1878.4]
  assign _GEN_432 = 6'h30 == _T_196 ? _T_68 : _GEN_431; // @[execute.scala 79:10:@1878.4]
  assign _GEN_433 = 6'h31 == _T_196 ? _T_69 : _GEN_432; // @[execute.scala 79:10:@1878.4]
  assign _GEN_434 = 6'h32 == _T_196 ? _T_70 : _GEN_433; // @[execute.scala 79:10:@1878.4]
  assign _GEN_435 = 6'h33 == _T_196 ? _T_71 : _GEN_434; // @[execute.scala 79:10:@1878.4]
  assign _GEN_436 = 6'h34 == _T_196 ? _T_72 : _GEN_435; // @[execute.scala 79:10:@1878.4]
  assign _GEN_437 = 6'h35 == _T_196 ? _T_73 : _GEN_436; // @[execute.scala 79:10:@1878.4]
  assign _GEN_438 = 6'h36 == _T_196 ? _T_74 : _GEN_437; // @[execute.scala 79:10:@1878.4]
  assign _GEN_439 = 6'h37 == _T_196 ? _T_75 : _GEN_438; // @[execute.scala 79:10:@1878.4]
  assign _GEN_440 = 6'h38 == _T_196 ? _T_76 : _GEN_439; // @[execute.scala 79:10:@1878.4]
  assign _GEN_441 = 6'h39 == _T_196 ? _T_77 : _GEN_440; // @[execute.scala 79:10:@1878.4]
  assign _GEN_442 = 6'h3a == _T_196 ? _T_78 : _GEN_441; // @[execute.scala 79:10:@1878.4]
  assign _GEN_443 = 6'h3b == _T_196 ? _T_79 : _GEN_442; // @[execute.scala 79:10:@1878.4]
  assign _GEN_444 = 6'h3c == _T_196 ? _T_80 : _GEN_443; // @[execute.scala 79:10:@1878.4]
  assign _GEN_445 = 6'h3d == _T_196 ? _T_81 : _GEN_444; // @[execute.scala 79:10:@1878.4]
  assign _GEN_446 = 6'h3e == _T_196 ? _T_82 : _GEN_445; // @[execute.scala 79:10:@1878.4]
  assign _GEN_447 = 6'h3f == _T_196 ? _T_83 : _GEN_446; // @[execute.scala 79:10:@1878.4]
  assign _GEN_449 = 6'h1 == _T_200 ? _T_21 : _T_20; // @[execute.scala 79:10:@1878.4]
  assign _GEN_450 = 6'h2 == _T_200 ? _T_22 : _GEN_449; // @[execute.scala 79:10:@1878.4]
  assign _GEN_451 = 6'h3 == _T_200 ? _T_23 : _GEN_450; // @[execute.scala 79:10:@1878.4]
  assign _GEN_452 = 6'h4 == _T_200 ? _T_24 : _GEN_451; // @[execute.scala 79:10:@1878.4]
  assign _GEN_453 = 6'h5 == _T_200 ? _T_25 : _GEN_452; // @[execute.scala 79:10:@1878.4]
  assign _GEN_454 = 6'h6 == _T_200 ? _T_26 : _GEN_453; // @[execute.scala 79:10:@1878.4]
  assign _GEN_455 = 6'h7 == _T_200 ? _T_27 : _GEN_454; // @[execute.scala 79:10:@1878.4]
  assign _GEN_456 = 6'h8 == _T_200 ? _T_28 : _GEN_455; // @[execute.scala 79:10:@1878.4]
  assign _GEN_457 = 6'h9 == _T_200 ? _T_29 : _GEN_456; // @[execute.scala 79:10:@1878.4]
  assign _GEN_458 = 6'ha == _T_200 ? _T_30 : _GEN_457; // @[execute.scala 79:10:@1878.4]
  assign _GEN_459 = 6'hb == _T_200 ? _T_31 : _GEN_458; // @[execute.scala 79:10:@1878.4]
  assign _GEN_460 = 6'hc == _T_200 ? _T_32 : _GEN_459; // @[execute.scala 79:10:@1878.4]
  assign _GEN_461 = 6'hd == _T_200 ? _T_33 : _GEN_460; // @[execute.scala 79:10:@1878.4]
  assign _GEN_462 = 6'he == _T_200 ? _T_34 : _GEN_461; // @[execute.scala 79:10:@1878.4]
  assign _GEN_463 = 6'hf == _T_200 ? _T_35 : _GEN_462; // @[execute.scala 79:10:@1878.4]
  assign _GEN_464 = 6'h10 == _T_200 ? _T_36 : _GEN_463; // @[execute.scala 79:10:@1878.4]
  assign _GEN_465 = 6'h11 == _T_200 ? _T_37 : _GEN_464; // @[execute.scala 79:10:@1878.4]
  assign _GEN_466 = 6'h12 == _T_200 ? _T_38 : _GEN_465; // @[execute.scala 79:10:@1878.4]
  assign _GEN_467 = 6'h13 == _T_200 ? _T_39 : _GEN_466; // @[execute.scala 79:10:@1878.4]
  assign _GEN_468 = 6'h14 == _T_200 ? _T_40 : _GEN_467; // @[execute.scala 79:10:@1878.4]
  assign _GEN_469 = 6'h15 == _T_200 ? _T_41 : _GEN_468; // @[execute.scala 79:10:@1878.4]
  assign _GEN_470 = 6'h16 == _T_200 ? _T_42 : _GEN_469; // @[execute.scala 79:10:@1878.4]
  assign _GEN_471 = 6'h17 == _T_200 ? _T_43 : _GEN_470; // @[execute.scala 79:10:@1878.4]
  assign _GEN_472 = 6'h18 == _T_200 ? _T_44 : _GEN_471; // @[execute.scala 79:10:@1878.4]
  assign _GEN_473 = 6'h19 == _T_200 ? _T_45 : _GEN_472; // @[execute.scala 79:10:@1878.4]
  assign _GEN_474 = 6'h1a == _T_200 ? _T_46 : _GEN_473; // @[execute.scala 79:10:@1878.4]
  assign _GEN_475 = 6'h1b == _T_200 ? _T_47 : _GEN_474; // @[execute.scala 79:10:@1878.4]
  assign _GEN_476 = 6'h1c == _T_200 ? _T_48 : _GEN_475; // @[execute.scala 79:10:@1878.4]
  assign _GEN_477 = 6'h1d == _T_200 ? _T_49 : _GEN_476; // @[execute.scala 79:10:@1878.4]
  assign _GEN_478 = 6'h1e == _T_200 ? _T_50 : _GEN_477; // @[execute.scala 79:10:@1878.4]
  assign _GEN_479 = 6'h1f == _T_200 ? _T_51 : _GEN_478; // @[execute.scala 79:10:@1878.4]
  assign _GEN_480 = 6'h20 == _T_200 ? _T_52 : _GEN_479; // @[execute.scala 79:10:@1878.4]
  assign _GEN_481 = 6'h21 == _T_200 ? _T_53 : _GEN_480; // @[execute.scala 79:10:@1878.4]
  assign _GEN_482 = 6'h22 == _T_200 ? _T_54 : _GEN_481; // @[execute.scala 79:10:@1878.4]
  assign _GEN_483 = 6'h23 == _T_200 ? _T_55 : _GEN_482; // @[execute.scala 79:10:@1878.4]
  assign _GEN_484 = 6'h24 == _T_200 ? _T_56 : _GEN_483; // @[execute.scala 79:10:@1878.4]
  assign _GEN_485 = 6'h25 == _T_200 ? _T_57 : _GEN_484; // @[execute.scala 79:10:@1878.4]
  assign _GEN_486 = 6'h26 == _T_200 ? _T_58 : _GEN_485; // @[execute.scala 79:10:@1878.4]
  assign _GEN_487 = 6'h27 == _T_200 ? _T_59 : _GEN_486; // @[execute.scala 79:10:@1878.4]
  assign _GEN_488 = 6'h28 == _T_200 ? _T_60 : _GEN_487; // @[execute.scala 79:10:@1878.4]
  assign _GEN_489 = 6'h29 == _T_200 ? _T_61 : _GEN_488; // @[execute.scala 79:10:@1878.4]
  assign _GEN_490 = 6'h2a == _T_200 ? _T_62 : _GEN_489; // @[execute.scala 79:10:@1878.4]
  assign _GEN_491 = 6'h2b == _T_200 ? _T_63 : _GEN_490; // @[execute.scala 79:10:@1878.4]
  assign _GEN_492 = 6'h2c == _T_200 ? _T_64 : _GEN_491; // @[execute.scala 79:10:@1878.4]
  assign _GEN_493 = 6'h2d == _T_200 ? _T_65 : _GEN_492; // @[execute.scala 79:10:@1878.4]
  assign _GEN_494 = 6'h2e == _T_200 ? _T_66 : _GEN_493; // @[execute.scala 79:10:@1878.4]
  assign _GEN_495 = 6'h2f == _T_200 ? _T_67 : _GEN_494; // @[execute.scala 79:10:@1878.4]
  assign _GEN_496 = 6'h30 == _T_200 ? _T_68 : _GEN_495; // @[execute.scala 79:10:@1878.4]
  assign _GEN_497 = 6'h31 == _T_200 ? _T_69 : _GEN_496; // @[execute.scala 79:10:@1878.4]
  assign _GEN_498 = 6'h32 == _T_200 ? _T_70 : _GEN_497; // @[execute.scala 79:10:@1878.4]
  assign _GEN_499 = 6'h33 == _T_200 ? _T_71 : _GEN_498; // @[execute.scala 79:10:@1878.4]
  assign _GEN_500 = 6'h34 == _T_200 ? _T_72 : _GEN_499; // @[execute.scala 79:10:@1878.4]
  assign _GEN_501 = 6'h35 == _T_200 ? _T_73 : _GEN_500; // @[execute.scala 79:10:@1878.4]
  assign _GEN_502 = 6'h36 == _T_200 ? _T_74 : _GEN_501; // @[execute.scala 79:10:@1878.4]
  assign _GEN_503 = 6'h37 == _T_200 ? _T_75 : _GEN_502; // @[execute.scala 79:10:@1878.4]
  assign _GEN_504 = 6'h38 == _T_200 ? _T_76 : _GEN_503; // @[execute.scala 79:10:@1878.4]
  assign _GEN_505 = 6'h39 == _T_200 ? _T_77 : _GEN_504; // @[execute.scala 79:10:@1878.4]
  assign _GEN_506 = 6'h3a == _T_200 ? _T_78 : _GEN_505; // @[execute.scala 79:10:@1878.4]
  assign _GEN_507 = 6'h3b == _T_200 ? _T_79 : _GEN_506; // @[execute.scala 79:10:@1878.4]
  assign _GEN_508 = 6'h3c == _T_200 ? _T_80 : _GEN_507; // @[execute.scala 79:10:@1878.4]
  assign _GEN_509 = 6'h3d == _T_200 ? _T_81 : _GEN_508; // @[execute.scala 79:10:@1878.4]
  assign _GEN_510 = 6'h3e == _T_200 ? _T_82 : _GEN_509; // @[execute.scala 79:10:@1878.4]
  assign _GEN_511 = 6'h3f == _T_200 ? _T_83 : _GEN_510; // @[execute.scala 79:10:@1878.4]
  assign _T_202 = _T_192 ? _GEN_447 : _GEN_511; // @[execute.scala 79:10:@1878.4]
  assign _T_204 = io_amount < 6'h3c; // @[execute.scala 79:15:@1879.4]
  assign _T_206 = io_amount - 6'h3c; // @[execute.scala 79:37:@1880.4]
  assign _T_207 = $unsigned(_T_206); // @[execute.scala 79:37:@1881.4]
  assign _T_208 = _T_207[5:0]; // @[execute.scala 79:37:@1882.4]
  assign _T_211 = 6'h4 + io_amount; // @[execute.scala 79:60:@1883.4]
  assign _T_212 = 6'h4 + io_amount; // @[execute.scala 79:60:@1884.4]
  assign _GEN_513 = 6'h1 == _T_208 ? _T_21 : _T_20; // @[execute.scala 79:10:@1885.4]
  assign _GEN_514 = 6'h2 == _T_208 ? _T_22 : _GEN_513; // @[execute.scala 79:10:@1885.4]
  assign _GEN_515 = 6'h3 == _T_208 ? _T_23 : _GEN_514; // @[execute.scala 79:10:@1885.4]
  assign _GEN_516 = 6'h4 == _T_208 ? _T_24 : _GEN_515; // @[execute.scala 79:10:@1885.4]
  assign _GEN_517 = 6'h5 == _T_208 ? _T_25 : _GEN_516; // @[execute.scala 79:10:@1885.4]
  assign _GEN_518 = 6'h6 == _T_208 ? _T_26 : _GEN_517; // @[execute.scala 79:10:@1885.4]
  assign _GEN_519 = 6'h7 == _T_208 ? _T_27 : _GEN_518; // @[execute.scala 79:10:@1885.4]
  assign _GEN_520 = 6'h8 == _T_208 ? _T_28 : _GEN_519; // @[execute.scala 79:10:@1885.4]
  assign _GEN_521 = 6'h9 == _T_208 ? _T_29 : _GEN_520; // @[execute.scala 79:10:@1885.4]
  assign _GEN_522 = 6'ha == _T_208 ? _T_30 : _GEN_521; // @[execute.scala 79:10:@1885.4]
  assign _GEN_523 = 6'hb == _T_208 ? _T_31 : _GEN_522; // @[execute.scala 79:10:@1885.4]
  assign _GEN_524 = 6'hc == _T_208 ? _T_32 : _GEN_523; // @[execute.scala 79:10:@1885.4]
  assign _GEN_525 = 6'hd == _T_208 ? _T_33 : _GEN_524; // @[execute.scala 79:10:@1885.4]
  assign _GEN_526 = 6'he == _T_208 ? _T_34 : _GEN_525; // @[execute.scala 79:10:@1885.4]
  assign _GEN_527 = 6'hf == _T_208 ? _T_35 : _GEN_526; // @[execute.scala 79:10:@1885.4]
  assign _GEN_528 = 6'h10 == _T_208 ? _T_36 : _GEN_527; // @[execute.scala 79:10:@1885.4]
  assign _GEN_529 = 6'h11 == _T_208 ? _T_37 : _GEN_528; // @[execute.scala 79:10:@1885.4]
  assign _GEN_530 = 6'h12 == _T_208 ? _T_38 : _GEN_529; // @[execute.scala 79:10:@1885.4]
  assign _GEN_531 = 6'h13 == _T_208 ? _T_39 : _GEN_530; // @[execute.scala 79:10:@1885.4]
  assign _GEN_532 = 6'h14 == _T_208 ? _T_40 : _GEN_531; // @[execute.scala 79:10:@1885.4]
  assign _GEN_533 = 6'h15 == _T_208 ? _T_41 : _GEN_532; // @[execute.scala 79:10:@1885.4]
  assign _GEN_534 = 6'h16 == _T_208 ? _T_42 : _GEN_533; // @[execute.scala 79:10:@1885.4]
  assign _GEN_535 = 6'h17 == _T_208 ? _T_43 : _GEN_534; // @[execute.scala 79:10:@1885.4]
  assign _GEN_536 = 6'h18 == _T_208 ? _T_44 : _GEN_535; // @[execute.scala 79:10:@1885.4]
  assign _GEN_537 = 6'h19 == _T_208 ? _T_45 : _GEN_536; // @[execute.scala 79:10:@1885.4]
  assign _GEN_538 = 6'h1a == _T_208 ? _T_46 : _GEN_537; // @[execute.scala 79:10:@1885.4]
  assign _GEN_539 = 6'h1b == _T_208 ? _T_47 : _GEN_538; // @[execute.scala 79:10:@1885.4]
  assign _GEN_540 = 6'h1c == _T_208 ? _T_48 : _GEN_539; // @[execute.scala 79:10:@1885.4]
  assign _GEN_541 = 6'h1d == _T_208 ? _T_49 : _GEN_540; // @[execute.scala 79:10:@1885.4]
  assign _GEN_542 = 6'h1e == _T_208 ? _T_50 : _GEN_541; // @[execute.scala 79:10:@1885.4]
  assign _GEN_543 = 6'h1f == _T_208 ? _T_51 : _GEN_542; // @[execute.scala 79:10:@1885.4]
  assign _GEN_544 = 6'h20 == _T_208 ? _T_52 : _GEN_543; // @[execute.scala 79:10:@1885.4]
  assign _GEN_545 = 6'h21 == _T_208 ? _T_53 : _GEN_544; // @[execute.scala 79:10:@1885.4]
  assign _GEN_546 = 6'h22 == _T_208 ? _T_54 : _GEN_545; // @[execute.scala 79:10:@1885.4]
  assign _GEN_547 = 6'h23 == _T_208 ? _T_55 : _GEN_546; // @[execute.scala 79:10:@1885.4]
  assign _GEN_548 = 6'h24 == _T_208 ? _T_56 : _GEN_547; // @[execute.scala 79:10:@1885.4]
  assign _GEN_549 = 6'h25 == _T_208 ? _T_57 : _GEN_548; // @[execute.scala 79:10:@1885.4]
  assign _GEN_550 = 6'h26 == _T_208 ? _T_58 : _GEN_549; // @[execute.scala 79:10:@1885.4]
  assign _GEN_551 = 6'h27 == _T_208 ? _T_59 : _GEN_550; // @[execute.scala 79:10:@1885.4]
  assign _GEN_552 = 6'h28 == _T_208 ? _T_60 : _GEN_551; // @[execute.scala 79:10:@1885.4]
  assign _GEN_553 = 6'h29 == _T_208 ? _T_61 : _GEN_552; // @[execute.scala 79:10:@1885.4]
  assign _GEN_554 = 6'h2a == _T_208 ? _T_62 : _GEN_553; // @[execute.scala 79:10:@1885.4]
  assign _GEN_555 = 6'h2b == _T_208 ? _T_63 : _GEN_554; // @[execute.scala 79:10:@1885.4]
  assign _GEN_556 = 6'h2c == _T_208 ? _T_64 : _GEN_555; // @[execute.scala 79:10:@1885.4]
  assign _GEN_557 = 6'h2d == _T_208 ? _T_65 : _GEN_556; // @[execute.scala 79:10:@1885.4]
  assign _GEN_558 = 6'h2e == _T_208 ? _T_66 : _GEN_557; // @[execute.scala 79:10:@1885.4]
  assign _GEN_559 = 6'h2f == _T_208 ? _T_67 : _GEN_558; // @[execute.scala 79:10:@1885.4]
  assign _GEN_560 = 6'h30 == _T_208 ? _T_68 : _GEN_559; // @[execute.scala 79:10:@1885.4]
  assign _GEN_561 = 6'h31 == _T_208 ? _T_69 : _GEN_560; // @[execute.scala 79:10:@1885.4]
  assign _GEN_562 = 6'h32 == _T_208 ? _T_70 : _GEN_561; // @[execute.scala 79:10:@1885.4]
  assign _GEN_563 = 6'h33 == _T_208 ? _T_71 : _GEN_562; // @[execute.scala 79:10:@1885.4]
  assign _GEN_564 = 6'h34 == _T_208 ? _T_72 : _GEN_563; // @[execute.scala 79:10:@1885.4]
  assign _GEN_565 = 6'h35 == _T_208 ? _T_73 : _GEN_564; // @[execute.scala 79:10:@1885.4]
  assign _GEN_566 = 6'h36 == _T_208 ? _T_74 : _GEN_565; // @[execute.scala 79:10:@1885.4]
  assign _GEN_567 = 6'h37 == _T_208 ? _T_75 : _GEN_566; // @[execute.scala 79:10:@1885.4]
  assign _GEN_568 = 6'h38 == _T_208 ? _T_76 : _GEN_567; // @[execute.scala 79:10:@1885.4]
  assign _GEN_569 = 6'h39 == _T_208 ? _T_77 : _GEN_568; // @[execute.scala 79:10:@1885.4]
  assign _GEN_570 = 6'h3a == _T_208 ? _T_78 : _GEN_569; // @[execute.scala 79:10:@1885.4]
  assign _GEN_571 = 6'h3b == _T_208 ? _T_79 : _GEN_570; // @[execute.scala 79:10:@1885.4]
  assign _GEN_572 = 6'h3c == _T_208 ? _T_80 : _GEN_571; // @[execute.scala 79:10:@1885.4]
  assign _GEN_573 = 6'h3d == _T_208 ? _T_81 : _GEN_572; // @[execute.scala 79:10:@1885.4]
  assign _GEN_574 = 6'h3e == _T_208 ? _T_82 : _GEN_573; // @[execute.scala 79:10:@1885.4]
  assign _GEN_575 = 6'h3f == _T_208 ? _T_83 : _GEN_574; // @[execute.scala 79:10:@1885.4]
  assign _GEN_577 = 6'h1 == _T_212 ? _T_21 : _T_20; // @[execute.scala 79:10:@1885.4]
  assign _GEN_578 = 6'h2 == _T_212 ? _T_22 : _GEN_577; // @[execute.scala 79:10:@1885.4]
  assign _GEN_579 = 6'h3 == _T_212 ? _T_23 : _GEN_578; // @[execute.scala 79:10:@1885.4]
  assign _GEN_580 = 6'h4 == _T_212 ? _T_24 : _GEN_579; // @[execute.scala 79:10:@1885.4]
  assign _GEN_581 = 6'h5 == _T_212 ? _T_25 : _GEN_580; // @[execute.scala 79:10:@1885.4]
  assign _GEN_582 = 6'h6 == _T_212 ? _T_26 : _GEN_581; // @[execute.scala 79:10:@1885.4]
  assign _GEN_583 = 6'h7 == _T_212 ? _T_27 : _GEN_582; // @[execute.scala 79:10:@1885.4]
  assign _GEN_584 = 6'h8 == _T_212 ? _T_28 : _GEN_583; // @[execute.scala 79:10:@1885.4]
  assign _GEN_585 = 6'h9 == _T_212 ? _T_29 : _GEN_584; // @[execute.scala 79:10:@1885.4]
  assign _GEN_586 = 6'ha == _T_212 ? _T_30 : _GEN_585; // @[execute.scala 79:10:@1885.4]
  assign _GEN_587 = 6'hb == _T_212 ? _T_31 : _GEN_586; // @[execute.scala 79:10:@1885.4]
  assign _GEN_588 = 6'hc == _T_212 ? _T_32 : _GEN_587; // @[execute.scala 79:10:@1885.4]
  assign _GEN_589 = 6'hd == _T_212 ? _T_33 : _GEN_588; // @[execute.scala 79:10:@1885.4]
  assign _GEN_590 = 6'he == _T_212 ? _T_34 : _GEN_589; // @[execute.scala 79:10:@1885.4]
  assign _GEN_591 = 6'hf == _T_212 ? _T_35 : _GEN_590; // @[execute.scala 79:10:@1885.4]
  assign _GEN_592 = 6'h10 == _T_212 ? _T_36 : _GEN_591; // @[execute.scala 79:10:@1885.4]
  assign _GEN_593 = 6'h11 == _T_212 ? _T_37 : _GEN_592; // @[execute.scala 79:10:@1885.4]
  assign _GEN_594 = 6'h12 == _T_212 ? _T_38 : _GEN_593; // @[execute.scala 79:10:@1885.4]
  assign _GEN_595 = 6'h13 == _T_212 ? _T_39 : _GEN_594; // @[execute.scala 79:10:@1885.4]
  assign _GEN_596 = 6'h14 == _T_212 ? _T_40 : _GEN_595; // @[execute.scala 79:10:@1885.4]
  assign _GEN_597 = 6'h15 == _T_212 ? _T_41 : _GEN_596; // @[execute.scala 79:10:@1885.4]
  assign _GEN_598 = 6'h16 == _T_212 ? _T_42 : _GEN_597; // @[execute.scala 79:10:@1885.4]
  assign _GEN_599 = 6'h17 == _T_212 ? _T_43 : _GEN_598; // @[execute.scala 79:10:@1885.4]
  assign _GEN_600 = 6'h18 == _T_212 ? _T_44 : _GEN_599; // @[execute.scala 79:10:@1885.4]
  assign _GEN_601 = 6'h19 == _T_212 ? _T_45 : _GEN_600; // @[execute.scala 79:10:@1885.4]
  assign _GEN_602 = 6'h1a == _T_212 ? _T_46 : _GEN_601; // @[execute.scala 79:10:@1885.4]
  assign _GEN_603 = 6'h1b == _T_212 ? _T_47 : _GEN_602; // @[execute.scala 79:10:@1885.4]
  assign _GEN_604 = 6'h1c == _T_212 ? _T_48 : _GEN_603; // @[execute.scala 79:10:@1885.4]
  assign _GEN_605 = 6'h1d == _T_212 ? _T_49 : _GEN_604; // @[execute.scala 79:10:@1885.4]
  assign _GEN_606 = 6'h1e == _T_212 ? _T_50 : _GEN_605; // @[execute.scala 79:10:@1885.4]
  assign _GEN_607 = 6'h1f == _T_212 ? _T_51 : _GEN_606; // @[execute.scala 79:10:@1885.4]
  assign _GEN_608 = 6'h20 == _T_212 ? _T_52 : _GEN_607; // @[execute.scala 79:10:@1885.4]
  assign _GEN_609 = 6'h21 == _T_212 ? _T_53 : _GEN_608; // @[execute.scala 79:10:@1885.4]
  assign _GEN_610 = 6'h22 == _T_212 ? _T_54 : _GEN_609; // @[execute.scala 79:10:@1885.4]
  assign _GEN_611 = 6'h23 == _T_212 ? _T_55 : _GEN_610; // @[execute.scala 79:10:@1885.4]
  assign _GEN_612 = 6'h24 == _T_212 ? _T_56 : _GEN_611; // @[execute.scala 79:10:@1885.4]
  assign _GEN_613 = 6'h25 == _T_212 ? _T_57 : _GEN_612; // @[execute.scala 79:10:@1885.4]
  assign _GEN_614 = 6'h26 == _T_212 ? _T_58 : _GEN_613; // @[execute.scala 79:10:@1885.4]
  assign _GEN_615 = 6'h27 == _T_212 ? _T_59 : _GEN_614; // @[execute.scala 79:10:@1885.4]
  assign _GEN_616 = 6'h28 == _T_212 ? _T_60 : _GEN_615; // @[execute.scala 79:10:@1885.4]
  assign _GEN_617 = 6'h29 == _T_212 ? _T_61 : _GEN_616; // @[execute.scala 79:10:@1885.4]
  assign _GEN_618 = 6'h2a == _T_212 ? _T_62 : _GEN_617; // @[execute.scala 79:10:@1885.4]
  assign _GEN_619 = 6'h2b == _T_212 ? _T_63 : _GEN_618; // @[execute.scala 79:10:@1885.4]
  assign _GEN_620 = 6'h2c == _T_212 ? _T_64 : _GEN_619; // @[execute.scala 79:10:@1885.4]
  assign _GEN_621 = 6'h2d == _T_212 ? _T_65 : _GEN_620; // @[execute.scala 79:10:@1885.4]
  assign _GEN_622 = 6'h2e == _T_212 ? _T_66 : _GEN_621; // @[execute.scala 79:10:@1885.4]
  assign _GEN_623 = 6'h2f == _T_212 ? _T_67 : _GEN_622; // @[execute.scala 79:10:@1885.4]
  assign _GEN_624 = 6'h30 == _T_212 ? _T_68 : _GEN_623; // @[execute.scala 79:10:@1885.4]
  assign _GEN_625 = 6'h31 == _T_212 ? _T_69 : _GEN_624; // @[execute.scala 79:10:@1885.4]
  assign _GEN_626 = 6'h32 == _T_212 ? _T_70 : _GEN_625; // @[execute.scala 79:10:@1885.4]
  assign _GEN_627 = 6'h33 == _T_212 ? _T_71 : _GEN_626; // @[execute.scala 79:10:@1885.4]
  assign _GEN_628 = 6'h34 == _T_212 ? _T_72 : _GEN_627; // @[execute.scala 79:10:@1885.4]
  assign _GEN_629 = 6'h35 == _T_212 ? _T_73 : _GEN_628; // @[execute.scala 79:10:@1885.4]
  assign _GEN_630 = 6'h36 == _T_212 ? _T_74 : _GEN_629; // @[execute.scala 79:10:@1885.4]
  assign _GEN_631 = 6'h37 == _T_212 ? _T_75 : _GEN_630; // @[execute.scala 79:10:@1885.4]
  assign _GEN_632 = 6'h38 == _T_212 ? _T_76 : _GEN_631; // @[execute.scala 79:10:@1885.4]
  assign _GEN_633 = 6'h39 == _T_212 ? _T_77 : _GEN_632; // @[execute.scala 79:10:@1885.4]
  assign _GEN_634 = 6'h3a == _T_212 ? _T_78 : _GEN_633; // @[execute.scala 79:10:@1885.4]
  assign _GEN_635 = 6'h3b == _T_212 ? _T_79 : _GEN_634; // @[execute.scala 79:10:@1885.4]
  assign _GEN_636 = 6'h3c == _T_212 ? _T_80 : _GEN_635; // @[execute.scala 79:10:@1885.4]
  assign _GEN_637 = 6'h3d == _T_212 ? _T_81 : _GEN_636; // @[execute.scala 79:10:@1885.4]
  assign _GEN_638 = 6'h3e == _T_212 ? _T_82 : _GEN_637; // @[execute.scala 79:10:@1885.4]
  assign _GEN_639 = 6'h3f == _T_212 ? _T_83 : _GEN_638; // @[execute.scala 79:10:@1885.4]
  assign _T_214 = _T_204 ? _GEN_575 : _GEN_639; // @[execute.scala 79:10:@1885.4]
  assign _T_216 = io_amount < 6'h3b; // @[execute.scala 79:15:@1886.4]
  assign _T_218 = io_amount - 6'h3b; // @[execute.scala 79:37:@1887.4]
  assign _T_219 = $unsigned(_T_218); // @[execute.scala 79:37:@1888.4]
  assign _T_220 = _T_219[5:0]; // @[execute.scala 79:37:@1889.4]
  assign _T_223 = 6'h5 + io_amount; // @[execute.scala 79:60:@1890.4]
  assign _T_224 = 6'h5 + io_amount; // @[execute.scala 79:60:@1891.4]
  assign _GEN_641 = 6'h1 == _T_220 ? _T_21 : _T_20; // @[execute.scala 79:10:@1892.4]
  assign _GEN_642 = 6'h2 == _T_220 ? _T_22 : _GEN_641; // @[execute.scala 79:10:@1892.4]
  assign _GEN_643 = 6'h3 == _T_220 ? _T_23 : _GEN_642; // @[execute.scala 79:10:@1892.4]
  assign _GEN_644 = 6'h4 == _T_220 ? _T_24 : _GEN_643; // @[execute.scala 79:10:@1892.4]
  assign _GEN_645 = 6'h5 == _T_220 ? _T_25 : _GEN_644; // @[execute.scala 79:10:@1892.4]
  assign _GEN_646 = 6'h6 == _T_220 ? _T_26 : _GEN_645; // @[execute.scala 79:10:@1892.4]
  assign _GEN_647 = 6'h7 == _T_220 ? _T_27 : _GEN_646; // @[execute.scala 79:10:@1892.4]
  assign _GEN_648 = 6'h8 == _T_220 ? _T_28 : _GEN_647; // @[execute.scala 79:10:@1892.4]
  assign _GEN_649 = 6'h9 == _T_220 ? _T_29 : _GEN_648; // @[execute.scala 79:10:@1892.4]
  assign _GEN_650 = 6'ha == _T_220 ? _T_30 : _GEN_649; // @[execute.scala 79:10:@1892.4]
  assign _GEN_651 = 6'hb == _T_220 ? _T_31 : _GEN_650; // @[execute.scala 79:10:@1892.4]
  assign _GEN_652 = 6'hc == _T_220 ? _T_32 : _GEN_651; // @[execute.scala 79:10:@1892.4]
  assign _GEN_653 = 6'hd == _T_220 ? _T_33 : _GEN_652; // @[execute.scala 79:10:@1892.4]
  assign _GEN_654 = 6'he == _T_220 ? _T_34 : _GEN_653; // @[execute.scala 79:10:@1892.4]
  assign _GEN_655 = 6'hf == _T_220 ? _T_35 : _GEN_654; // @[execute.scala 79:10:@1892.4]
  assign _GEN_656 = 6'h10 == _T_220 ? _T_36 : _GEN_655; // @[execute.scala 79:10:@1892.4]
  assign _GEN_657 = 6'h11 == _T_220 ? _T_37 : _GEN_656; // @[execute.scala 79:10:@1892.4]
  assign _GEN_658 = 6'h12 == _T_220 ? _T_38 : _GEN_657; // @[execute.scala 79:10:@1892.4]
  assign _GEN_659 = 6'h13 == _T_220 ? _T_39 : _GEN_658; // @[execute.scala 79:10:@1892.4]
  assign _GEN_660 = 6'h14 == _T_220 ? _T_40 : _GEN_659; // @[execute.scala 79:10:@1892.4]
  assign _GEN_661 = 6'h15 == _T_220 ? _T_41 : _GEN_660; // @[execute.scala 79:10:@1892.4]
  assign _GEN_662 = 6'h16 == _T_220 ? _T_42 : _GEN_661; // @[execute.scala 79:10:@1892.4]
  assign _GEN_663 = 6'h17 == _T_220 ? _T_43 : _GEN_662; // @[execute.scala 79:10:@1892.4]
  assign _GEN_664 = 6'h18 == _T_220 ? _T_44 : _GEN_663; // @[execute.scala 79:10:@1892.4]
  assign _GEN_665 = 6'h19 == _T_220 ? _T_45 : _GEN_664; // @[execute.scala 79:10:@1892.4]
  assign _GEN_666 = 6'h1a == _T_220 ? _T_46 : _GEN_665; // @[execute.scala 79:10:@1892.4]
  assign _GEN_667 = 6'h1b == _T_220 ? _T_47 : _GEN_666; // @[execute.scala 79:10:@1892.4]
  assign _GEN_668 = 6'h1c == _T_220 ? _T_48 : _GEN_667; // @[execute.scala 79:10:@1892.4]
  assign _GEN_669 = 6'h1d == _T_220 ? _T_49 : _GEN_668; // @[execute.scala 79:10:@1892.4]
  assign _GEN_670 = 6'h1e == _T_220 ? _T_50 : _GEN_669; // @[execute.scala 79:10:@1892.4]
  assign _GEN_671 = 6'h1f == _T_220 ? _T_51 : _GEN_670; // @[execute.scala 79:10:@1892.4]
  assign _GEN_672 = 6'h20 == _T_220 ? _T_52 : _GEN_671; // @[execute.scala 79:10:@1892.4]
  assign _GEN_673 = 6'h21 == _T_220 ? _T_53 : _GEN_672; // @[execute.scala 79:10:@1892.4]
  assign _GEN_674 = 6'h22 == _T_220 ? _T_54 : _GEN_673; // @[execute.scala 79:10:@1892.4]
  assign _GEN_675 = 6'h23 == _T_220 ? _T_55 : _GEN_674; // @[execute.scala 79:10:@1892.4]
  assign _GEN_676 = 6'h24 == _T_220 ? _T_56 : _GEN_675; // @[execute.scala 79:10:@1892.4]
  assign _GEN_677 = 6'h25 == _T_220 ? _T_57 : _GEN_676; // @[execute.scala 79:10:@1892.4]
  assign _GEN_678 = 6'h26 == _T_220 ? _T_58 : _GEN_677; // @[execute.scala 79:10:@1892.4]
  assign _GEN_679 = 6'h27 == _T_220 ? _T_59 : _GEN_678; // @[execute.scala 79:10:@1892.4]
  assign _GEN_680 = 6'h28 == _T_220 ? _T_60 : _GEN_679; // @[execute.scala 79:10:@1892.4]
  assign _GEN_681 = 6'h29 == _T_220 ? _T_61 : _GEN_680; // @[execute.scala 79:10:@1892.4]
  assign _GEN_682 = 6'h2a == _T_220 ? _T_62 : _GEN_681; // @[execute.scala 79:10:@1892.4]
  assign _GEN_683 = 6'h2b == _T_220 ? _T_63 : _GEN_682; // @[execute.scala 79:10:@1892.4]
  assign _GEN_684 = 6'h2c == _T_220 ? _T_64 : _GEN_683; // @[execute.scala 79:10:@1892.4]
  assign _GEN_685 = 6'h2d == _T_220 ? _T_65 : _GEN_684; // @[execute.scala 79:10:@1892.4]
  assign _GEN_686 = 6'h2e == _T_220 ? _T_66 : _GEN_685; // @[execute.scala 79:10:@1892.4]
  assign _GEN_687 = 6'h2f == _T_220 ? _T_67 : _GEN_686; // @[execute.scala 79:10:@1892.4]
  assign _GEN_688 = 6'h30 == _T_220 ? _T_68 : _GEN_687; // @[execute.scala 79:10:@1892.4]
  assign _GEN_689 = 6'h31 == _T_220 ? _T_69 : _GEN_688; // @[execute.scala 79:10:@1892.4]
  assign _GEN_690 = 6'h32 == _T_220 ? _T_70 : _GEN_689; // @[execute.scala 79:10:@1892.4]
  assign _GEN_691 = 6'h33 == _T_220 ? _T_71 : _GEN_690; // @[execute.scala 79:10:@1892.4]
  assign _GEN_692 = 6'h34 == _T_220 ? _T_72 : _GEN_691; // @[execute.scala 79:10:@1892.4]
  assign _GEN_693 = 6'h35 == _T_220 ? _T_73 : _GEN_692; // @[execute.scala 79:10:@1892.4]
  assign _GEN_694 = 6'h36 == _T_220 ? _T_74 : _GEN_693; // @[execute.scala 79:10:@1892.4]
  assign _GEN_695 = 6'h37 == _T_220 ? _T_75 : _GEN_694; // @[execute.scala 79:10:@1892.4]
  assign _GEN_696 = 6'h38 == _T_220 ? _T_76 : _GEN_695; // @[execute.scala 79:10:@1892.4]
  assign _GEN_697 = 6'h39 == _T_220 ? _T_77 : _GEN_696; // @[execute.scala 79:10:@1892.4]
  assign _GEN_698 = 6'h3a == _T_220 ? _T_78 : _GEN_697; // @[execute.scala 79:10:@1892.4]
  assign _GEN_699 = 6'h3b == _T_220 ? _T_79 : _GEN_698; // @[execute.scala 79:10:@1892.4]
  assign _GEN_700 = 6'h3c == _T_220 ? _T_80 : _GEN_699; // @[execute.scala 79:10:@1892.4]
  assign _GEN_701 = 6'h3d == _T_220 ? _T_81 : _GEN_700; // @[execute.scala 79:10:@1892.4]
  assign _GEN_702 = 6'h3e == _T_220 ? _T_82 : _GEN_701; // @[execute.scala 79:10:@1892.4]
  assign _GEN_703 = 6'h3f == _T_220 ? _T_83 : _GEN_702; // @[execute.scala 79:10:@1892.4]
  assign _GEN_705 = 6'h1 == _T_224 ? _T_21 : _T_20; // @[execute.scala 79:10:@1892.4]
  assign _GEN_706 = 6'h2 == _T_224 ? _T_22 : _GEN_705; // @[execute.scala 79:10:@1892.4]
  assign _GEN_707 = 6'h3 == _T_224 ? _T_23 : _GEN_706; // @[execute.scala 79:10:@1892.4]
  assign _GEN_708 = 6'h4 == _T_224 ? _T_24 : _GEN_707; // @[execute.scala 79:10:@1892.4]
  assign _GEN_709 = 6'h5 == _T_224 ? _T_25 : _GEN_708; // @[execute.scala 79:10:@1892.4]
  assign _GEN_710 = 6'h6 == _T_224 ? _T_26 : _GEN_709; // @[execute.scala 79:10:@1892.4]
  assign _GEN_711 = 6'h7 == _T_224 ? _T_27 : _GEN_710; // @[execute.scala 79:10:@1892.4]
  assign _GEN_712 = 6'h8 == _T_224 ? _T_28 : _GEN_711; // @[execute.scala 79:10:@1892.4]
  assign _GEN_713 = 6'h9 == _T_224 ? _T_29 : _GEN_712; // @[execute.scala 79:10:@1892.4]
  assign _GEN_714 = 6'ha == _T_224 ? _T_30 : _GEN_713; // @[execute.scala 79:10:@1892.4]
  assign _GEN_715 = 6'hb == _T_224 ? _T_31 : _GEN_714; // @[execute.scala 79:10:@1892.4]
  assign _GEN_716 = 6'hc == _T_224 ? _T_32 : _GEN_715; // @[execute.scala 79:10:@1892.4]
  assign _GEN_717 = 6'hd == _T_224 ? _T_33 : _GEN_716; // @[execute.scala 79:10:@1892.4]
  assign _GEN_718 = 6'he == _T_224 ? _T_34 : _GEN_717; // @[execute.scala 79:10:@1892.4]
  assign _GEN_719 = 6'hf == _T_224 ? _T_35 : _GEN_718; // @[execute.scala 79:10:@1892.4]
  assign _GEN_720 = 6'h10 == _T_224 ? _T_36 : _GEN_719; // @[execute.scala 79:10:@1892.4]
  assign _GEN_721 = 6'h11 == _T_224 ? _T_37 : _GEN_720; // @[execute.scala 79:10:@1892.4]
  assign _GEN_722 = 6'h12 == _T_224 ? _T_38 : _GEN_721; // @[execute.scala 79:10:@1892.4]
  assign _GEN_723 = 6'h13 == _T_224 ? _T_39 : _GEN_722; // @[execute.scala 79:10:@1892.4]
  assign _GEN_724 = 6'h14 == _T_224 ? _T_40 : _GEN_723; // @[execute.scala 79:10:@1892.4]
  assign _GEN_725 = 6'h15 == _T_224 ? _T_41 : _GEN_724; // @[execute.scala 79:10:@1892.4]
  assign _GEN_726 = 6'h16 == _T_224 ? _T_42 : _GEN_725; // @[execute.scala 79:10:@1892.4]
  assign _GEN_727 = 6'h17 == _T_224 ? _T_43 : _GEN_726; // @[execute.scala 79:10:@1892.4]
  assign _GEN_728 = 6'h18 == _T_224 ? _T_44 : _GEN_727; // @[execute.scala 79:10:@1892.4]
  assign _GEN_729 = 6'h19 == _T_224 ? _T_45 : _GEN_728; // @[execute.scala 79:10:@1892.4]
  assign _GEN_730 = 6'h1a == _T_224 ? _T_46 : _GEN_729; // @[execute.scala 79:10:@1892.4]
  assign _GEN_731 = 6'h1b == _T_224 ? _T_47 : _GEN_730; // @[execute.scala 79:10:@1892.4]
  assign _GEN_732 = 6'h1c == _T_224 ? _T_48 : _GEN_731; // @[execute.scala 79:10:@1892.4]
  assign _GEN_733 = 6'h1d == _T_224 ? _T_49 : _GEN_732; // @[execute.scala 79:10:@1892.4]
  assign _GEN_734 = 6'h1e == _T_224 ? _T_50 : _GEN_733; // @[execute.scala 79:10:@1892.4]
  assign _GEN_735 = 6'h1f == _T_224 ? _T_51 : _GEN_734; // @[execute.scala 79:10:@1892.4]
  assign _GEN_736 = 6'h20 == _T_224 ? _T_52 : _GEN_735; // @[execute.scala 79:10:@1892.4]
  assign _GEN_737 = 6'h21 == _T_224 ? _T_53 : _GEN_736; // @[execute.scala 79:10:@1892.4]
  assign _GEN_738 = 6'h22 == _T_224 ? _T_54 : _GEN_737; // @[execute.scala 79:10:@1892.4]
  assign _GEN_739 = 6'h23 == _T_224 ? _T_55 : _GEN_738; // @[execute.scala 79:10:@1892.4]
  assign _GEN_740 = 6'h24 == _T_224 ? _T_56 : _GEN_739; // @[execute.scala 79:10:@1892.4]
  assign _GEN_741 = 6'h25 == _T_224 ? _T_57 : _GEN_740; // @[execute.scala 79:10:@1892.4]
  assign _GEN_742 = 6'h26 == _T_224 ? _T_58 : _GEN_741; // @[execute.scala 79:10:@1892.4]
  assign _GEN_743 = 6'h27 == _T_224 ? _T_59 : _GEN_742; // @[execute.scala 79:10:@1892.4]
  assign _GEN_744 = 6'h28 == _T_224 ? _T_60 : _GEN_743; // @[execute.scala 79:10:@1892.4]
  assign _GEN_745 = 6'h29 == _T_224 ? _T_61 : _GEN_744; // @[execute.scala 79:10:@1892.4]
  assign _GEN_746 = 6'h2a == _T_224 ? _T_62 : _GEN_745; // @[execute.scala 79:10:@1892.4]
  assign _GEN_747 = 6'h2b == _T_224 ? _T_63 : _GEN_746; // @[execute.scala 79:10:@1892.4]
  assign _GEN_748 = 6'h2c == _T_224 ? _T_64 : _GEN_747; // @[execute.scala 79:10:@1892.4]
  assign _GEN_749 = 6'h2d == _T_224 ? _T_65 : _GEN_748; // @[execute.scala 79:10:@1892.4]
  assign _GEN_750 = 6'h2e == _T_224 ? _T_66 : _GEN_749; // @[execute.scala 79:10:@1892.4]
  assign _GEN_751 = 6'h2f == _T_224 ? _T_67 : _GEN_750; // @[execute.scala 79:10:@1892.4]
  assign _GEN_752 = 6'h30 == _T_224 ? _T_68 : _GEN_751; // @[execute.scala 79:10:@1892.4]
  assign _GEN_753 = 6'h31 == _T_224 ? _T_69 : _GEN_752; // @[execute.scala 79:10:@1892.4]
  assign _GEN_754 = 6'h32 == _T_224 ? _T_70 : _GEN_753; // @[execute.scala 79:10:@1892.4]
  assign _GEN_755 = 6'h33 == _T_224 ? _T_71 : _GEN_754; // @[execute.scala 79:10:@1892.4]
  assign _GEN_756 = 6'h34 == _T_224 ? _T_72 : _GEN_755; // @[execute.scala 79:10:@1892.4]
  assign _GEN_757 = 6'h35 == _T_224 ? _T_73 : _GEN_756; // @[execute.scala 79:10:@1892.4]
  assign _GEN_758 = 6'h36 == _T_224 ? _T_74 : _GEN_757; // @[execute.scala 79:10:@1892.4]
  assign _GEN_759 = 6'h37 == _T_224 ? _T_75 : _GEN_758; // @[execute.scala 79:10:@1892.4]
  assign _GEN_760 = 6'h38 == _T_224 ? _T_76 : _GEN_759; // @[execute.scala 79:10:@1892.4]
  assign _GEN_761 = 6'h39 == _T_224 ? _T_77 : _GEN_760; // @[execute.scala 79:10:@1892.4]
  assign _GEN_762 = 6'h3a == _T_224 ? _T_78 : _GEN_761; // @[execute.scala 79:10:@1892.4]
  assign _GEN_763 = 6'h3b == _T_224 ? _T_79 : _GEN_762; // @[execute.scala 79:10:@1892.4]
  assign _GEN_764 = 6'h3c == _T_224 ? _T_80 : _GEN_763; // @[execute.scala 79:10:@1892.4]
  assign _GEN_765 = 6'h3d == _T_224 ? _T_81 : _GEN_764; // @[execute.scala 79:10:@1892.4]
  assign _GEN_766 = 6'h3e == _T_224 ? _T_82 : _GEN_765; // @[execute.scala 79:10:@1892.4]
  assign _GEN_767 = 6'h3f == _T_224 ? _T_83 : _GEN_766; // @[execute.scala 79:10:@1892.4]
  assign _T_226 = _T_216 ? _GEN_703 : _GEN_767; // @[execute.scala 79:10:@1892.4]
  assign _T_228 = io_amount < 6'h3a; // @[execute.scala 79:15:@1893.4]
  assign _T_230 = io_amount - 6'h3a; // @[execute.scala 79:37:@1894.4]
  assign _T_231 = $unsigned(_T_230); // @[execute.scala 79:37:@1895.4]
  assign _T_232 = _T_231[5:0]; // @[execute.scala 79:37:@1896.4]
  assign _T_235 = 6'h6 + io_amount; // @[execute.scala 79:60:@1897.4]
  assign _T_236 = 6'h6 + io_amount; // @[execute.scala 79:60:@1898.4]
  assign _GEN_769 = 6'h1 == _T_232 ? _T_21 : _T_20; // @[execute.scala 79:10:@1899.4]
  assign _GEN_770 = 6'h2 == _T_232 ? _T_22 : _GEN_769; // @[execute.scala 79:10:@1899.4]
  assign _GEN_771 = 6'h3 == _T_232 ? _T_23 : _GEN_770; // @[execute.scala 79:10:@1899.4]
  assign _GEN_772 = 6'h4 == _T_232 ? _T_24 : _GEN_771; // @[execute.scala 79:10:@1899.4]
  assign _GEN_773 = 6'h5 == _T_232 ? _T_25 : _GEN_772; // @[execute.scala 79:10:@1899.4]
  assign _GEN_774 = 6'h6 == _T_232 ? _T_26 : _GEN_773; // @[execute.scala 79:10:@1899.4]
  assign _GEN_775 = 6'h7 == _T_232 ? _T_27 : _GEN_774; // @[execute.scala 79:10:@1899.4]
  assign _GEN_776 = 6'h8 == _T_232 ? _T_28 : _GEN_775; // @[execute.scala 79:10:@1899.4]
  assign _GEN_777 = 6'h9 == _T_232 ? _T_29 : _GEN_776; // @[execute.scala 79:10:@1899.4]
  assign _GEN_778 = 6'ha == _T_232 ? _T_30 : _GEN_777; // @[execute.scala 79:10:@1899.4]
  assign _GEN_779 = 6'hb == _T_232 ? _T_31 : _GEN_778; // @[execute.scala 79:10:@1899.4]
  assign _GEN_780 = 6'hc == _T_232 ? _T_32 : _GEN_779; // @[execute.scala 79:10:@1899.4]
  assign _GEN_781 = 6'hd == _T_232 ? _T_33 : _GEN_780; // @[execute.scala 79:10:@1899.4]
  assign _GEN_782 = 6'he == _T_232 ? _T_34 : _GEN_781; // @[execute.scala 79:10:@1899.4]
  assign _GEN_783 = 6'hf == _T_232 ? _T_35 : _GEN_782; // @[execute.scala 79:10:@1899.4]
  assign _GEN_784 = 6'h10 == _T_232 ? _T_36 : _GEN_783; // @[execute.scala 79:10:@1899.4]
  assign _GEN_785 = 6'h11 == _T_232 ? _T_37 : _GEN_784; // @[execute.scala 79:10:@1899.4]
  assign _GEN_786 = 6'h12 == _T_232 ? _T_38 : _GEN_785; // @[execute.scala 79:10:@1899.4]
  assign _GEN_787 = 6'h13 == _T_232 ? _T_39 : _GEN_786; // @[execute.scala 79:10:@1899.4]
  assign _GEN_788 = 6'h14 == _T_232 ? _T_40 : _GEN_787; // @[execute.scala 79:10:@1899.4]
  assign _GEN_789 = 6'h15 == _T_232 ? _T_41 : _GEN_788; // @[execute.scala 79:10:@1899.4]
  assign _GEN_790 = 6'h16 == _T_232 ? _T_42 : _GEN_789; // @[execute.scala 79:10:@1899.4]
  assign _GEN_791 = 6'h17 == _T_232 ? _T_43 : _GEN_790; // @[execute.scala 79:10:@1899.4]
  assign _GEN_792 = 6'h18 == _T_232 ? _T_44 : _GEN_791; // @[execute.scala 79:10:@1899.4]
  assign _GEN_793 = 6'h19 == _T_232 ? _T_45 : _GEN_792; // @[execute.scala 79:10:@1899.4]
  assign _GEN_794 = 6'h1a == _T_232 ? _T_46 : _GEN_793; // @[execute.scala 79:10:@1899.4]
  assign _GEN_795 = 6'h1b == _T_232 ? _T_47 : _GEN_794; // @[execute.scala 79:10:@1899.4]
  assign _GEN_796 = 6'h1c == _T_232 ? _T_48 : _GEN_795; // @[execute.scala 79:10:@1899.4]
  assign _GEN_797 = 6'h1d == _T_232 ? _T_49 : _GEN_796; // @[execute.scala 79:10:@1899.4]
  assign _GEN_798 = 6'h1e == _T_232 ? _T_50 : _GEN_797; // @[execute.scala 79:10:@1899.4]
  assign _GEN_799 = 6'h1f == _T_232 ? _T_51 : _GEN_798; // @[execute.scala 79:10:@1899.4]
  assign _GEN_800 = 6'h20 == _T_232 ? _T_52 : _GEN_799; // @[execute.scala 79:10:@1899.4]
  assign _GEN_801 = 6'h21 == _T_232 ? _T_53 : _GEN_800; // @[execute.scala 79:10:@1899.4]
  assign _GEN_802 = 6'h22 == _T_232 ? _T_54 : _GEN_801; // @[execute.scala 79:10:@1899.4]
  assign _GEN_803 = 6'h23 == _T_232 ? _T_55 : _GEN_802; // @[execute.scala 79:10:@1899.4]
  assign _GEN_804 = 6'h24 == _T_232 ? _T_56 : _GEN_803; // @[execute.scala 79:10:@1899.4]
  assign _GEN_805 = 6'h25 == _T_232 ? _T_57 : _GEN_804; // @[execute.scala 79:10:@1899.4]
  assign _GEN_806 = 6'h26 == _T_232 ? _T_58 : _GEN_805; // @[execute.scala 79:10:@1899.4]
  assign _GEN_807 = 6'h27 == _T_232 ? _T_59 : _GEN_806; // @[execute.scala 79:10:@1899.4]
  assign _GEN_808 = 6'h28 == _T_232 ? _T_60 : _GEN_807; // @[execute.scala 79:10:@1899.4]
  assign _GEN_809 = 6'h29 == _T_232 ? _T_61 : _GEN_808; // @[execute.scala 79:10:@1899.4]
  assign _GEN_810 = 6'h2a == _T_232 ? _T_62 : _GEN_809; // @[execute.scala 79:10:@1899.4]
  assign _GEN_811 = 6'h2b == _T_232 ? _T_63 : _GEN_810; // @[execute.scala 79:10:@1899.4]
  assign _GEN_812 = 6'h2c == _T_232 ? _T_64 : _GEN_811; // @[execute.scala 79:10:@1899.4]
  assign _GEN_813 = 6'h2d == _T_232 ? _T_65 : _GEN_812; // @[execute.scala 79:10:@1899.4]
  assign _GEN_814 = 6'h2e == _T_232 ? _T_66 : _GEN_813; // @[execute.scala 79:10:@1899.4]
  assign _GEN_815 = 6'h2f == _T_232 ? _T_67 : _GEN_814; // @[execute.scala 79:10:@1899.4]
  assign _GEN_816 = 6'h30 == _T_232 ? _T_68 : _GEN_815; // @[execute.scala 79:10:@1899.4]
  assign _GEN_817 = 6'h31 == _T_232 ? _T_69 : _GEN_816; // @[execute.scala 79:10:@1899.4]
  assign _GEN_818 = 6'h32 == _T_232 ? _T_70 : _GEN_817; // @[execute.scala 79:10:@1899.4]
  assign _GEN_819 = 6'h33 == _T_232 ? _T_71 : _GEN_818; // @[execute.scala 79:10:@1899.4]
  assign _GEN_820 = 6'h34 == _T_232 ? _T_72 : _GEN_819; // @[execute.scala 79:10:@1899.4]
  assign _GEN_821 = 6'h35 == _T_232 ? _T_73 : _GEN_820; // @[execute.scala 79:10:@1899.4]
  assign _GEN_822 = 6'h36 == _T_232 ? _T_74 : _GEN_821; // @[execute.scala 79:10:@1899.4]
  assign _GEN_823 = 6'h37 == _T_232 ? _T_75 : _GEN_822; // @[execute.scala 79:10:@1899.4]
  assign _GEN_824 = 6'h38 == _T_232 ? _T_76 : _GEN_823; // @[execute.scala 79:10:@1899.4]
  assign _GEN_825 = 6'h39 == _T_232 ? _T_77 : _GEN_824; // @[execute.scala 79:10:@1899.4]
  assign _GEN_826 = 6'h3a == _T_232 ? _T_78 : _GEN_825; // @[execute.scala 79:10:@1899.4]
  assign _GEN_827 = 6'h3b == _T_232 ? _T_79 : _GEN_826; // @[execute.scala 79:10:@1899.4]
  assign _GEN_828 = 6'h3c == _T_232 ? _T_80 : _GEN_827; // @[execute.scala 79:10:@1899.4]
  assign _GEN_829 = 6'h3d == _T_232 ? _T_81 : _GEN_828; // @[execute.scala 79:10:@1899.4]
  assign _GEN_830 = 6'h3e == _T_232 ? _T_82 : _GEN_829; // @[execute.scala 79:10:@1899.4]
  assign _GEN_831 = 6'h3f == _T_232 ? _T_83 : _GEN_830; // @[execute.scala 79:10:@1899.4]
  assign _GEN_833 = 6'h1 == _T_236 ? _T_21 : _T_20; // @[execute.scala 79:10:@1899.4]
  assign _GEN_834 = 6'h2 == _T_236 ? _T_22 : _GEN_833; // @[execute.scala 79:10:@1899.4]
  assign _GEN_835 = 6'h3 == _T_236 ? _T_23 : _GEN_834; // @[execute.scala 79:10:@1899.4]
  assign _GEN_836 = 6'h4 == _T_236 ? _T_24 : _GEN_835; // @[execute.scala 79:10:@1899.4]
  assign _GEN_837 = 6'h5 == _T_236 ? _T_25 : _GEN_836; // @[execute.scala 79:10:@1899.4]
  assign _GEN_838 = 6'h6 == _T_236 ? _T_26 : _GEN_837; // @[execute.scala 79:10:@1899.4]
  assign _GEN_839 = 6'h7 == _T_236 ? _T_27 : _GEN_838; // @[execute.scala 79:10:@1899.4]
  assign _GEN_840 = 6'h8 == _T_236 ? _T_28 : _GEN_839; // @[execute.scala 79:10:@1899.4]
  assign _GEN_841 = 6'h9 == _T_236 ? _T_29 : _GEN_840; // @[execute.scala 79:10:@1899.4]
  assign _GEN_842 = 6'ha == _T_236 ? _T_30 : _GEN_841; // @[execute.scala 79:10:@1899.4]
  assign _GEN_843 = 6'hb == _T_236 ? _T_31 : _GEN_842; // @[execute.scala 79:10:@1899.4]
  assign _GEN_844 = 6'hc == _T_236 ? _T_32 : _GEN_843; // @[execute.scala 79:10:@1899.4]
  assign _GEN_845 = 6'hd == _T_236 ? _T_33 : _GEN_844; // @[execute.scala 79:10:@1899.4]
  assign _GEN_846 = 6'he == _T_236 ? _T_34 : _GEN_845; // @[execute.scala 79:10:@1899.4]
  assign _GEN_847 = 6'hf == _T_236 ? _T_35 : _GEN_846; // @[execute.scala 79:10:@1899.4]
  assign _GEN_848 = 6'h10 == _T_236 ? _T_36 : _GEN_847; // @[execute.scala 79:10:@1899.4]
  assign _GEN_849 = 6'h11 == _T_236 ? _T_37 : _GEN_848; // @[execute.scala 79:10:@1899.4]
  assign _GEN_850 = 6'h12 == _T_236 ? _T_38 : _GEN_849; // @[execute.scala 79:10:@1899.4]
  assign _GEN_851 = 6'h13 == _T_236 ? _T_39 : _GEN_850; // @[execute.scala 79:10:@1899.4]
  assign _GEN_852 = 6'h14 == _T_236 ? _T_40 : _GEN_851; // @[execute.scala 79:10:@1899.4]
  assign _GEN_853 = 6'h15 == _T_236 ? _T_41 : _GEN_852; // @[execute.scala 79:10:@1899.4]
  assign _GEN_854 = 6'h16 == _T_236 ? _T_42 : _GEN_853; // @[execute.scala 79:10:@1899.4]
  assign _GEN_855 = 6'h17 == _T_236 ? _T_43 : _GEN_854; // @[execute.scala 79:10:@1899.4]
  assign _GEN_856 = 6'h18 == _T_236 ? _T_44 : _GEN_855; // @[execute.scala 79:10:@1899.4]
  assign _GEN_857 = 6'h19 == _T_236 ? _T_45 : _GEN_856; // @[execute.scala 79:10:@1899.4]
  assign _GEN_858 = 6'h1a == _T_236 ? _T_46 : _GEN_857; // @[execute.scala 79:10:@1899.4]
  assign _GEN_859 = 6'h1b == _T_236 ? _T_47 : _GEN_858; // @[execute.scala 79:10:@1899.4]
  assign _GEN_860 = 6'h1c == _T_236 ? _T_48 : _GEN_859; // @[execute.scala 79:10:@1899.4]
  assign _GEN_861 = 6'h1d == _T_236 ? _T_49 : _GEN_860; // @[execute.scala 79:10:@1899.4]
  assign _GEN_862 = 6'h1e == _T_236 ? _T_50 : _GEN_861; // @[execute.scala 79:10:@1899.4]
  assign _GEN_863 = 6'h1f == _T_236 ? _T_51 : _GEN_862; // @[execute.scala 79:10:@1899.4]
  assign _GEN_864 = 6'h20 == _T_236 ? _T_52 : _GEN_863; // @[execute.scala 79:10:@1899.4]
  assign _GEN_865 = 6'h21 == _T_236 ? _T_53 : _GEN_864; // @[execute.scala 79:10:@1899.4]
  assign _GEN_866 = 6'h22 == _T_236 ? _T_54 : _GEN_865; // @[execute.scala 79:10:@1899.4]
  assign _GEN_867 = 6'h23 == _T_236 ? _T_55 : _GEN_866; // @[execute.scala 79:10:@1899.4]
  assign _GEN_868 = 6'h24 == _T_236 ? _T_56 : _GEN_867; // @[execute.scala 79:10:@1899.4]
  assign _GEN_869 = 6'h25 == _T_236 ? _T_57 : _GEN_868; // @[execute.scala 79:10:@1899.4]
  assign _GEN_870 = 6'h26 == _T_236 ? _T_58 : _GEN_869; // @[execute.scala 79:10:@1899.4]
  assign _GEN_871 = 6'h27 == _T_236 ? _T_59 : _GEN_870; // @[execute.scala 79:10:@1899.4]
  assign _GEN_872 = 6'h28 == _T_236 ? _T_60 : _GEN_871; // @[execute.scala 79:10:@1899.4]
  assign _GEN_873 = 6'h29 == _T_236 ? _T_61 : _GEN_872; // @[execute.scala 79:10:@1899.4]
  assign _GEN_874 = 6'h2a == _T_236 ? _T_62 : _GEN_873; // @[execute.scala 79:10:@1899.4]
  assign _GEN_875 = 6'h2b == _T_236 ? _T_63 : _GEN_874; // @[execute.scala 79:10:@1899.4]
  assign _GEN_876 = 6'h2c == _T_236 ? _T_64 : _GEN_875; // @[execute.scala 79:10:@1899.4]
  assign _GEN_877 = 6'h2d == _T_236 ? _T_65 : _GEN_876; // @[execute.scala 79:10:@1899.4]
  assign _GEN_878 = 6'h2e == _T_236 ? _T_66 : _GEN_877; // @[execute.scala 79:10:@1899.4]
  assign _GEN_879 = 6'h2f == _T_236 ? _T_67 : _GEN_878; // @[execute.scala 79:10:@1899.4]
  assign _GEN_880 = 6'h30 == _T_236 ? _T_68 : _GEN_879; // @[execute.scala 79:10:@1899.4]
  assign _GEN_881 = 6'h31 == _T_236 ? _T_69 : _GEN_880; // @[execute.scala 79:10:@1899.4]
  assign _GEN_882 = 6'h32 == _T_236 ? _T_70 : _GEN_881; // @[execute.scala 79:10:@1899.4]
  assign _GEN_883 = 6'h33 == _T_236 ? _T_71 : _GEN_882; // @[execute.scala 79:10:@1899.4]
  assign _GEN_884 = 6'h34 == _T_236 ? _T_72 : _GEN_883; // @[execute.scala 79:10:@1899.4]
  assign _GEN_885 = 6'h35 == _T_236 ? _T_73 : _GEN_884; // @[execute.scala 79:10:@1899.4]
  assign _GEN_886 = 6'h36 == _T_236 ? _T_74 : _GEN_885; // @[execute.scala 79:10:@1899.4]
  assign _GEN_887 = 6'h37 == _T_236 ? _T_75 : _GEN_886; // @[execute.scala 79:10:@1899.4]
  assign _GEN_888 = 6'h38 == _T_236 ? _T_76 : _GEN_887; // @[execute.scala 79:10:@1899.4]
  assign _GEN_889 = 6'h39 == _T_236 ? _T_77 : _GEN_888; // @[execute.scala 79:10:@1899.4]
  assign _GEN_890 = 6'h3a == _T_236 ? _T_78 : _GEN_889; // @[execute.scala 79:10:@1899.4]
  assign _GEN_891 = 6'h3b == _T_236 ? _T_79 : _GEN_890; // @[execute.scala 79:10:@1899.4]
  assign _GEN_892 = 6'h3c == _T_236 ? _T_80 : _GEN_891; // @[execute.scala 79:10:@1899.4]
  assign _GEN_893 = 6'h3d == _T_236 ? _T_81 : _GEN_892; // @[execute.scala 79:10:@1899.4]
  assign _GEN_894 = 6'h3e == _T_236 ? _T_82 : _GEN_893; // @[execute.scala 79:10:@1899.4]
  assign _GEN_895 = 6'h3f == _T_236 ? _T_83 : _GEN_894; // @[execute.scala 79:10:@1899.4]
  assign _T_238 = _T_228 ? _GEN_831 : _GEN_895; // @[execute.scala 79:10:@1899.4]
  assign _T_240 = io_amount < 6'h39; // @[execute.scala 79:15:@1900.4]
  assign _T_242 = io_amount - 6'h39; // @[execute.scala 79:37:@1901.4]
  assign _T_243 = $unsigned(_T_242); // @[execute.scala 79:37:@1902.4]
  assign _T_244 = _T_243[5:0]; // @[execute.scala 79:37:@1903.4]
  assign _T_247 = 6'h7 + io_amount; // @[execute.scala 79:60:@1904.4]
  assign _T_248 = 6'h7 + io_amount; // @[execute.scala 79:60:@1905.4]
  assign _GEN_897 = 6'h1 == _T_244 ? _T_21 : _T_20; // @[execute.scala 79:10:@1906.4]
  assign _GEN_898 = 6'h2 == _T_244 ? _T_22 : _GEN_897; // @[execute.scala 79:10:@1906.4]
  assign _GEN_899 = 6'h3 == _T_244 ? _T_23 : _GEN_898; // @[execute.scala 79:10:@1906.4]
  assign _GEN_900 = 6'h4 == _T_244 ? _T_24 : _GEN_899; // @[execute.scala 79:10:@1906.4]
  assign _GEN_901 = 6'h5 == _T_244 ? _T_25 : _GEN_900; // @[execute.scala 79:10:@1906.4]
  assign _GEN_902 = 6'h6 == _T_244 ? _T_26 : _GEN_901; // @[execute.scala 79:10:@1906.4]
  assign _GEN_903 = 6'h7 == _T_244 ? _T_27 : _GEN_902; // @[execute.scala 79:10:@1906.4]
  assign _GEN_904 = 6'h8 == _T_244 ? _T_28 : _GEN_903; // @[execute.scala 79:10:@1906.4]
  assign _GEN_905 = 6'h9 == _T_244 ? _T_29 : _GEN_904; // @[execute.scala 79:10:@1906.4]
  assign _GEN_906 = 6'ha == _T_244 ? _T_30 : _GEN_905; // @[execute.scala 79:10:@1906.4]
  assign _GEN_907 = 6'hb == _T_244 ? _T_31 : _GEN_906; // @[execute.scala 79:10:@1906.4]
  assign _GEN_908 = 6'hc == _T_244 ? _T_32 : _GEN_907; // @[execute.scala 79:10:@1906.4]
  assign _GEN_909 = 6'hd == _T_244 ? _T_33 : _GEN_908; // @[execute.scala 79:10:@1906.4]
  assign _GEN_910 = 6'he == _T_244 ? _T_34 : _GEN_909; // @[execute.scala 79:10:@1906.4]
  assign _GEN_911 = 6'hf == _T_244 ? _T_35 : _GEN_910; // @[execute.scala 79:10:@1906.4]
  assign _GEN_912 = 6'h10 == _T_244 ? _T_36 : _GEN_911; // @[execute.scala 79:10:@1906.4]
  assign _GEN_913 = 6'h11 == _T_244 ? _T_37 : _GEN_912; // @[execute.scala 79:10:@1906.4]
  assign _GEN_914 = 6'h12 == _T_244 ? _T_38 : _GEN_913; // @[execute.scala 79:10:@1906.4]
  assign _GEN_915 = 6'h13 == _T_244 ? _T_39 : _GEN_914; // @[execute.scala 79:10:@1906.4]
  assign _GEN_916 = 6'h14 == _T_244 ? _T_40 : _GEN_915; // @[execute.scala 79:10:@1906.4]
  assign _GEN_917 = 6'h15 == _T_244 ? _T_41 : _GEN_916; // @[execute.scala 79:10:@1906.4]
  assign _GEN_918 = 6'h16 == _T_244 ? _T_42 : _GEN_917; // @[execute.scala 79:10:@1906.4]
  assign _GEN_919 = 6'h17 == _T_244 ? _T_43 : _GEN_918; // @[execute.scala 79:10:@1906.4]
  assign _GEN_920 = 6'h18 == _T_244 ? _T_44 : _GEN_919; // @[execute.scala 79:10:@1906.4]
  assign _GEN_921 = 6'h19 == _T_244 ? _T_45 : _GEN_920; // @[execute.scala 79:10:@1906.4]
  assign _GEN_922 = 6'h1a == _T_244 ? _T_46 : _GEN_921; // @[execute.scala 79:10:@1906.4]
  assign _GEN_923 = 6'h1b == _T_244 ? _T_47 : _GEN_922; // @[execute.scala 79:10:@1906.4]
  assign _GEN_924 = 6'h1c == _T_244 ? _T_48 : _GEN_923; // @[execute.scala 79:10:@1906.4]
  assign _GEN_925 = 6'h1d == _T_244 ? _T_49 : _GEN_924; // @[execute.scala 79:10:@1906.4]
  assign _GEN_926 = 6'h1e == _T_244 ? _T_50 : _GEN_925; // @[execute.scala 79:10:@1906.4]
  assign _GEN_927 = 6'h1f == _T_244 ? _T_51 : _GEN_926; // @[execute.scala 79:10:@1906.4]
  assign _GEN_928 = 6'h20 == _T_244 ? _T_52 : _GEN_927; // @[execute.scala 79:10:@1906.4]
  assign _GEN_929 = 6'h21 == _T_244 ? _T_53 : _GEN_928; // @[execute.scala 79:10:@1906.4]
  assign _GEN_930 = 6'h22 == _T_244 ? _T_54 : _GEN_929; // @[execute.scala 79:10:@1906.4]
  assign _GEN_931 = 6'h23 == _T_244 ? _T_55 : _GEN_930; // @[execute.scala 79:10:@1906.4]
  assign _GEN_932 = 6'h24 == _T_244 ? _T_56 : _GEN_931; // @[execute.scala 79:10:@1906.4]
  assign _GEN_933 = 6'h25 == _T_244 ? _T_57 : _GEN_932; // @[execute.scala 79:10:@1906.4]
  assign _GEN_934 = 6'h26 == _T_244 ? _T_58 : _GEN_933; // @[execute.scala 79:10:@1906.4]
  assign _GEN_935 = 6'h27 == _T_244 ? _T_59 : _GEN_934; // @[execute.scala 79:10:@1906.4]
  assign _GEN_936 = 6'h28 == _T_244 ? _T_60 : _GEN_935; // @[execute.scala 79:10:@1906.4]
  assign _GEN_937 = 6'h29 == _T_244 ? _T_61 : _GEN_936; // @[execute.scala 79:10:@1906.4]
  assign _GEN_938 = 6'h2a == _T_244 ? _T_62 : _GEN_937; // @[execute.scala 79:10:@1906.4]
  assign _GEN_939 = 6'h2b == _T_244 ? _T_63 : _GEN_938; // @[execute.scala 79:10:@1906.4]
  assign _GEN_940 = 6'h2c == _T_244 ? _T_64 : _GEN_939; // @[execute.scala 79:10:@1906.4]
  assign _GEN_941 = 6'h2d == _T_244 ? _T_65 : _GEN_940; // @[execute.scala 79:10:@1906.4]
  assign _GEN_942 = 6'h2e == _T_244 ? _T_66 : _GEN_941; // @[execute.scala 79:10:@1906.4]
  assign _GEN_943 = 6'h2f == _T_244 ? _T_67 : _GEN_942; // @[execute.scala 79:10:@1906.4]
  assign _GEN_944 = 6'h30 == _T_244 ? _T_68 : _GEN_943; // @[execute.scala 79:10:@1906.4]
  assign _GEN_945 = 6'h31 == _T_244 ? _T_69 : _GEN_944; // @[execute.scala 79:10:@1906.4]
  assign _GEN_946 = 6'h32 == _T_244 ? _T_70 : _GEN_945; // @[execute.scala 79:10:@1906.4]
  assign _GEN_947 = 6'h33 == _T_244 ? _T_71 : _GEN_946; // @[execute.scala 79:10:@1906.4]
  assign _GEN_948 = 6'h34 == _T_244 ? _T_72 : _GEN_947; // @[execute.scala 79:10:@1906.4]
  assign _GEN_949 = 6'h35 == _T_244 ? _T_73 : _GEN_948; // @[execute.scala 79:10:@1906.4]
  assign _GEN_950 = 6'h36 == _T_244 ? _T_74 : _GEN_949; // @[execute.scala 79:10:@1906.4]
  assign _GEN_951 = 6'h37 == _T_244 ? _T_75 : _GEN_950; // @[execute.scala 79:10:@1906.4]
  assign _GEN_952 = 6'h38 == _T_244 ? _T_76 : _GEN_951; // @[execute.scala 79:10:@1906.4]
  assign _GEN_953 = 6'h39 == _T_244 ? _T_77 : _GEN_952; // @[execute.scala 79:10:@1906.4]
  assign _GEN_954 = 6'h3a == _T_244 ? _T_78 : _GEN_953; // @[execute.scala 79:10:@1906.4]
  assign _GEN_955 = 6'h3b == _T_244 ? _T_79 : _GEN_954; // @[execute.scala 79:10:@1906.4]
  assign _GEN_956 = 6'h3c == _T_244 ? _T_80 : _GEN_955; // @[execute.scala 79:10:@1906.4]
  assign _GEN_957 = 6'h3d == _T_244 ? _T_81 : _GEN_956; // @[execute.scala 79:10:@1906.4]
  assign _GEN_958 = 6'h3e == _T_244 ? _T_82 : _GEN_957; // @[execute.scala 79:10:@1906.4]
  assign _GEN_959 = 6'h3f == _T_244 ? _T_83 : _GEN_958; // @[execute.scala 79:10:@1906.4]
  assign _GEN_961 = 6'h1 == _T_248 ? _T_21 : _T_20; // @[execute.scala 79:10:@1906.4]
  assign _GEN_962 = 6'h2 == _T_248 ? _T_22 : _GEN_961; // @[execute.scala 79:10:@1906.4]
  assign _GEN_963 = 6'h3 == _T_248 ? _T_23 : _GEN_962; // @[execute.scala 79:10:@1906.4]
  assign _GEN_964 = 6'h4 == _T_248 ? _T_24 : _GEN_963; // @[execute.scala 79:10:@1906.4]
  assign _GEN_965 = 6'h5 == _T_248 ? _T_25 : _GEN_964; // @[execute.scala 79:10:@1906.4]
  assign _GEN_966 = 6'h6 == _T_248 ? _T_26 : _GEN_965; // @[execute.scala 79:10:@1906.4]
  assign _GEN_967 = 6'h7 == _T_248 ? _T_27 : _GEN_966; // @[execute.scala 79:10:@1906.4]
  assign _GEN_968 = 6'h8 == _T_248 ? _T_28 : _GEN_967; // @[execute.scala 79:10:@1906.4]
  assign _GEN_969 = 6'h9 == _T_248 ? _T_29 : _GEN_968; // @[execute.scala 79:10:@1906.4]
  assign _GEN_970 = 6'ha == _T_248 ? _T_30 : _GEN_969; // @[execute.scala 79:10:@1906.4]
  assign _GEN_971 = 6'hb == _T_248 ? _T_31 : _GEN_970; // @[execute.scala 79:10:@1906.4]
  assign _GEN_972 = 6'hc == _T_248 ? _T_32 : _GEN_971; // @[execute.scala 79:10:@1906.4]
  assign _GEN_973 = 6'hd == _T_248 ? _T_33 : _GEN_972; // @[execute.scala 79:10:@1906.4]
  assign _GEN_974 = 6'he == _T_248 ? _T_34 : _GEN_973; // @[execute.scala 79:10:@1906.4]
  assign _GEN_975 = 6'hf == _T_248 ? _T_35 : _GEN_974; // @[execute.scala 79:10:@1906.4]
  assign _GEN_976 = 6'h10 == _T_248 ? _T_36 : _GEN_975; // @[execute.scala 79:10:@1906.4]
  assign _GEN_977 = 6'h11 == _T_248 ? _T_37 : _GEN_976; // @[execute.scala 79:10:@1906.4]
  assign _GEN_978 = 6'h12 == _T_248 ? _T_38 : _GEN_977; // @[execute.scala 79:10:@1906.4]
  assign _GEN_979 = 6'h13 == _T_248 ? _T_39 : _GEN_978; // @[execute.scala 79:10:@1906.4]
  assign _GEN_980 = 6'h14 == _T_248 ? _T_40 : _GEN_979; // @[execute.scala 79:10:@1906.4]
  assign _GEN_981 = 6'h15 == _T_248 ? _T_41 : _GEN_980; // @[execute.scala 79:10:@1906.4]
  assign _GEN_982 = 6'h16 == _T_248 ? _T_42 : _GEN_981; // @[execute.scala 79:10:@1906.4]
  assign _GEN_983 = 6'h17 == _T_248 ? _T_43 : _GEN_982; // @[execute.scala 79:10:@1906.4]
  assign _GEN_984 = 6'h18 == _T_248 ? _T_44 : _GEN_983; // @[execute.scala 79:10:@1906.4]
  assign _GEN_985 = 6'h19 == _T_248 ? _T_45 : _GEN_984; // @[execute.scala 79:10:@1906.4]
  assign _GEN_986 = 6'h1a == _T_248 ? _T_46 : _GEN_985; // @[execute.scala 79:10:@1906.4]
  assign _GEN_987 = 6'h1b == _T_248 ? _T_47 : _GEN_986; // @[execute.scala 79:10:@1906.4]
  assign _GEN_988 = 6'h1c == _T_248 ? _T_48 : _GEN_987; // @[execute.scala 79:10:@1906.4]
  assign _GEN_989 = 6'h1d == _T_248 ? _T_49 : _GEN_988; // @[execute.scala 79:10:@1906.4]
  assign _GEN_990 = 6'h1e == _T_248 ? _T_50 : _GEN_989; // @[execute.scala 79:10:@1906.4]
  assign _GEN_991 = 6'h1f == _T_248 ? _T_51 : _GEN_990; // @[execute.scala 79:10:@1906.4]
  assign _GEN_992 = 6'h20 == _T_248 ? _T_52 : _GEN_991; // @[execute.scala 79:10:@1906.4]
  assign _GEN_993 = 6'h21 == _T_248 ? _T_53 : _GEN_992; // @[execute.scala 79:10:@1906.4]
  assign _GEN_994 = 6'h22 == _T_248 ? _T_54 : _GEN_993; // @[execute.scala 79:10:@1906.4]
  assign _GEN_995 = 6'h23 == _T_248 ? _T_55 : _GEN_994; // @[execute.scala 79:10:@1906.4]
  assign _GEN_996 = 6'h24 == _T_248 ? _T_56 : _GEN_995; // @[execute.scala 79:10:@1906.4]
  assign _GEN_997 = 6'h25 == _T_248 ? _T_57 : _GEN_996; // @[execute.scala 79:10:@1906.4]
  assign _GEN_998 = 6'h26 == _T_248 ? _T_58 : _GEN_997; // @[execute.scala 79:10:@1906.4]
  assign _GEN_999 = 6'h27 == _T_248 ? _T_59 : _GEN_998; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1000 = 6'h28 == _T_248 ? _T_60 : _GEN_999; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1001 = 6'h29 == _T_248 ? _T_61 : _GEN_1000; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1002 = 6'h2a == _T_248 ? _T_62 : _GEN_1001; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1003 = 6'h2b == _T_248 ? _T_63 : _GEN_1002; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1004 = 6'h2c == _T_248 ? _T_64 : _GEN_1003; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1005 = 6'h2d == _T_248 ? _T_65 : _GEN_1004; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1006 = 6'h2e == _T_248 ? _T_66 : _GEN_1005; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1007 = 6'h2f == _T_248 ? _T_67 : _GEN_1006; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1008 = 6'h30 == _T_248 ? _T_68 : _GEN_1007; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1009 = 6'h31 == _T_248 ? _T_69 : _GEN_1008; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1010 = 6'h32 == _T_248 ? _T_70 : _GEN_1009; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1011 = 6'h33 == _T_248 ? _T_71 : _GEN_1010; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1012 = 6'h34 == _T_248 ? _T_72 : _GEN_1011; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1013 = 6'h35 == _T_248 ? _T_73 : _GEN_1012; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1014 = 6'h36 == _T_248 ? _T_74 : _GEN_1013; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1015 = 6'h37 == _T_248 ? _T_75 : _GEN_1014; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1016 = 6'h38 == _T_248 ? _T_76 : _GEN_1015; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1017 = 6'h39 == _T_248 ? _T_77 : _GEN_1016; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1018 = 6'h3a == _T_248 ? _T_78 : _GEN_1017; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1019 = 6'h3b == _T_248 ? _T_79 : _GEN_1018; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1020 = 6'h3c == _T_248 ? _T_80 : _GEN_1019; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1021 = 6'h3d == _T_248 ? _T_81 : _GEN_1020; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1022 = 6'h3e == _T_248 ? _T_82 : _GEN_1021; // @[execute.scala 79:10:@1906.4]
  assign _GEN_1023 = 6'h3f == _T_248 ? _T_83 : _GEN_1022; // @[execute.scala 79:10:@1906.4]
  assign _T_250 = _T_240 ? _GEN_959 : _GEN_1023; // @[execute.scala 79:10:@1906.4]
  assign _T_252 = io_amount < 6'h38; // @[execute.scala 79:15:@1907.4]
  assign _T_254 = io_amount - 6'h38; // @[execute.scala 79:37:@1908.4]
  assign _T_255 = $unsigned(_T_254); // @[execute.scala 79:37:@1909.4]
  assign _T_256 = _T_255[5:0]; // @[execute.scala 79:37:@1910.4]
  assign _T_259 = 6'h8 + io_amount; // @[execute.scala 79:60:@1911.4]
  assign _T_260 = 6'h8 + io_amount; // @[execute.scala 79:60:@1912.4]
  assign _GEN_1025 = 6'h1 == _T_256 ? _T_21 : _T_20; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1026 = 6'h2 == _T_256 ? _T_22 : _GEN_1025; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1027 = 6'h3 == _T_256 ? _T_23 : _GEN_1026; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1028 = 6'h4 == _T_256 ? _T_24 : _GEN_1027; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1029 = 6'h5 == _T_256 ? _T_25 : _GEN_1028; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1030 = 6'h6 == _T_256 ? _T_26 : _GEN_1029; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1031 = 6'h7 == _T_256 ? _T_27 : _GEN_1030; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1032 = 6'h8 == _T_256 ? _T_28 : _GEN_1031; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1033 = 6'h9 == _T_256 ? _T_29 : _GEN_1032; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1034 = 6'ha == _T_256 ? _T_30 : _GEN_1033; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1035 = 6'hb == _T_256 ? _T_31 : _GEN_1034; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1036 = 6'hc == _T_256 ? _T_32 : _GEN_1035; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1037 = 6'hd == _T_256 ? _T_33 : _GEN_1036; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1038 = 6'he == _T_256 ? _T_34 : _GEN_1037; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1039 = 6'hf == _T_256 ? _T_35 : _GEN_1038; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1040 = 6'h10 == _T_256 ? _T_36 : _GEN_1039; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1041 = 6'h11 == _T_256 ? _T_37 : _GEN_1040; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1042 = 6'h12 == _T_256 ? _T_38 : _GEN_1041; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1043 = 6'h13 == _T_256 ? _T_39 : _GEN_1042; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1044 = 6'h14 == _T_256 ? _T_40 : _GEN_1043; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1045 = 6'h15 == _T_256 ? _T_41 : _GEN_1044; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1046 = 6'h16 == _T_256 ? _T_42 : _GEN_1045; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1047 = 6'h17 == _T_256 ? _T_43 : _GEN_1046; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1048 = 6'h18 == _T_256 ? _T_44 : _GEN_1047; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1049 = 6'h19 == _T_256 ? _T_45 : _GEN_1048; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1050 = 6'h1a == _T_256 ? _T_46 : _GEN_1049; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1051 = 6'h1b == _T_256 ? _T_47 : _GEN_1050; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1052 = 6'h1c == _T_256 ? _T_48 : _GEN_1051; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1053 = 6'h1d == _T_256 ? _T_49 : _GEN_1052; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1054 = 6'h1e == _T_256 ? _T_50 : _GEN_1053; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1055 = 6'h1f == _T_256 ? _T_51 : _GEN_1054; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1056 = 6'h20 == _T_256 ? _T_52 : _GEN_1055; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1057 = 6'h21 == _T_256 ? _T_53 : _GEN_1056; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1058 = 6'h22 == _T_256 ? _T_54 : _GEN_1057; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1059 = 6'h23 == _T_256 ? _T_55 : _GEN_1058; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1060 = 6'h24 == _T_256 ? _T_56 : _GEN_1059; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1061 = 6'h25 == _T_256 ? _T_57 : _GEN_1060; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1062 = 6'h26 == _T_256 ? _T_58 : _GEN_1061; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1063 = 6'h27 == _T_256 ? _T_59 : _GEN_1062; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1064 = 6'h28 == _T_256 ? _T_60 : _GEN_1063; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1065 = 6'h29 == _T_256 ? _T_61 : _GEN_1064; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1066 = 6'h2a == _T_256 ? _T_62 : _GEN_1065; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1067 = 6'h2b == _T_256 ? _T_63 : _GEN_1066; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1068 = 6'h2c == _T_256 ? _T_64 : _GEN_1067; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1069 = 6'h2d == _T_256 ? _T_65 : _GEN_1068; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1070 = 6'h2e == _T_256 ? _T_66 : _GEN_1069; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1071 = 6'h2f == _T_256 ? _T_67 : _GEN_1070; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1072 = 6'h30 == _T_256 ? _T_68 : _GEN_1071; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1073 = 6'h31 == _T_256 ? _T_69 : _GEN_1072; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1074 = 6'h32 == _T_256 ? _T_70 : _GEN_1073; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1075 = 6'h33 == _T_256 ? _T_71 : _GEN_1074; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1076 = 6'h34 == _T_256 ? _T_72 : _GEN_1075; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1077 = 6'h35 == _T_256 ? _T_73 : _GEN_1076; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1078 = 6'h36 == _T_256 ? _T_74 : _GEN_1077; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1079 = 6'h37 == _T_256 ? _T_75 : _GEN_1078; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1080 = 6'h38 == _T_256 ? _T_76 : _GEN_1079; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1081 = 6'h39 == _T_256 ? _T_77 : _GEN_1080; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1082 = 6'h3a == _T_256 ? _T_78 : _GEN_1081; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1083 = 6'h3b == _T_256 ? _T_79 : _GEN_1082; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1084 = 6'h3c == _T_256 ? _T_80 : _GEN_1083; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1085 = 6'h3d == _T_256 ? _T_81 : _GEN_1084; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1086 = 6'h3e == _T_256 ? _T_82 : _GEN_1085; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1087 = 6'h3f == _T_256 ? _T_83 : _GEN_1086; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1089 = 6'h1 == _T_260 ? _T_21 : _T_20; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1090 = 6'h2 == _T_260 ? _T_22 : _GEN_1089; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1091 = 6'h3 == _T_260 ? _T_23 : _GEN_1090; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1092 = 6'h4 == _T_260 ? _T_24 : _GEN_1091; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1093 = 6'h5 == _T_260 ? _T_25 : _GEN_1092; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1094 = 6'h6 == _T_260 ? _T_26 : _GEN_1093; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1095 = 6'h7 == _T_260 ? _T_27 : _GEN_1094; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1096 = 6'h8 == _T_260 ? _T_28 : _GEN_1095; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1097 = 6'h9 == _T_260 ? _T_29 : _GEN_1096; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1098 = 6'ha == _T_260 ? _T_30 : _GEN_1097; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1099 = 6'hb == _T_260 ? _T_31 : _GEN_1098; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1100 = 6'hc == _T_260 ? _T_32 : _GEN_1099; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1101 = 6'hd == _T_260 ? _T_33 : _GEN_1100; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1102 = 6'he == _T_260 ? _T_34 : _GEN_1101; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1103 = 6'hf == _T_260 ? _T_35 : _GEN_1102; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1104 = 6'h10 == _T_260 ? _T_36 : _GEN_1103; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1105 = 6'h11 == _T_260 ? _T_37 : _GEN_1104; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1106 = 6'h12 == _T_260 ? _T_38 : _GEN_1105; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1107 = 6'h13 == _T_260 ? _T_39 : _GEN_1106; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1108 = 6'h14 == _T_260 ? _T_40 : _GEN_1107; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1109 = 6'h15 == _T_260 ? _T_41 : _GEN_1108; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1110 = 6'h16 == _T_260 ? _T_42 : _GEN_1109; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1111 = 6'h17 == _T_260 ? _T_43 : _GEN_1110; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1112 = 6'h18 == _T_260 ? _T_44 : _GEN_1111; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1113 = 6'h19 == _T_260 ? _T_45 : _GEN_1112; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1114 = 6'h1a == _T_260 ? _T_46 : _GEN_1113; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1115 = 6'h1b == _T_260 ? _T_47 : _GEN_1114; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1116 = 6'h1c == _T_260 ? _T_48 : _GEN_1115; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1117 = 6'h1d == _T_260 ? _T_49 : _GEN_1116; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1118 = 6'h1e == _T_260 ? _T_50 : _GEN_1117; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1119 = 6'h1f == _T_260 ? _T_51 : _GEN_1118; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1120 = 6'h20 == _T_260 ? _T_52 : _GEN_1119; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1121 = 6'h21 == _T_260 ? _T_53 : _GEN_1120; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1122 = 6'h22 == _T_260 ? _T_54 : _GEN_1121; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1123 = 6'h23 == _T_260 ? _T_55 : _GEN_1122; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1124 = 6'h24 == _T_260 ? _T_56 : _GEN_1123; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1125 = 6'h25 == _T_260 ? _T_57 : _GEN_1124; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1126 = 6'h26 == _T_260 ? _T_58 : _GEN_1125; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1127 = 6'h27 == _T_260 ? _T_59 : _GEN_1126; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1128 = 6'h28 == _T_260 ? _T_60 : _GEN_1127; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1129 = 6'h29 == _T_260 ? _T_61 : _GEN_1128; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1130 = 6'h2a == _T_260 ? _T_62 : _GEN_1129; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1131 = 6'h2b == _T_260 ? _T_63 : _GEN_1130; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1132 = 6'h2c == _T_260 ? _T_64 : _GEN_1131; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1133 = 6'h2d == _T_260 ? _T_65 : _GEN_1132; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1134 = 6'h2e == _T_260 ? _T_66 : _GEN_1133; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1135 = 6'h2f == _T_260 ? _T_67 : _GEN_1134; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1136 = 6'h30 == _T_260 ? _T_68 : _GEN_1135; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1137 = 6'h31 == _T_260 ? _T_69 : _GEN_1136; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1138 = 6'h32 == _T_260 ? _T_70 : _GEN_1137; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1139 = 6'h33 == _T_260 ? _T_71 : _GEN_1138; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1140 = 6'h34 == _T_260 ? _T_72 : _GEN_1139; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1141 = 6'h35 == _T_260 ? _T_73 : _GEN_1140; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1142 = 6'h36 == _T_260 ? _T_74 : _GEN_1141; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1143 = 6'h37 == _T_260 ? _T_75 : _GEN_1142; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1144 = 6'h38 == _T_260 ? _T_76 : _GEN_1143; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1145 = 6'h39 == _T_260 ? _T_77 : _GEN_1144; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1146 = 6'h3a == _T_260 ? _T_78 : _GEN_1145; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1147 = 6'h3b == _T_260 ? _T_79 : _GEN_1146; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1148 = 6'h3c == _T_260 ? _T_80 : _GEN_1147; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1149 = 6'h3d == _T_260 ? _T_81 : _GEN_1148; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1150 = 6'h3e == _T_260 ? _T_82 : _GEN_1149; // @[execute.scala 79:10:@1913.4]
  assign _GEN_1151 = 6'h3f == _T_260 ? _T_83 : _GEN_1150; // @[execute.scala 79:10:@1913.4]
  assign _T_262 = _T_252 ? _GEN_1087 : _GEN_1151; // @[execute.scala 79:10:@1913.4]
  assign _T_264 = io_amount < 6'h37; // @[execute.scala 79:15:@1914.4]
  assign _T_266 = io_amount - 6'h37; // @[execute.scala 79:37:@1915.4]
  assign _T_267 = $unsigned(_T_266); // @[execute.scala 79:37:@1916.4]
  assign _T_268 = _T_267[5:0]; // @[execute.scala 79:37:@1917.4]
  assign _T_271 = 6'h9 + io_amount; // @[execute.scala 79:60:@1918.4]
  assign _T_272 = 6'h9 + io_amount; // @[execute.scala 79:60:@1919.4]
  assign _GEN_1153 = 6'h1 == _T_268 ? _T_21 : _T_20; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1154 = 6'h2 == _T_268 ? _T_22 : _GEN_1153; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1155 = 6'h3 == _T_268 ? _T_23 : _GEN_1154; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1156 = 6'h4 == _T_268 ? _T_24 : _GEN_1155; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1157 = 6'h5 == _T_268 ? _T_25 : _GEN_1156; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1158 = 6'h6 == _T_268 ? _T_26 : _GEN_1157; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1159 = 6'h7 == _T_268 ? _T_27 : _GEN_1158; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1160 = 6'h8 == _T_268 ? _T_28 : _GEN_1159; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1161 = 6'h9 == _T_268 ? _T_29 : _GEN_1160; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1162 = 6'ha == _T_268 ? _T_30 : _GEN_1161; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1163 = 6'hb == _T_268 ? _T_31 : _GEN_1162; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1164 = 6'hc == _T_268 ? _T_32 : _GEN_1163; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1165 = 6'hd == _T_268 ? _T_33 : _GEN_1164; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1166 = 6'he == _T_268 ? _T_34 : _GEN_1165; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1167 = 6'hf == _T_268 ? _T_35 : _GEN_1166; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1168 = 6'h10 == _T_268 ? _T_36 : _GEN_1167; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1169 = 6'h11 == _T_268 ? _T_37 : _GEN_1168; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1170 = 6'h12 == _T_268 ? _T_38 : _GEN_1169; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1171 = 6'h13 == _T_268 ? _T_39 : _GEN_1170; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1172 = 6'h14 == _T_268 ? _T_40 : _GEN_1171; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1173 = 6'h15 == _T_268 ? _T_41 : _GEN_1172; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1174 = 6'h16 == _T_268 ? _T_42 : _GEN_1173; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1175 = 6'h17 == _T_268 ? _T_43 : _GEN_1174; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1176 = 6'h18 == _T_268 ? _T_44 : _GEN_1175; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1177 = 6'h19 == _T_268 ? _T_45 : _GEN_1176; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1178 = 6'h1a == _T_268 ? _T_46 : _GEN_1177; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1179 = 6'h1b == _T_268 ? _T_47 : _GEN_1178; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1180 = 6'h1c == _T_268 ? _T_48 : _GEN_1179; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1181 = 6'h1d == _T_268 ? _T_49 : _GEN_1180; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1182 = 6'h1e == _T_268 ? _T_50 : _GEN_1181; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1183 = 6'h1f == _T_268 ? _T_51 : _GEN_1182; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1184 = 6'h20 == _T_268 ? _T_52 : _GEN_1183; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1185 = 6'h21 == _T_268 ? _T_53 : _GEN_1184; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1186 = 6'h22 == _T_268 ? _T_54 : _GEN_1185; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1187 = 6'h23 == _T_268 ? _T_55 : _GEN_1186; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1188 = 6'h24 == _T_268 ? _T_56 : _GEN_1187; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1189 = 6'h25 == _T_268 ? _T_57 : _GEN_1188; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1190 = 6'h26 == _T_268 ? _T_58 : _GEN_1189; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1191 = 6'h27 == _T_268 ? _T_59 : _GEN_1190; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1192 = 6'h28 == _T_268 ? _T_60 : _GEN_1191; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1193 = 6'h29 == _T_268 ? _T_61 : _GEN_1192; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1194 = 6'h2a == _T_268 ? _T_62 : _GEN_1193; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1195 = 6'h2b == _T_268 ? _T_63 : _GEN_1194; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1196 = 6'h2c == _T_268 ? _T_64 : _GEN_1195; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1197 = 6'h2d == _T_268 ? _T_65 : _GEN_1196; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1198 = 6'h2e == _T_268 ? _T_66 : _GEN_1197; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1199 = 6'h2f == _T_268 ? _T_67 : _GEN_1198; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1200 = 6'h30 == _T_268 ? _T_68 : _GEN_1199; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1201 = 6'h31 == _T_268 ? _T_69 : _GEN_1200; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1202 = 6'h32 == _T_268 ? _T_70 : _GEN_1201; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1203 = 6'h33 == _T_268 ? _T_71 : _GEN_1202; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1204 = 6'h34 == _T_268 ? _T_72 : _GEN_1203; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1205 = 6'h35 == _T_268 ? _T_73 : _GEN_1204; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1206 = 6'h36 == _T_268 ? _T_74 : _GEN_1205; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1207 = 6'h37 == _T_268 ? _T_75 : _GEN_1206; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1208 = 6'h38 == _T_268 ? _T_76 : _GEN_1207; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1209 = 6'h39 == _T_268 ? _T_77 : _GEN_1208; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1210 = 6'h3a == _T_268 ? _T_78 : _GEN_1209; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1211 = 6'h3b == _T_268 ? _T_79 : _GEN_1210; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1212 = 6'h3c == _T_268 ? _T_80 : _GEN_1211; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1213 = 6'h3d == _T_268 ? _T_81 : _GEN_1212; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1214 = 6'h3e == _T_268 ? _T_82 : _GEN_1213; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1215 = 6'h3f == _T_268 ? _T_83 : _GEN_1214; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1217 = 6'h1 == _T_272 ? _T_21 : _T_20; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1218 = 6'h2 == _T_272 ? _T_22 : _GEN_1217; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1219 = 6'h3 == _T_272 ? _T_23 : _GEN_1218; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1220 = 6'h4 == _T_272 ? _T_24 : _GEN_1219; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1221 = 6'h5 == _T_272 ? _T_25 : _GEN_1220; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1222 = 6'h6 == _T_272 ? _T_26 : _GEN_1221; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1223 = 6'h7 == _T_272 ? _T_27 : _GEN_1222; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1224 = 6'h8 == _T_272 ? _T_28 : _GEN_1223; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1225 = 6'h9 == _T_272 ? _T_29 : _GEN_1224; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1226 = 6'ha == _T_272 ? _T_30 : _GEN_1225; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1227 = 6'hb == _T_272 ? _T_31 : _GEN_1226; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1228 = 6'hc == _T_272 ? _T_32 : _GEN_1227; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1229 = 6'hd == _T_272 ? _T_33 : _GEN_1228; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1230 = 6'he == _T_272 ? _T_34 : _GEN_1229; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1231 = 6'hf == _T_272 ? _T_35 : _GEN_1230; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1232 = 6'h10 == _T_272 ? _T_36 : _GEN_1231; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1233 = 6'h11 == _T_272 ? _T_37 : _GEN_1232; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1234 = 6'h12 == _T_272 ? _T_38 : _GEN_1233; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1235 = 6'h13 == _T_272 ? _T_39 : _GEN_1234; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1236 = 6'h14 == _T_272 ? _T_40 : _GEN_1235; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1237 = 6'h15 == _T_272 ? _T_41 : _GEN_1236; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1238 = 6'h16 == _T_272 ? _T_42 : _GEN_1237; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1239 = 6'h17 == _T_272 ? _T_43 : _GEN_1238; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1240 = 6'h18 == _T_272 ? _T_44 : _GEN_1239; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1241 = 6'h19 == _T_272 ? _T_45 : _GEN_1240; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1242 = 6'h1a == _T_272 ? _T_46 : _GEN_1241; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1243 = 6'h1b == _T_272 ? _T_47 : _GEN_1242; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1244 = 6'h1c == _T_272 ? _T_48 : _GEN_1243; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1245 = 6'h1d == _T_272 ? _T_49 : _GEN_1244; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1246 = 6'h1e == _T_272 ? _T_50 : _GEN_1245; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1247 = 6'h1f == _T_272 ? _T_51 : _GEN_1246; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1248 = 6'h20 == _T_272 ? _T_52 : _GEN_1247; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1249 = 6'h21 == _T_272 ? _T_53 : _GEN_1248; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1250 = 6'h22 == _T_272 ? _T_54 : _GEN_1249; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1251 = 6'h23 == _T_272 ? _T_55 : _GEN_1250; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1252 = 6'h24 == _T_272 ? _T_56 : _GEN_1251; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1253 = 6'h25 == _T_272 ? _T_57 : _GEN_1252; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1254 = 6'h26 == _T_272 ? _T_58 : _GEN_1253; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1255 = 6'h27 == _T_272 ? _T_59 : _GEN_1254; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1256 = 6'h28 == _T_272 ? _T_60 : _GEN_1255; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1257 = 6'h29 == _T_272 ? _T_61 : _GEN_1256; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1258 = 6'h2a == _T_272 ? _T_62 : _GEN_1257; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1259 = 6'h2b == _T_272 ? _T_63 : _GEN_1258; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1260 = 6'h2c == _T_272 ? _T_64 : _GEN_1259; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1261 = 6'h2d == _T_272 ? _T_65 : _GEN_1260; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1262 = 6'h2e == _T_272 ? _T_66 : _GEN_1261; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1263 = 6'h2f == _T_272 ? _T_67 : _GEN_1262; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1264 = 6'h30 == _T_272 ? _T_68 : _GEN_1263; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1265 = 6'h31 == _T_272 ? _T_69 : _GEN_1264; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1266 = 6'h32 == _T_272 ? _T_70 : _GEN_1265; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1267 = 6'h33 == _T_272 ? _T_71 : _GEN_1266; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1268 = 6'h34 == _T_272 ? _T_72 : _GEN_1267; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1269 = 6'h35 == _T_272 ? _T_73 : _GEN_1268; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1270 = 6'h36 == _T_272 ? _T_74 : _GEN_1269; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1271 = 6'h37 == _T_272 ? _T_75 : _GEN_1270; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1272 = 6'h38 == _T_272 ? _T_76 : _GEN_1271; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1273 = 6'h39 == _T_272 ? _T_77 : _GEN_1272; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1274 = 6'h3a == _T_272 ? _T_78 : _GEN_1273; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1275 = 6'h3b == _T_272 ? _T_79 : _GEN_1274; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1276 = 6'h3c == _T_272 ? _T_80 : _GEN_1275; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1277 = 6'h3d == _T_272 ? _T_81 : _GEN_1276; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1278 = 6'h3e == _T_272 ? _T_82 : _GEN_1277; // @[execute.scala 79:10:@1920.4]
  assign _GEN_1279 = 6'h3f == _T_272 ? _T_83 : _GEN_1278; // @[execute.scala 79:10:@1920.4]
  assign _T_274 = _T_264 ? _GEN_1215 : _GEN_1279; // @[execute.scala 79:10:@1920.4]
  assign _T_276 = io_amount < 6'h36; // @[execute.scala 79:15:@1921.4]
  assign _T_278 = io_amount - 6'h36; // @[execute.scala 79:37:@1922.4]
  assign _T_279 = $unsigned(_T_278); // @[execute.scala 79:37:@1923.4]
  assign _T_280 = _T_279[5:0]; // @[execute.scala 79:37:@1924.4]
  assign _T_283 = 6'ha + io_amount; // @[execute.scala 79:60:@1925.4]
  assign _T_284 = 6'ha + io_amount; // @[execute.scala 79:60:@1926.4]
  assign _GEN_1281 = 6'h1 == _T_280 ? _T_21 : _T_20; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1282 = 6'h2 == _T_280 ? _T_22 : _GEN_1281; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1283 = 6'h3 == _T_280 ? _T_23 : _GEN_1282; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1284 = 6'h4 == _T_280 ? _T_24 : _GEN_1283; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1285 = 6'h5 == _T_280 ? _T_25 : _GEN_1284; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1286 = 6'h6 == _T_280 ? _T_26 : _GEN_1285; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1287 = 6'h7 == _T_280 ? _T_27 : _GEN_1286; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1288 = 6'h8 == _T_280 ? _T_28 : _GEN_1287; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1289 = 6'h9 == _T_280 ? _T_29 : _GEN_1288; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1290 = 6'ha == _T_280 ? _T_30 : _GEN_1289; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1291 = 6'hb == _T_280 ? _T_31 : _GEN_1290; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1292 = 6'hc == _T_280 ? _T_32 : _GEN_1291; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1293 = 6'hd == _T_280 ? _T_33 : _GEN_1292; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1294 = 6'he == _T_280 ? _T_34 : _GEN_1293; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1295 = 6'hf == _T_280 ? _T_35 : _GEN_1294; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1296 = 6'h10 == _T_280 ? _T_36 : _GEN_1295; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1297 = 6'h11 == _T_280 ? _T_37 : _GEN_1296; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1298 = 6'h12 == _T_280 ? _T_38 : _GEN_1297; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1299 = 6'h13 == _T_280 ? _T_39 : _GEN_1298; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1300 = 6'h14 == _T_280 ? _T_40 : _GEN_1299; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1301 = 6'h15 == _T_280 ? _T_41 : _GEN_1300; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1302 = 6'h16 == _T_280 ? _T_42 : _GEN_1301; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1303 = 6'h17 == _T_280 ? _T_43 : _GEN_1302; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1304 = 6'h18 == _T_280 ? _T_44 : _GEN_1303; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1305 = 6'h19 == _T_280 ? _T_45 : _GEN_1304; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1306 = 6'h1a == _T_280 ? _T_46 : _GEN_1305; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1307 = 6'h1b == _T_280 ? _T_47 : _GEN_1306; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1308 = 6'h1c == _T_280 ? _T_48 : _GEN_1307; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1309 = 6'h1d == _T_280 ? _T_49 : _GEN_1308; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1310 = 6'h1e == _T_280 ? _T_50 : _GEN_1309; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1311 = 6'h1f == _T_280 ? _T_51 : _GEN_1310; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1312 = 6'h20 == _T_280 ? _T_52 : _GEN_1311; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1313 = 6'h21 == _T_280 ? _T_53 : _GEN_1312; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1314 = 6'h22 == _T_280 ? _T_54 : _GEN_1313; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1315 = 6'h23 == _T_280 ? _T_55 : _GEN_1314; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1316 = 6'h24 == _T_280 ? _T_56 : _GEN_1315; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1317 = 6'h25 == _T_280 ? _T_57 : _GEN_1316; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1318 = 6'h26 == _T_280 ? _T_58 : _GEN_1317; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1319 = 6'h27 == _T_280 ? _T_59 : _GEN_1318; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1320 = 6'h28 == _T_280 ? _T_60 : _GEN_1319; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1321 = 6'h29 == _T_280 ? _T_61 : _GEN_1320; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1322 = 6'h2a == _T_280 ? _T_62 : _GEN_1321; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1323 = 6'h2b == _T_280 ? _T_63 : _GEN_1322; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1324 = 6'h2c == _T_280 ? _T_64 : _GEN_1323; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1325 = 6'h2d == _T_280 ? _T_65 : _GEN_1324; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1326 = 6'h2e == _T_280 ? _T_66 : _GEN_1325; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1327 = 6'h2f == _T_280 ? _T_67 : _GEN_1326; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1328 = 6'h30 == _T_280 ? _T_68 : _GEN_1327; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1329 = 6'h31 == _T_280 ? _T_69 : _GEN_1328; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1330 = 6'h32 == _T_280 ? _T_70 : _GEN_1329; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1331 = 6'h33 == _T_280 ? _T_71 : _GEN_1330; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1332 = 6'h34 == _T_280 ? _T_72 : _GEN_1331; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1333 = 6'h35 == _T_280 ? _T_73 : _GEN_1332; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1334 = 6'h36 == _T_280 ? _T_74 : _GEN_1333; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1335 = 6'h37 == _T_280 ? _T_75 : _GEN_1334; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1336 = 6'h38 == _T_280 ? _T_76 : _GEN_1335; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1337 = 6'h39 == _T_280 ? _T_77 : _GEN_1336; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1338 = 6'h3a == _T_280 ? _T_78 : _GEN_1337; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1339 = 6'h3b == _T_280 ? _T_79 : _GEN_1338; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1340 = 6'h3c == _T_280 ? _T_80 : _GEN_1339; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1341 = 6'h3d == _T_280 ? _T_81 : _GEN_1340; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1342 = 6'h3e == _T_280 ? _T_82 : _GEN_1341; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1343 = 6'h3f == _T_280 ? _T_83 : _GEN_1342; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1345 = 6'h1 == _T_284 ? _T_21 : _T_20; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1346 = 6'h2 == _T_284 ? _T_22 : _GEN_1345; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1347 = 6'h3 == _T_284 ? _T_23 : _GEN_1346; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1348 = 6'h4 == _T_284 ? _T_24 : _GEN_1347; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1349 = 6'h5 == _T_284 ? _T_25 : _GEN_1348; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1350 = 6'h6 == _T_284 ? _T_26 : _GEN_1349; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1351 = 6'h7 == _T_284 ? _T_27 : _GEN_1350; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1352 = 6'h8 == _T_284 ? _T_28 : _GEN_1351; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1353 = 6'h9 == _T_284 ? _T_29 : _GEN_1352; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1354 = 6'ha == _T_284 ? _T_30 : _GEN_1353; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1355 = 6'hb == _T_284 ? _T_31 : _GEN_1354; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1356 = 6'hc == _T_284 ? _T_32 : _GEN_1355; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1357 = 6'hd == _T_284 ? _T_33 : _GEN_1356; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1358 = 6'he == _T_284 ? _T_34 : _GEN_1357; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1359 = 6'hf == _T_284 ? _T_35 : _GEN_1358; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1360 = 6'h10 == _T_284 ? _T_36 : _GEN_1359; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1361 = 6'h11 == _T_284 ? _T_37 : _GEN_1360; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1362 = 6'h12 == _T_284 ? _T_38 : _GEN_1361; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1363 = 6'h13 == _T_284 ? _T_39 : _GEN_1362; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1364 = 6'h14 == _T_284 ? _T_40 : _GEN_1363; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1365 = 6'h15 == _T_284 ? _T_41 : _GEN_1364; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1366 = 6'h16 == _T_284 ? _T_42 : _GEN_1365; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1367 = 6'h17 == _T_284 ? _T_43 : _GEN_1366; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1368 = 6'h18 == _T_284 ? _T_44 : _GEN_1367; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1369 = 6'h19 == _T_284 ? _T_45 : _GEN_1368; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1370 = 6'h1a == _T_284 ? _T_46 : _GEN_1369; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1371 = 6'h1b == _T_284 ? _T_47 : _GEN_1370; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1372 = 6'h1c == _T_284 ? _T_48 : _GEN_1371; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1373 = 6'h1d == _T_284 ? _T_49 : _GEN_1372; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1374 = 6'h1e == _T_284 ? _T_50 : _GEN_1373; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1375 = 6'h1f == _T_284 ? _T_51 : _GEN_1374; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1376 = 6'h20 == _T_284 ? _T_52 : _GEN_1375; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1377 = 6'h21 == _T_284 ? _T_53 : _GEN_1376; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1378 = 6'h22 == _T_284 ? _T_54 : _GEN_1377; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1379 = 6'h23 == _T_284 ? _T_55 : _GEN_1378; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1380 = 6'h24 == _T_284 ? _T_56 : _GEN_1379; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1381 = 6'h25 == _T_284 ? _T_57 : _GEN_1380; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1382 = 6'h26 == _T_284 ? _T_58 : _GEN_1381; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1383 = 6'h27 == _T_284 ? _T_59 : _GEN_1382; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1384 = 6'h28 == _T_284 ? _T_60 : _GEN_1383; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1385 = 6'h29 == _T_284 ? _T_61 : _GEN_1384; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1386 = 6'h2a == _T_284 ? _T_62 : _GEN_1385; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1387 = 6'h2b == _T_284 ? _T_63 : _GEN_1386; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1388 = 6'h2c == _T_284 ? _T_64 : _GEN_1387; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1389 = 6'h2d == _T_284 ? _T_65 : _GEN_1388; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1390 = 6'h2e == _T_284 ? _T_66 : _GEN_1389; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1391 = 6'h2f == _T_284 ? _T_67 : _GEN_1390; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1392 = 6'h30 == _T_284 ? _T_68 : _GEN_1391; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1393 = 6'h31 == _T_284 ? _T_69 : _GEN_1392; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1394 = 6'h32 == _T_284 ? _T_70 : _GEN_1393; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1395 = 6'h33 == _T_284 ? _T_71 : _GEN_1394; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1396 = 6'h34 == _T_284 ? _T_72 : _GEN_1395; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1397 = 6'h35 == _T_284 ? _T_73 : _GEN_1396; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1398 = 6'h36 == _T_284 ? _T_74 : _GEN_1397; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1399 = 6'h37 == _T_284 ? _T_75 : _GEN_1398; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1400 = 6'h38 == _T_284 ? _T_76 : _GEN_1399; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1401 = 6'h39 == _T_284 ? _T_77 : _GEN_1400; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1402 = 6'h3a == _T_284 ? _T_78 : _GEN_1401; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1403 = 6'h3b == _T_284 ? _T_79 : _GEN_1402; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1404 = 6'h3c == _T_284 ? _T_80 : _GEN_1403; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1405 = 6'h3d == _T_284 ? _T_81 : _GEN_1404; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1406 = 6'h3e == _T_284 ? _T_82 : _GEN_1405; // @[execute.scala 79:10:@1927.4]
  assign _GEN_1407 = 6'h3f == _T_284 ? _T_83 : _GEN_1406; // @[execute.scala 79:10:@1927.4]
  assign _T_286 = _T_276 ? _GEN_1343 : _GEN_1407; // @[execute.scala 79:10:@1927.4]
  assign _T_288 = io_amount < 6'h35; // @[execute.scala 79:15:@1928.4]
  assign _T_290 = io_amount - 6'h35; // @[execute.scala 79:37:@1929.4]
  assign _T_291 = $unsigned(_T_290); // @[execute.scala 79:37:@1930.4]
  assign _T_292 = _T_291[5:0]; // @[execute.scala 79:37:@1931.4]
  assign _T_295 = 6'hb + io_amount; // @[execute.scala 79:60:@1932.4]
  assign _T_296 = 6'hb + io_amount; // @[execute.scala 79:60:@1933.4]
  assign _GEN_1409 = 6'h1 == _T_292 ? _T_21 : _T_20; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1410 = 6'h2 == _T_292 ? _T_22 : _GEN_1409; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1411 = 6'h3 == _T_292 ? _T_23 : _GEN_1410; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1412 = 6'h4 == _T_292 ? _T_24 : _GEN_1411; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1413 = 6'h5 == _T_292 ? _T_25 : _GEN_1412; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1414 = 6'h6 == _T_292 ? _T_26 : _GEN_1413; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1415 = 6'h7 == _T_292 ? _T_27 : _GEN_1414; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1416 = 6'h8 == _T_292 ? _T_28 : _GEN_1415; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1417 = 6'h9 == _T_292 ? _T_29 : _GEN_1416; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1418 = 6'ha == _T_292 ? _T_30 : _GEN_1417; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1419 = 6'hb == _T_292 ? _T_31 : _GEN_1418; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1420 = 6'hc == _T_292 ? _T_32 : _GEN_1419; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1421 = 6'hd == _T_292 ? _T_33 : _GEN_1420; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1422 = 6'he == _T_292 ? _T_34 : _GEN_1421; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1423 = 6'hf == _T_292 ? _T_35 : _GEN_1422; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1424 = 6'h10 == _T_292 ? _T_36 : _GEN_1423; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1425 = 6'h11 == _T_292 ? _T_37 : _GEN_1424; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1426 = 6'h12 == _T_292 ? _T_38 : _GEN_1425; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1427 = 6'h13 == _T_292 ? _T_39 : _GEN_1426; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1428 = 6'h14 == _T_292 ? _T_40 : _GEN_1427; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1429 = 6'h15 == _T_292 ? _T_41 : _GEN_1428; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1430 = 6'h16 == _T_292 ? _T_42 : _GEN_1429; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1431 = 6'h17 == _T_292 ? _T_43 : _GEN_1430; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1432 = 6'h18 == _T_292 ? _T_44 : _GEN_1431; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1433 = 6'h19 == _T_292 ? _T_45 : _GEN_1432; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1434 = 6'h1a == _T_292 ? _T_46 : _GEN_1433; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1435 = 6'h1b == _T_292 ? _T_47 : _GEN_1434; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1436 = 6'h1c == _T_292 ? _T_48 : _GEN_1435; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1437 = 6'h1d == _T_292 ? _T_49 : _GEN_1436; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1438 = 6'h1e == _T_292 ? _T_50 : _GEN_1437; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1439 = 6'h1f == _T_292 ? _T_51 : _GEN_1438; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1440 = 6'h20 == _T_292 ? _T_52 : _GEN_1439; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1441 = 6'h21 == _T_292 ? _T_53 : _GEN_1440; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1442 = 6'h22 == _T_292 ? _T_54 : _GEN_1441; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1443 = 6'h23 == _T_292 ? _T_55 : _GEN_1442; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1444 = 6'h24 == _T_292 ? _T_56 : _GEN_1443; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1445 = 6'h25 == _T_292 ? _T_57 : _GEN_1444; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1446 = 6'h26 == _T_292 ? _T_58 : _GEN_1445; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1447 = 6'h27 == _T_292 ? _T_59 : _GEN_1446; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1448 = 6'h28 == _T_292 ? _T_60 : _GEN_1447; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1449 = 6'h29 == _T_292 ? _T_61 : _GEN_1448; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1450 = 6'h2a == _T_292 ? _T_62 : _GEN_1449; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1451 = 6'h2b == _T_292 ? _T_63 : _GEN_1450; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1452 = 6'h2c == _T_292 ? _T_64 : _GEN_1451; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1453 = 6'h2d == _T_292 ? _T_65 : _GEN_1452; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1454 = 6'h2e == _T_292 ? _T_66 : _GEN_1453; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1455 = 6'h2f == _T_292 ? _T_67 : _GEN_1454; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1456 = 6'h30 == _T_292 ? _T_68 : _GEN_1455; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1457 = 6'h31 == _T_292 ? _T_69 : _GEN_1456; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1458 = 6'h32 == _T_292 ? _T_70 : _GEN_1457; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1459 = 6'h33 == _T_292 ? _T_71 : _GEN_1458; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1460 = 6'h34 == _T_292 ? _T_72 : _GEN_1459; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1461 = 6'h35 == _T_292 ? _T_73 : _GEN_1460; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1462 = 6'h36 == _T_292 ? _T_74 : _GEN_1461; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1463 = 6'h37 == _T_292 ? _T_75 : _GEN_1462; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1464 = 6'h38 == _T_292 ? _T_76 : _GEN_1463; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1465 = 6'h39 == _T_292 ? _T_77 : _GEN_1464; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1466 = 6'h3a == _T_292 ? _T_78 : _GEN_1465; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1467 = 6'h3b == _T_292 ? _T_79 : _GEN_1466; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1468 = 6'h3c == _T_292 ? _T_80 : _GEN_1467; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1469 = 6'h3d == _T_292 ? _T_81 : _GEN_1468; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1470 = 6'h3e == _T_292 ? _T_82 : _GEN_1469; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1471 = 6'h3f == _T_292 ? _T_83 : _GEN_1470; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1473 = 6'h1 == _T_296 ? _T_21 : _T_20; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1474 = 6'h2 == _T_296 ? _T_22 : _GEN_1473; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1475 = 6'h3 == _T_296 ? _T_23 : _GEN_1474; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1476 = 6'h4 == _T_296 ? _T_24 : _GEN_1475; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1477 = 6'h5 == _T_296 ? _T_25 : _GEN_1476; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1478 = 6'h6 == _T_296 ? _T_26 : _GEN_1477; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1479 = 6'h7 == _T_296 ? _T_27 : _GEN_1478; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1480 = 6'h8 == _T_296 ? _T_28 : _GEN_1479; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1481 = 6'h9 == _T_296 ? _T_29 : _GEN_1480; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1482 = 6'ha == _T_296 ? _T_30 : _GEN_1481; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1483 = 6'hb == _T_296 ? _T_31 : _GEN_1482; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1484 = 6'hc == _T_296 ? _T_32 : _GEN_1483; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1485 = 6'hd == _T_296 ? _T_33 : _GEN_1484; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1486 = 6'he == _T_296 ? _T_34 : _GEN_1485; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1487 = 6'hf == _T_296 ? _T_35 : _GEN_1486; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1488 = 6'h10 == _T_296 ? _T_36 : _GEN_1487; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1489 = 6'h11 == _T_296 ? _T_37 : _GEN_1488; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1490 = 6'h12 == _T_296 ? _T_38 : _GEN_1489; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1491 = 6'h13 == _T_296 ? _T_39 : _GEN_1490; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1492 = 6'h14 == _T_296 ? _T_40 : _GEN_1491; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1493 = 6'h15 == _T_296 ? _T_41 : _GEN_1492; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1494 = 6'h16 == _T_296 ? _T_42 : _GEN_1493; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1495 = 6'h17 == _T_296 ? _T_43 : _GEN_1494; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1496 = 6'h18 == _T_296 ? _T_44 : _GEN_1495; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1497 = 6'h19 == _T_296 ? _T_45 : _GEN_1496; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1498 = 6'h1a == _T_296 ? _T_46 : _GEN_1497; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1499 = 6'h1b == _T_296 ? _T_47 : _GEN_1498; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1500 = 6'h1c == _T_296 ? _T_48 : _GEN_1499; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1501 = 6'h1d == _T_296 ? _T_49 : _GEN_1500; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1502 = 6'h1e == _T_296 ? _T_50 : _GEN_1501; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1503 = 6'h1f == _T_296 ? _T_51 : _GEN_1502; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1504 = 6'h20 == _T_296 ? _T_52 : _GEN_1503; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1505 = 6'h21 == _T_296 ? _T_53 : _GEN_1504; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1506 = 6'h22 == _T_296 ? _T_54 : _GEN_1505; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1507 = 6'h23 == _T_296 ? _T_55 : _GEN_1506; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1508 = 6'h24 == _T_296 ? _T_56 : _GEN_1507; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1509 = 6'h25 == _T_296 ? _T_57 : _GEN_1508; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1510 = 6'h26 == _T_296 ? _T_58 : _GEN_1509; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1511 = 6'h27 == _T_296 ? _T_59 : _GEN_1510; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1512 = 6'h28 == _T_296 ? _T_60 : _GEN_1511; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1513 = 6'h29 == _T_296 ? _T_61 : _GEN_1512; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1514 = 6'h2a == _T_296 ? _T_62 : _GEN_1513; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1515 = 6'h2b == _T_296 ? _T_63 : _GEN_1514; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1516 = 6'h2c == _T_296 ? _T_64 : _GEN_1515; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1517 = 6'h2d == _T_296 ? _T_65 : _GEN_1516; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1518 = 6'h2e == _T_296 ? _T_66 : _GEN_1517; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1519 = 6'h2f == _T_296 ? _T_67 : _GEN_1518; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1520 = 6'h30 == _T_296 ? _T_68 : _GEN_1519; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1521 = 6'h31 == _T_296 ? _T_69 : _GEN_1520; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1522 = 6'h32 == _T_296 ? _T_70 : _GEN_1521; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1523 = 6'h33 == _T_296 ? _T_71 : _GEN_1522; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1524 = 6'h34 == _T_296 ? _T_72 : _GEN_1523; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1525 = 6'h35 == _T_296 ? _T_73 : _GEN_1524; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1526 = 6'h36 == _T_296 ? _T_74 : _GEN_1525; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1527 = 6'h37 == _T_296 ? _T_75 : _GEN_1526; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1528 = 6'h38 == _T_296 ? _T_76 : _GEN_1527; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1529 = 6'h39 == _T_296 ? _T_77 : _GEN_1528; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1530 = 6'h3a == _T_296 ? _T_78 : _GEN_1529; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1531 = 6'h3b == _T_296 ? _T_79 : _GEN_1530; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1532 = 6'h3c == _T_296 ? _T_80 : _GEN_1531; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1533 = 6'h3d == _T_296 ? _T_81 : _GEN_1532; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1534 = 6'h3e == _T_296 ? _T_82 : _GEN_1533; // @[execute.scala 79:10:@1934.4]
  assign _GEN_1535 = 6'h3f == _T_296 ? _T_83 : _GEN_1534; // @[execute.scala 79:10:@1934.4]
  assign _T_298 = _T_288 ? _GEN_1471 : _GEN_1535; // @[execute.scala 79:10:@1934.4]
  assign _T_300 = io_amount < 6'h34; // @[execute.scala 79:15:@1935.4]
  assign _T_302 = io_amount - 6'h34; // @[execute.scala 79:37:@1936.4]
  assign _T_303 = $unsigned(_T_302); // @[execute.scala 79:37:@1937.4]
  assign _T_304 = _T_303[5:0]; // @[execute.scala 79:37:@1938.4]
  assign _T_307 = 6'hc + io_amount; // @[execute.scala 79:60:@1939.4]
  assign _T_308 = 6'hc + io_amount; // @[execute.scala 79:60:@1940.4]
  assign _GEN_1537 = 6'h1 == _T_304 ? _T_21 : _T_20; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1538 = 6'h2 == _T_304 ? _T_22 : _GEN_1537; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1539 = 6'h3 == _T_304 ? _T_23 : _GEN_1538; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1540 = 6'h4 == _T_304 ? _T_24 : _GEN_1539; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1541 = 6'h5 == _T_304 ? _T_25 : _GEN_1540; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1542 = 6'h6 == _T_304 ? _T_26 : _GEN_1541; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1543 = 6'h7 == _T_304 ? _T_27 : _GEN_1542; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1544 = 6'h8 == _T_304 ? _T_28 : _GEN_1543; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1545 = 6'h9 == _T_304 ? _T_29 : _GEN_1544; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1546 = 6'ha == _T_304 ? _T_30 : _GEN_1545; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1547 = 6'hb == _T_304 ? _T_31 : _GEN_1546; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1548 = 6'hc == _T_304 ? _T_32 : _GEN_1547; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1549 = 6'hd == _T_304 ? _T_33 : _GEN_1548; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1550 = 6'he == _T_304 ? _T_34 : _GEN_1549; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1551 = 6'hf == _T_304 ? _T_35 : _GEN_1550; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1552 = 6'h10 == _T_304 ? _T_36 : _GEN_1551; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1553 = 6'h11 == _T_304 ? _T_37 : _GEN_1552; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1554 = 6'h12 == _T_304 ? _T_38 : _GEN_1553; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1555 = 6'h13 == _T_304 ? _T_39 : _GEN_1554; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1556 = 6'h14 == _T_304 ? _T_40 : _GEN_1555; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1557 = 6'h15 == _T_304 ? _T_41 : _GEN_1556; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1558 = 6'h16 == _T_304 ? _T_42 : _GEN_1557; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1559 = 6'h17 == _T_304 ? _T_43 : _GEN_1558; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1560 = 6'h18 == _T_304 ? _T_44 : _GEN_1559; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1561 = 6'h19 == _T_304 ? _T_45 : _GEN_1560; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1562 = 6'h1a == _T_304 ? _T_46 : _GEN_1561; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1563 = 6'h1b == _T_304 ? _T_47 : _GEN_1562; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1564 = 6'h1c == _T_304 ? _T_48 : _GEN_1563; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1565 = 6'h1d == _T_304 ? _T_49 : _GEN_1564; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1566 = 6'h1e == _T_304 ? _T_50 : _GEN_1565; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1567 = 6'h1f == _T_304 ? _T_51 : _GEN_1566; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1568 = 6'h20 == _T_304 ? _T_52 : _GEN_1567; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1569 = 6'h21 == _T_304 ? _T_53 : _GEN_1568; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1570 = 6'h22 == _T_304 ? _T_54 : _GEN_1569; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1571 = 6'h23 == _T_304 ? _T_55 : _GEN_1570; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1572 = 6'h24 == _T_304 ? _T_56 : _GEN_1571; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1573 = 6'h25 == _T_304 ? _T_57 : _GEN_1572; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1574 = 6'h26 == _T_304 ? _T_58 : _GEN_1573; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1575 = 6'h27 == _T_304 ? _T_59 : _GEN_1574; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1576 = 6'h28 == _T_304 ? _T_60 : _GEN_1575; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1577 = 6'h29 == _T_304 ? _T_61 : _GEN_1576; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1578 = 6'h2a == _T_304 ? _T_62 : _GEN_1577; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1579 = 6'h2b == _T_304 ? _T_63 : _GEN_1578; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1580 = 6'h2c == _T_304 ? _T_64 : _GEN_1579; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1581 = 6'h2d == _T_304 ? _T_65 : _GEN_1580; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1582 = 6'h2e == _T_304 ? _T_66 : _GEN_1581; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1583 = 6'h2f == _T_304 ? _T_67 : _GEN_1582; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1584 = 6'h30 == _T_304 ? _T_68 : _GEN_1583; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1585 = 6'h31 == _T_304 ? _T_69 : _GEN_1584; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1586 = 6'h32 == _T_304 ? _T_70 : _GEN_1585; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1587 = 6'h33 == _T_304 ? _T_71 : _GEN_1586; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1588 = 6'h34 == _T_304 ? _T_72 : _GEN_1587; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1589 = 6'h35 == _T_304 ? _T_73 : _GEN_1588; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1590 = 6'h36 == _T_304 ? _T_74 : _GEN_1589; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1591 = 6'h37 == _T_304 ? _T_75 : _GEN_1590; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1592 = 6'h38 == _T_304 ? _T_76 : _GEN_1591; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1593 = 6'h39 == _T_304 ? _T_77 : _GEN_1592; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1594 = 6'h3a == _T_304 ? _T_78 : _GEN_1593; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1595 = 6'h3b == _T_304 ? _T_79 : _GEN_1594; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1596 = 6'h3c == _T_304 ? _T_80 : _GEN_1595; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1597 = 6'h3d == _T_304 ? _T_81 : _GEN_1596; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1598 = 6'h3e == _T_304 ? _T_82 : _GEN_1597; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1599 = 6'h3f == _T_304 ? _T_83 : _GEN_1598; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1601 = 6'h1 == _T_308 ? _T_21 : _T_20; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1602 = 6'h2 == _T_308 ? _T_22 : _GEN_1601; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1603 = 6'h3 == _T_308 ? _T_23 : _GEN_1602; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1604 = 6'h4 == _T_308 ? _T_24 : _GEN_1603; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1605 = 6'h5 == _T_308 ? _T_25 : _GEN_1604; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1606 = 6'h6 == _T_308 ? _T_26 : _GEN_1605; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1607 = 6'h7 == _T_308 ? _T_27 : _GEN_1606; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1608 = 6'h8 == _T_308 ? _T_28 : _GEN_1607; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1609 = 6'h9 == _T_308 ? _T_29 : _GEN_1608; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1610 = 6'ha == _T_308 ? _T_30 : _GEN_1609; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1611 = 6'hb == _T_308 ? _T_31 : _GEN_1610; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1612 = 6'hc == _T_308 ? _T_32 : _GEN_1611; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1613 = 6'hd == _T_308 ? _T_33 : _GEN_1612; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1614 = 6'he == _T_308 ? _T_34 : _GEN_1613; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1615 = 6'hf == _T_308 ? _T_35 : _GEN_1614; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1616 = 6'h10 == _T_308 ? _T_36 : _GEN_1615; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1617 = 6'h11 == _T_308 ? _T_37 : _GEN_1616; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1618 = 6'h12 == _T_308 ? _T_38 : _GEN_1617; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1619 = 6'h13 == _T_308 ? _T_39 : _GEN_1618; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1620 = 6'h14 == _T_308 ? _T_40 : _GEN_1619; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1621 = 6'h15 == _T_308 ? _T_41 : _GEN_1620; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1622 = 6'h16 == _T_308 ? _T_42 : _GEN_1621; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1623 = 6'h17 == _T_308 ? _T_43 : _GEN_1622; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1624 = 6'h18 == _T_308 ? _T_44 : _GEN_1623; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1625 = 6'h19 == _T_308 ? _T_45 : _GEN_1624; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1626 = 6'h1a == _T_308 ? _T_46 : _GEN_1625; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1627 = 6'h1b == _T_308 ? _T_47 : _GEN_1626; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1628 = 6'h1c == _T_308 ? _T_48 : _GEN_1627; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1629 = 6'h1d == _T_308 ? _T_49 : _GEN_1628; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1630 = 6'h1e == _T_308 ? _T_50 : _GEN_1629; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1631 = 6'h1f == _T_308 ? _T_51 : _GEN_1630; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1632 = 6'h20 == _T_308 ? _T_52 : _GEN_1631; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1633 = 6'h21 == _T_308 ? _T_53 : _GEN_1632; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1634 = 6'h22 == _T_308 ? _T_54 : _GEN_1633; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1635 = 6'h23 == _T_308 ? _T_55 : _GEN_1634; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1636 = 6'h24 == _T_308 ? _T_56 : _GEN_1635; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1637 = 6'h25 == _T_308 ? _T_57 : _GEN_1636; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1638 = 6'h26 == _T_308 ? _T_58 : _GEN_1637; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1639 = 6'h27 == _T_308 ? _T_59 : _GEN_1638; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1640 = 6'h28 == _T_308 ? _T_60 : _GEN_1639; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1641 = 6'h29 == _T_308 ? _T_61 : _GEN_1640; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1642 = 6'h2a == _T_308 ? _T_62 : _GEN_1641; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1643 = 6'h2b == _T_308 ? _T_63 : _GEN_1642; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1644 = 6'h2c == _T_308 ? _T_64 : _GEN_1643; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1645 = 6'h2d == _T_308 ? _T_65 : _GEN_1644; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1646 = 6'h2e == _T_308 ? _T_66 : _GEN_1645; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1647 = 6'h2f == _T_308 ? _T_67 : _GEN_1646; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1648 = 6'h30 == _T_308 ? _T_68 : _GEN_1647; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1649 = 6'h31 == _T_308 ? _T_69 : _GEN_1648; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1650 = 6'h32 == _T_308 ? _T_70 : _GEN_1649; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1651 = 6'h33 == _T_308 ? _T_71 : _GEN_1650; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1652 = 6'h34 == _T_308 ? _T_72 : _GEN_1651; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1653 = 6'h35 == _T_308 ? _T_73 : _GEN_1652; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1654 = 6'h36 == _T_308 ? _T_74 : _GEN_1653; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1655 = 6'h37 == _T_308 ? _T_75 : _GEN_1654; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1656 = 6'h38 == _T_308 ? _T_76 : _GEN_1655; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1657 = 6'h39 == _T_308 ? _T_77 : _GEN_1656; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1658 = 6'h3a == _T_308 ? _T_78 : _GEN_1657; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1659 = 6'h3b == _T_308 ? _T_79 : _GEN_1658; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1660 = 6'h3c == _T_308 ? _T_80 : _GEN_1659; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1661 = 6'h3d == _T_308 ? _T_81 : _GEN_1660; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1662 = 6'h3e == _T_308 ? _T_82 : _GEN_1661; // @[execute.scala 79:10:@1941.4]
  assign _GEN_1663 = 6'h3f == _T_308 ? _T_83 : _GEN_1662; // @[execute.scala 79:10:@1941.4]
  assign _T_310 = _T_300 ? _GEN_1599 : _GEN_1663; // @[execute.scala 79:10:@1941.4]
  assign _T_312 = io_amount < 6'h33; // @[execute.scala 79:15:@1942.4]
  assign _T_314 = io_amount - 6'h33; // @[execute.scala 79:37:@1943.4]
  assign _T_315 = $unsigned(_T_314); // @[execute.scala 79:37:@1944.4]
  assign _T_316 = _T_315[5:0]; // @[execute.scala 79:37:@1945.4]
  assign _T_319 = 6'hd + io_amount; // @[execute.scala 79:60:@1946.4]
  assign _T_320 = 6'hd + io_amount; // @[execute.scala 79:60:@1947.4]
  assign _GEN_1665 = 6'h1 == _T_316 ? _T_21 : _T_20; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1666 = 6'h2 == _T_316 ? _T_22 : _GEN_1665; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1667 = 6'h3 == _T_316 ? _T_23 : _GEN_1666; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1668 = 6'h4 == _T_316 ? _T_24 : _GEN_1667; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1669 = 6'h5 == _T_316 ? _T_25 : _GEN_1668; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1670 = 6'h6 == _T_316 ? _T_26 : _GEN_1669; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1671 = 6'h7 == _T_316 ? _T_27 : _GEN_1670; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1672 = 6'h8 == _T_316 ? _T_28 : _GEN_1671; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1673 = 6'h9 == _T_316 ? _T_29 : _GEN_1672; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1674 = 6'ha == _T_316 ? _T_30 : _GEN_1673; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1675 = 6'hb == _T_316 ? _T_31 : _GEN_1674; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1676 = 6'hc == _T_316 ? _T_32 : _GEN_1675; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1677 = 6'hd == _T_316 ? _T_33 : _GEN_1676; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1678 = 6'he == _T_316 ? _T_34 : _GEN_1677; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1679 = 6'hf == _T_316 ? _T_35 : _GEN_1678; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1680 = 6'h10 == _T_316 ? _T_36 : _GEN_1679; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1681 = 6'h11 == _T_316 ? _T_37 : _GEN_1680; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1682 = 6'h12 == _T_316 ? _T_38 : _GEN_1681; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1683 = 6'h13 == _T_316 ? _T_39 : _GEN_1682; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1684 = 6'h14 == _T_316 ? _T_40 : _GEN_1683; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1685 = 6'h15 == _T_316 ? _T_41 : _GEN_1684; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1686 = 6'h16 == _T_316 ? _T_42 : _GEN_1685; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1687 = 6'h17 == _T_316 ? _T_43 : _GEN_1686; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1688 = 6'h18 == _T_316 ? _T_44 : _GEN_1687; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1689 = 6'h19 == _T_316 ? _T_45 : _GEN_1688; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1690 = 6'h1a == _T_316 ? _T_46 : _GEN_1689; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1691 = 6'h1b == _T_316 ? _T_47 : _GEN_1690; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1692 = 6'h1c == _T_316 ? _T_48 : _GEN_1691; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1693 = 6'h1d == _T_316 ? _T_49 : _GEN_1692; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1694 = 6'h1e == _T_316 ? _T_50 : _GEN_1693; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1695 = 6'h1f == _T_316 ? _T_51 : _GEN_1694; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1696 = 6'h20 == _T_316 ? _T_52 : _GEN_1695; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1697 = 6'h21 == _T_316 ? _T_53 : _GEN_1696; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1698 = 6'h22 == _T_316 ? _T_54 : _GEN_1697; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1699 = 6'h23 == _T_316 ? _T_55 : _GEN_1698; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1700 = 6'h24 == _T_316 ? _T_56 : _GEN_1699; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1701 = 6'h25 == _T_316 ? _T_57 : _GEN_1700; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1702 = 6'h26 == _T_316 ? _T_58 : _GEN_1701; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1703 = 6'h27 == _T_316 ? _T_59 : _GEN_1702; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1704 = 6'h28 == _T_316 ? _T_60 : _GEN_1703; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1705 = 6'h29 == _T_316 ? _T_61 : _GEN_1704; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1706 = 6'h2a == _T_316 ? _T_62 : _GEN_1705; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1707 = 6'h2b == _T_316 ? _T_63 : _GEN_1706; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1708 = 6'h2c == _T_316 ? _T_64 : _GEN_1707; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1709 = 6'h2d == _T_316 ? _T_65 : _GEN_1708; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1710 = 6'h2e == _T_316 ? _T_66 : _GEN_1709; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1711 = 6'h2f == _T_316 ? _T_67 : _GEN_1710; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1712 = 6'h30 == _T_316 ? _T_68 : _GEN_1711; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1713 = 6'h31 == _T_316 ? _T_69 : _GEN_1712; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1714 = 6'h32 == _T_316 ? _T_70 : _GEN_1713; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1715 = 6'h33 == _T_316 ? _T_71 : _GEN_1714; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1716 = 6'h34 == _T_316 ? _T_72 : _GEN_1715; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1717 = 6'h35 == _T_316 ? _T_73 : _GEN_1716; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1718 = 6'h36 == _T_316 ? _T_74 : _GEN_1717; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1719 = 6'h37 == _T_316 ? _T_75 : _GEN_1718; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1720 = 6'h38 == _T_316 ? _T_76 : _GEN_1719; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1721 = 6'h39 == _T_316 ? _T_77 : _GEN_1720; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1722 = 6'h3a == _T_316 ? _T_78 : _GEN_1721; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1723 = 6'h3b == _T_316 ? _T_79 : _GEN_1722; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1724 = 6'h3c == _T_316 ? _T_80 : _GEN_1723; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1725 = 6'h3d == _T_316 ? _T_81 : _GEN_1724; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1726 = 6'h3e == _T_316 ? _T_82 : _GEN_1725; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1727 = 6'h3f == _T_316 ? _T_83 : _GEN_1726; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1729 = 6'h1 == _T_320 ? _T_21 : _T_20; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1730 = 6'h2 == _T_320 ? _T_22 : _GEN_1729; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1731 = 6'h3 == _T_320 ? _T_23 : _GEN_1730; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1732 = 6'h4 == _T_320 ? _T_24 : _GEN_1731; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1733 = 6'h5 == _T_320 ? _T_25 : _GEN_1732; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1734 = 6'h6 == _T_320 ? _T_26 : _GEN_1733; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1735 = 6'h7 == _T_320 ? _T_27 : _GEN_1734; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1736 = 6'h8 == _T_320 ? _T_28 : _GEN_1735; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1737 = 6'h9 == _T_320 ? _T_29 : _GEN_1736; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1738 = 6'ha == _T_320 ? _T_30 : _GEN_1737; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1739 = 6'hb == _T_320 ? _T_31 : _GEN_1738; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1740 = 6'hc == _T_320 ? _T_32 : _GEN_1739; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1741 = 6'hd == _T_320 ? _T_33 : _GEN_1740; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1742 = 6'he == _T_320 ? _T_34 : _GEN_1741; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1743 = 6'hf == _T_320 ? _T_35 : _GEN_1742; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1744 = 6'h10 == _T_320 ? _T_36 : _GEN_1743; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1745 = 6'h11 == _T_320 ? _T_37 : _GEN_1744; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1746 = 6'h12 == _T_320 ? _T_38 : _GEN_1745; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1747 = 6'h13 == _T_320 ? _T_39 : _GEN_1746; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1748 = 6'h14 == _T_320 ? _T_40 : _GEN_1747; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1749 = 6'h15 == _T_320 ? _T_41 : _GEN_1748; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1750 = 6'h16 == _T_320 ? _T_42 : _GEN_1749; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1751 = 6'h17 == _T_320 ? _T_43 : _GEN_1750; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1752 = 6'h18 == _T_320 ? _T_44 : _GEN_1751; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1753 = 6'h19 == _T_320 ? _T_45 : _GEN_1752; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1754 = 6'h1a == _T_320 ? _T_46 : _GEN_1753; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1755 = 6'h1b == _T_320 ? _T_47 : _GEN_1754; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1756 = 6'h1c == _T_320 ? _T_48 : _GEN_1755; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1757 = 6'h1d == _T_320 ? _T_49 : _GEN_1756; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1758 = 6'h1e == _T_320 ? _T_50 : _GEN_1757; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1759 = 6'h1f == _T_320 ? _T_51 : _GEN_1758; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1760 = 6'h20 == _T_320 ? _T_52 : _GEN_1759; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1761 = 6'h21 == _T_320 ? _T_53 : _GEN_1760; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1762 = 6'h22 == _T_320 ? _T_54 : _GEN_1761; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1763 = 6'h23 == _T_320 ? _T_55 : _GEN_1762; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1764 = 6'h24 == _T_320 ? _T_56 : _GEN_1763; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1765 = 6'h25 == _T_320 ? _T_57 : _GEN_1764; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1766 = 6'h26 == _T_320 ? _T_58 : _GEN_1765; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1767 = 6'h27 == _T_320 ? _T_59 : _GEN_1766; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1768 = 6'h28 == _T_320 ? _T_60 : _GEN_1767; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1769 = 6'h29 == _T_320 ? _T_61 : _GEN_1768; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1770 = 6'h2a == _T_320 ? _T_62 : _GEN_1769; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1771 = 6'h2b == _T_320 ? _T_63 : _GEN_1770; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1772 = 6'h2c == _T_320 ? _T_64 : _GEN_1771; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1773 = 6'h2d == _T_320 ? _T_65 : _GEN_1772; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1774 = 6'h2e == _T_320 ? _T_66 : _GEN_1773; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1775 = 6'h2f == _T_320 ? _T_67 : _GEN_1774; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1776 = 6'h30 == _T_320 ? _T_68 : _GEN_1775; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1777 = 6'h31 == _T_320 ? _T_69 : _GEN_1776; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1778 = 6'h32 == _T_320 ? _T_70 : _GEN_1777; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1779 = 6'h33 == _T_320 ? _T_71 : _GEN_1778; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1780 = 6'h34 == _T_320 ? _T_72 : _GEN_1779; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1781 = 6'h35 == _T_320 ? _T_73 : _GEN_1780; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1782 = 6'h36 == _T_320 ? _T_74 : _GEN_1781; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1783 = 6'h37 == _T_320 ? _T_75 : _GEN_1782; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1784 = 6'h38 == _T_320 ? _T_76 : _GEN_1783; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1785 = 6'h39 == _T_320 ? _T_77 : _GEN_1784; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1786 = 6'h3a == _T_320 ? _T_78 : _GEN_1785; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1787 = 6'h3b == _T_320 ? _T_79 : _GEN_1786; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1788 = 6'h3c == _T_320 ? _T_80 : _GEN_1787; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1789 = 6'h3d == _T_320 ? _T_81 : _GEN_1788; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1790 = 6'h3e == _T_320 ? _T_82 : _GEN_1789; // @[execute.scala 79:10:@1948.4]
  assign _GEN_1791 = 6'h3f == _T_320 ? _T_83 : _GEN_1790; // @[execute.scala 79:10:@1948.4]
  assign _T_322 = _T_312 ? _GEN_1727 : _GEN_1791; // @[execute.scala 79:10:@1948.4]
  assign _T_324 = io_amount < 6'h32; // @[execute.scala 79:15:@1949.4]
  assign _T_326 = io_amount - 6'h32; // @[execute.scala 79:37:@1950.4]
  assign _T_327 = $unsigned(_T_326); // @[execute.scala 79:37:@1951.4]
  assign _T_328 = _T_327[5:0]; // @[execute.scala 79:37:@1952.4]
  assign _T_331 = 6'he + io_amount; // @[execute.scala 79:60:@1953.4]
  assign _T_332 = 6'he + io_amount; // @[execute.scala 79:60:@1954.4]
  assign _GEN_1793 = 6'h1 == _T_328 ? _T_21 : _T_20; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1794 = 6'h2 == _T_328 ? _T_22 : _GEN_1793; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1795 = 6'h3 == _T_328 ? _T_23 : _GEN_1794; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1796 = 6'h4 == _T_328 ? _T_24 : _GEN_1795; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1797 = 6'h5 == _T_328 ? _T_25 : _GEN_1796; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1798 = 6'h6 == _T_328 ? _T_26 : _GEN_1797; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1799 = 6'h7 == _T_328 ? _T_27 : _GEN_1798; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1800 = 6'h8 == _T_328 ? _T_28 : _GEN_1799; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1801 = 6'h9 == _T_328 ? _T_29 : _GEN_1800; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1802 = 6'ha == _T_328 ? _T_30 : _GEN_1801; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1803 = 6'hb == _T_328 ? _T_31 : _GEN_1802; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1804 = 6'hc == _T_328 ? _T_32 : _GEN_1803; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1805 = 6'hd == _T_328 ? _T_33 : _GEN_1804; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1806 = 6'he == _T_328 ? _T_34 : _GEN_1805; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1807 = 6'hf == _T_328 ? _T_35 : _GEN_1806; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1808 = 6'h10 == _T_328 ? _T_36 : _GEN_1807; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1809 = 6'h11 == _T_328 ? _T_37 : _GEN_1808; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1810 = 6'h12 == _T_328 ? _T_38 : _GEN_1809; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1811 = 6'h13 == _T_328 ? _T_39 : _GEN_1810; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1812 = 6'h14 == _T_328 ? _T_40 : _GEN_1811; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1813 = 6'h15 == _T_328 ? _T_41 : _GEN_1812; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1814 = 6'h16 == _T_328 ? _T_42 : _GEN_1813; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1815 = 6'h17 == _T_328 ? _T_43 : _GEN_1814; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1816 = 6'h18 == _T_328 ? _T_44 : _GEN_1815; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1817 = 6'h19 == _T_328 ? _T_45 : _GEN_1816; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1818 = 6'h1a == _T_328 ? _T_46 : _GEN_1817; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1819 = 6'h1b == _T_328 ? _T_47 : _GEN_1818; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1820 = 6'h1c == _T_328 ? _T_48 : _GEN_1819; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1821 = 6'h1d == _T_328 ? _T_49 : _GEN_1820; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1822 = 6'h1e == _T_328 ? _T_50 : _GEN_1821; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1823 = 6'h1f == _T_328 ? _T_51 : _GEN_1822; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1824 = 6'h20 == _T_328 ? _T_52 : _GEN_1823; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1825 = 6'h21 == _T_328 ? _T_53 : _GEN_1824; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1826 = 6'h22 == _T_328 ? _T_54 : _GEN_1825; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1827 = 6'h23 == _T_328 ? _T_55 : _GEN_1826; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1828 = 6'h24 == _T_328 ? _T_56 : _GEN_1827; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1829 = 6'h25 == _T_328 ? _T_57 : _GEN_1828; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1830 = 6'h26 == _T_328 ? _T_58 : _GEN_1829; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1831 = 6'h27 == _T_328 ? _T_59 : _GEN_1830; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1832 = 6'h28 == _T_328 ? _T_60 : _GEN_1831; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1833 = 6'h29 == _T_328 ? _T_61 : _GEN_1832; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1834 = 6'h2a == _T_328 ? _T_62 : _GEN_1833; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1835 = 6'h2b == _T_328 ? _T_63 : _GEN_1834; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1836 = 6'h2c == _T_328 ? _T_64 : _GEN_1835; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1837 = 6'h2d == _T_328 ? _T_65 : _GEN_1836; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1838 = 6'h2e == _T_328 ? _T_66 : _GEN_1837; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1839 = 6'h2f == _T_328 ? _T_67 : _GEN_1838; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1840 = 6'h30 == _T_328 ? _T_68 : _GEN_1839; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1841 = 6'h31 == _T_328 ? _T_69 : _GEN_1840; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1842 = 6'h32 == _T_328 ? _T_70 : _GEN_1841; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1843 = 6'h33 == _T_328 ? _T_71 : _GEN_1842; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1844 = 6'h34 == _T_328 ? _T_72 : _GEN_1843; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1845 = 6'h35 == _T_328 ? _T_73 : _GEN_1844; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1846 = 6'h36 == _T_328 ? _T_74 : _GEN_1845; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1847 = 6'h37 == _T_328 ? _T_75 : _GEN_1846; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1848 = 6'h38 == _T_328 ? _T_76 : _GEN_1847; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1849 = 6'h39 == _T_328 ? _T_77 : _GEN_1848; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1850 = 6'h3a == _T_328 ? _T_78 : _GEN_1849; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1851 = 6'h3b == _T_328 ? _T_79 : _GEN_1850; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1852 = 6'h3c == _T_328 ? _T_80 : _GEN_1851; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1853 = 6'h3d == _T_328 ? _T_81 : _GEN_1852; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1854 = 6'h3e == _T_328 ? _T_82 : _GEN_1853; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1855 = 6'h3f == _T_328 ? _T_83 : _GEN_1854; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1857 = 6'h1 == _T_332 ? _T_21 : _T_20; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1858 = 6'h2 == _T_332 ? _T_22 : _GEN_1857; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1859 = 6'h3 == _T_332 ? _T_23 : _GEN_1858; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1860 = 6'h4 == _T_332 ? _T_24 : _GEN_1859; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1861 = 6'h5 == _T_332 ? _T_25 : _GEN_1860; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1862 = 6'h6 == _T_332 ? _T_26 : _GEN_1861; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1863 = 6'h7 == _T_332 ? _T_27 : _GEN_1862; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1864 = 6'h8 == _T_332 ? _T_28 : _GEN_1863; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1865 = 6'h9 == _T_332 ? _T_29 : _GEN_1864; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1866 = 6'ha == _T_332 ? _T_30 : _GEN_1865; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1867 = 6'hb == _T_332 ? _T_31 : _GEN_1866; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1868 = 6'hc == _T_332 ? _T_32 : _GEN_1867; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1869 = 6'hd == _T_332 ? _T_33 : _GEN_1868; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1870 = 6'he == _T_332 ? _T_34 : _GEN_1869; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1871 = 6'hf == _T_332 ? _T_35 : _GEN_1870; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1872 = 6'h10 == _T_332 ? _T_36 : _GEN_1871; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1873 = 6'h11 == _T_332 ? _T_37 : _GEN_1872; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1874 = 6'h12 == _T_332 ? _T_38 : _GEN_1873; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1875 = 6'h13 == _T_332 ? _T_39 : _GEN_1874; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1876 = 6'h14 == _T_332 ? _T_40 : _GEN_1875; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1877 = 6'h15 == _T_332 ? _T_41 : _GEN_1876; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1878 = 6'h16 == _T_332 ? _T_42 : _GEN_1877; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1879 = 6'h17 == _T_332 ? _T_43 : _GEN_1878; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1880 = 6'h18 == _T_332 ? _T_44 : _GEN_1879; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1881 = 6'h19 == _T_332 ? _T_45 : _GEN_1880; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1882 = 6'h1a == _T_332 ? _T_46 : _GEN_1881; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1883 = 6'h1b == _T_332 ? _T_47 : _GEN_1882; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1884 = 6'h1c == _T_332 ? _T_48 : _GEN_1883; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1885 = 6'h1d == _T_332 ? _T_49 : _GEN_1884; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1886 = 6'h1e == _T_332 ? _T_50 : _GEN_1885; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1887 = 6'h1f == _T_332 ? _T_51 : _GEN_1886; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1888 = 6'h20 == _T_332 ? _T_52 : _GEN_1887; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1889 = 6'h21 == _T_332 ? _T_53 : _GEN_1888; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1890 = 6'h22 == _T_332 ? _T_54 : _GEN_1889; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1891 = 6'h23 == _T_332 ? _T_55 : _GEN_1890; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1892 = 6'h24 == _T_332 ? _T_56 : _GEN_1891; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1893 = 6'h25 == _T_332 ? _T_57 : _GEN_1892; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1894 = 6'h26 == _T_332 ? _T_58 : _GEN_1893; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1895 = 6'h27 == _T_332 ? _T_59 : _GEN_1894; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1896 = 6'h28 == _T_332 ? _T_60 : _GEN_1895; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1897 = 6'h29 == _T_332 ? _T_61 : _GEN_1896; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1898 = 6'h2a == _T_332 ? _T_62 : _GEN_1897; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1899 = 6'h2b == _T_332 ? _T_63 : _GEN_1898; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1900 = 6'h2c == _T_332 ? _T_64 : _GEN_1899; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1901 = 6'h2d == _T_332 ? _T_65 : _GEN_1900; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1902 = 6'h2e == _T_332 ? _T_66 : _GEN_1901; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1903 = 6'h2f == _T_332 ? _T_67 : _GEN_1902; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1904 = 6'h30 == _T_332 ? _T_68 : _GEN_1903; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1905 = 6'h31 == _T_332 ? _T_69 : _GEN_1904; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1906 = 6'h32 == _T_332 ? _T_70 : _GEN_1905; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1907 = 6'h33 == _T_332 ? _T_71 : _GEN_1906; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1908 = 6'h34 == _T_332 ? _T_72 : _GEN_1907; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1909 = 6'h35 == _T_332 ? _T_73 : _GEN_1908; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1910 = 6'h36 == _T_332 ? _T_74 : _GEN_1909; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1911 = 6'h37 == _T_332 ? _T_75 : _GEN_1910; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1912 = 6'h38 == _T_332 ? _T_76 : _GEN_1911; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1913 = 6'h39 == _T_332 ? _T_77 : _GEN_1912; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1914 = 6'h3a == _T_332 ? _T_78 : _GEN_1913; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1915 = 6'h3b == _T_332 ? _T_79 : _GEN_1914; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1916 = 6'h3c == _T_332 ? _T_80 : _GEN_1915; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1917 = 6'h3d == _T_332 ? _T_81 : _GEN_1916; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1918 = 6'h3e == _T_332 ? _T_82 : _GEN_1917; // @[execute.scala 79:10:@1955.4]
  assign _GEN_1919 = 6'h3f == _T_332 ? _T_83 : _GEN_1918; // @[execute.scala 79:10:@1955.4]
  assign _T_334 = _T_324 ? _GEN_1855 : _GEN_1919; // @[execute.scala 79:10:@1955.4]
  assign _T_336 = io_amount < 6'h31; // @[execute.scala 79:15:@1956.4]
  assign _T_338 = io_amount - 6'h31; // @[execute.scala 79:37:@1957.4]
  assign _T_339 = $unsigned(_T_338); // @[execute.scala 79:37:@1958.4]
  assign _T_340 = _T_339[5:0]; // @[execute.scala 79:37:@1959.4]
  assign _T_343 = 6'hf + io_amount; // @[execute.scala 79:60:@1960.4]
  assign _T_344 = 6'hf + io_amount; // @[execute.scala 79:60:@1961.4]
  assign _GEN_1921 = 6'h1 == _T_340 ? _T_21 : _T_20; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1922 = 6'h2 == _T_340 ? _T_22 : _GEN_1921; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1923 = 6'h3 == _T_340 ? _T_23 : _GEN_1922; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1924 = 6'h4 == _T_340 ? _T_24 : _GEN_1923; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1925 = 6'h5 == _T_340 ? _T_25 : _GEN_1924; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1926 = 6'h6 == _T_340 ? _T_26 : _GEN_1925; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1927 = 6'h7 == _T_340 ? _T_27 : _GEN_1926; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1928 = 6'h8 == _T_340 ? _T_28 : _GEN_1927; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1929 = 6'h9 == _T_340 ? _T_29 : _GEN_1928; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1930 = 6'ha == _T_340 ? _T_30 : _GEN_1929; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1931 = 6'hb == _T_340 ? _T_31 : _GEN_1930; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1932 = 6'hc == _T_340 ? _T_32 : _GEN_1931; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1933 = 6'hd == _T_340 ? _T_33 : _GEN_1932; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1934 = 6'he == _T_340 ? _T_34 : _GEN_1933; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1935 = 6'hf == _T_340 ? _T_35 : _GEN_1934; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1936 = 6'h10 == _T_340 ? _T_36 : _GEN_1935; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1937 = 6'h11 == _T_340 ? _T_37 : _GEN_1936; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1938 = 6'h12 == _T_340 ? _T_38 : _GEN_1937; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1939 = 6'h13 == _T_340 ? _T_39 : _GEN_1938; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1940 = 6'h14 == _T_340 ? _T_40 : _GEN_1939; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1941 = 6'h15 == _T_340 ? _T_41 : _GEN_1940; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1942 = 6'h16 == _T_340 ? _T_42 : _GEN_1941; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1943 = 6'h17 == _T_340 ? _T_43 : _GEN_1942; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1944 = 6'h18 == _T_340 ? _T_44 : _GEN_1943; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1945 = 6'h19 == _T_340 ? _T_45 : _GEN_1944; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1946 = 6'h1a == _T_340 ? _T_46 : _GEN_1945; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1947 = 6'h1b == _T_340 ? _T_47 : _GEN_1946; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1948 = 6'h1c == _T_340 ? _T_48 : _GEN_1947; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1949 = 6'h1d == _T_340 ? _T_49 : _GEN_1948; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1950 = 6'h1e == _T_340 ? _T_50 : _GEN_1949; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1951 = 6'h1f == _T_340 ? _T_51 : _GEN_1950; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1952 = 6'h20 == _T_340 ? _T_52 : _GEN_1951; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1953 = 6'h21 == _T_340 ? _T_53 : _GEN_1952; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1954 = 6'h22 == _T_340 ? _T_54 : _GEN_1953; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1955 = 6'h23 == _T_340 ? _T_55 : _GEN_1954; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1956 = 6'h24 == _T_340 ? _T_56 : _GEN_1955; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1957 = 6'h25 == _T_340 ? _T_57 : _GEN_1956; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1958 = 6'h26 == _T_340 ? _T_58 : _GEN_1957; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1959 = 6'h27 == _T_340 ? _T_59 : _GEN_1958; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1960 = 6'h28 == _T_340 ? _T_60 : _GEN_1959; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1961 = 6'h29 == _T_340 ? _T_61 : _GEN_1960; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1962 = 6'h2a == _T_340 ? _T_62 : _GEN_1961; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1963 = 6'h2b == _T_340 ? _T_63 : _GEN_1962; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1964 = 6'h2c == _T_340 ? _T_64 : _GEN_1963; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1965 = 6'h2d == _T_340 ? _T_65 : _GEN_1964; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1966 = 6'h2e == _T_340 ? _T_66 : _GEN_1965; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1967 = 6'h2f == _T_340 ? _T_67 : _GEN_1966; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1968 = 6'h30 == _T_340 ? _T_68 : _GEN_1967; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1969 = 6'h31 == _T_340 ? _T_69 : _GEN_1968; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1970 = 6'h32 == _T_340 ? _T_70 : _GEN_1969; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1971 = 6'h33 == _T_340 ? _T_71 : _GEN_1970; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1972 = 6'h34 == _T_340 ? _T_72 : _GEN_1971; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1973 = 6'h35 == _T_340 ? _T_73 : _GEN_1972; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1974 = 6'h36 == _T_340 ? _T_74 : _GEN_1973; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1975 = 6'h37 == _T_340 ? _T_75 : _GEN_1974; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1976 = 6'h38 == _T_340 ? _T_76 : _GEN_1975; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1977 = 6'h39 == _T_340 ? _T_77 : _GEN_1976; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1978 = 6'h3a == _T_340 ? _T_78 : _GEN_1977; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1979 = 6'h3b == _T_340 ? _T_79 : _GEN_1978; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1980 = 6'h3c == _T_340 ? _T_80 : _GEN_1979; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1981 = 6'h3d == _T_340 ? _T_81 : _GEN_1980; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1982 = 6'h3e == _T_340 ? _T_82 : _GEN_1981; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1983 = 6'h3f == _T_340 ? _T_83 : _GEN_1982; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1985 = 6'h1 == _T_344 ? _T_21 : _T_20; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1986 = 6'h2 == _T_344 ? _T_22 : _GEN_1985; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1987 = 6'h3 == _T_344 ? _T_23 : _GEN_1986; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1988 = 6'h4 == _T_344 ? _T_24 : _GEN_1987; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1989 = 6'h5 == _T_344 ? _T_25 : _GEN_1988; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1990 = 6'h6 == _T_344 ? _T_26 : _GEN_1989; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1991 = 6'h7 == _T_344 ? _T_27 : _GEN_1990; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1992 = 6'h8 == _T_344 ? _T_28 : _GEN_1991; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1993 = 6'h9 == _T_344 ? _T_29 : _GEN_1992; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1994 = 6'ha == _T_344 ? _T_30 : _GEN_1993; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1995 = 6'hb == _T_344 ? _T_31 : _GEN_1994; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1996 = 6'hc == _T_344 ? _T_32 : _GEN_1995; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1997 = 6'hd == _T_344 ? _T_33 : _GEN_1996; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1998 = 6'he == _T_344 ? _T_34 : _GEN_1997; // @[execute.scala 79:10:@1962.4]
  assign _GEN_1999 = 6'hf == _T_344 ? _T_35 : _GEN_1998; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2000 = 6'h10 == _T_344 ? _T_36 : _GEN_1999; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2001 = 6'h11 == _T_344 ? _T_37 : _GEN_2000; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2002 = 6'h12 == _T_344 ? _T_38 : _GEN_2001; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2003 = 6'h13 == _T_344 ? _T_39 : _GEN_2002; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2004 = 6'h14 == _T_344 ? _T_40 : _GEN_2003; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2005 = 6'h15 == _T_344 ? _T_41 : _GEN_2004; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2006 = 6'h16 == _T_344 ? _T_42 : _GEN_2005; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2007 = 6'h17 == _T_344 ? _T_43 : _GEN_2006; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2008 = 6'h18 == _T_344 ? _T_44 : _GEN_2007; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2009 = 6'h19 == _T_344 ? _T_45 : _GEN_2008; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2010 = 6'h1a == _T_344 ? _T_46 : _GEN_2009; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2011 = 6'h1b == _T_344 ? _T_47 : _GEN_2010; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2012 = 6'h1c == _T_344 ? _T_48 : _GEN_2011; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2013 = 6'h1d == _T_344 ? _T_49 : _GEN_2012; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2014 = 6'h1e == _T_344 ? _T_50 : _GEN_2013; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2015 = 6'h1f == _T_344 ? _T_51 : _GEN_2014; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2016 = 6'h20 == _T_344 ? _T_52 : _GEN_2015; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2017 = 6'h21 == _T_344 ? _T_53 : _GEN_2016; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2018 = 6'h22 == _T_344 ? _T_54 : _GEN_2017; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2019 = 6'h23 == _T_344 ? _T_55 : _GEN_2018; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2020 = 6'h24 == _T_344 ? _T_56 : _GEN_2019; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2021 = 6'h25 == _T_344 ? _T_57 : _GEN_2020; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2022 = 6'h26 == _T_344 ? _T_58 : _GEN_2021; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2023 = 6'h27 == _T_344 ? _T_59 : _GEN_2022; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2024 = 6'h28 == _T_344 ? _T_60 : _GEN_2023; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2025 = 6'h29 == _T_344 ? _T_61 : _GEN_2024; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2026 = 6'h2a == _T_344 ? _T_62 : _GEN_2025; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2027 = 6'h2b == _T_344 ? _T_63 : _GEN_2026; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2028 = 6'h2c == _T_344 ? _T_64 : _GEN_2027; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2029 = 6'h2d == _T_344 ? _T_65 : _GEN_2028; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2030 = 6'h2e == _T_344 ? _T_66 : _GEN_2029; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2031 = 6'h2f == _T_344 ? _T_67 : _GEN_2030; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2032 = 6'h30 == _T_344 ? _T_68 : _GEN_2031; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2033 = 6'h31 == _T_344 ? _T_69 : _GEN_2032; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2034 = 6'h32 == _T_344 ? _T_70 : _GEN_2033; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2035 = 6'h33 == _T_344 ? _T_71 : _GEN_2034; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2036 = 6'h34 == _T_344 ? _T_72 : _GEN_2035; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2037 = 6'h35 == _T_344 ? _T_73 : _GEN_2036; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2038 = 6'h36 == _T_344 ? _T_74 : _GEN_2037; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2039 = 6'h37 == _T_344 ? _T_75 : _GEN_2038; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2040 = 6'h38 == _T_344 ? _T_76 : _GEN_2039; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2041 = 6'h39 == _T_344 ? _T_77 : _GEN_2040; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2042 = 6'h3a == _T_344 ? _T_78 : _GEN_2041; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2043 = 6'h3b == _T_344 ? _T_79 : _GEN_2042; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2044 = 6'h3c == _T_344 ? _T_80 : _GEN_2043; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2045 = 6'h3d == _T_344 ? _T_81 : _GEN_2044; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2046 = 6'h3e == _T_344 ? _T_82 : _GEN_2045; // @[execute.scala 79:10:@1962.4]
  assign _GEN_2047 = 6'h3f == _T_344 ? _T_83 : _GEN_2046; // @[execute.scala 79:10:@1962.4]
  assign _T_346 = _T_336 ? _GEN_1983 : _GEN_2047; // @[execute.scala 79:10:@1962.4]
  assign _T_348 = io_amount < 6'h30; // @[execute.scala 79:15:@1963.4]
  assign _T_350 = io_amount - 6'h30; // @[execute.scala 79:37:@1964.4]
  assign _T_351 = $unsigned(_T_350); // @[execute.scala 79:37:@1965.4]
  assign _T_352 = _T_351[5:0]; // @[execute.scala 79:37:@1966.4]
  assign _T_355 = 6'h10 + io_amount; // @[execute.scala 79:60:@1967.4]
  assign _T_356 = 6'h10 + io_amount; // @[execute.scala 79:60:@1968.4]
  assign _GEN_2049 = 6'h1 == _T_352 ? _T_21 : _T_20; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2050 = 6'h2 == _T_352 ? _T_22 : _GEN_2049; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2051 = 6'h3 == _T_352 ? _T_23 : _GEN_2050; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2052 = 6'h4 == _T_352 ? _T_24 : _GEN_2051; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2053 = 6'h5 == _T_352 ? _T_25 : _GEN_2052; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2054 = 6'h6 == _T_352 ? _T_26 : _GEN_2053; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2055 = 6'h7 == _T_352 ? _T_27 : _GEN_2054; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2056 = 6'h8 == _T_352 ? _T_28 : _GEN_2055; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2057 = 6'h9 == _T_352 ? _T_29 : _GEN_2056; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2058 = 6'ha == _T_352 ? _T_30 : _GEN_2057; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2059 = 6'hb == _T_352 ? _T_31 : _GEN_2058; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2060 = 6'hc == _T_352 ? _T_32 : _GEN_2059; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2061 = 6'hd == _T_352 ? _T_33 : _GEN_2060; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2062 = 6'he == _T_352 ? _T_34 : _GEN_2061; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2063 = 6'hf == _T_352 ? _T_35 : _GEN_2062; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2064 = 6'h10 == _T_352 ? _T_36 : _GEN_2063; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2065 = 6'h11 == _T_352 ? _T_37 : _GEN_2064; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2066 = 6'h12 == _T_352 ? _T_38 : _GEN_2065; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2067 = 6'h13 == _T_352 ? _T_39 : _GEN_2066; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2068 = 6'h14 == _T_352 ? _T_40 : _GEN_2067; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2069 = 6'h15 == _T_352 ? _T_41 : _GEN_2068; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2070 = 6'h16 == _T_352 ? _T_42 : _GEN_2069; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2071 = 6'h17 == _T_352 ? _T_43 : _GEN_2070; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2072 = 6'h18 == _T_352 ? _T_44 : _GEN_2071; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2073 = 6'h19 == _T_352 ? _T_45 : _GEN_2072; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2074 = 6'h1a == _T_352 ? _T_46 : _GEN_2073; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2075 = 6'h1b == _T_352 ? _T_47 : _GEN_2074; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2076 = 6'h1c == _T_352 ? _T_48 : _GEN_2075; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2077 = 6'h1d == _T_352 ? _T_49 : _GEN_2076; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2078 = 6'h1e == _T_352 ? _T_50 : _GEN_2077; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2079 = 6'h1f == _T_352 ? _T_51 : _GEN_2078; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2080 = 6'h20 == _T_352 ? _T_52 : _GEN_2079; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2081 = 6'h21 == _T_352 ? _T_53 : _GEN_2080; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2082 = 6'h22 == _T_352 ? _T_54 : _GEN_2081; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2083 = 6'h23 == _T_352 ? _T_55 : _GEN_2082; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2084 = 6'h24 == _T_352 ? _T_56 : _GEN_2083; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2085 = 6'h25 == _T_352 ? _T_57 : _GEN_2084; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2086 = 6'h26 == _T_352 ? _T_58 : _GEN_2085; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2087 = 6'h27 == _T_352 ? _T_59 : _GEN_2086; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2088 = 6'h28 == _T_352 ? _T_60 : _GEN_2087; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2089 = 6'h29 == _T_352 ? _T_61 : _GEN_2088; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2090 = 6'h2a == _T_352 ? _T_62 : _GEN_2089; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2091 = 6'h2b == _T_352 ? _T_63 : _GEN_2090; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2092 = 6'h2c == _T_352 ? _T_64 : _GEN_2091; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2093 = 6'h2d == _T_352 ? _T_65 : _GEN_2092; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2094 = 6'h2e == _T_352 ? _T_66 : _GEN_2093; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2095 = 6'h2f == _T_352 ? _T_67 : _GEN_2094; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2096 = 6'h30 == _T_352 ? _T_68 : _GEN_2095; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2097 = 6'h31 == _T_352 ? _T_69 : _GEN_2096; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2098 = 6'h32 == _T_352 ? _T_70 : _GEN_2097; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2099 = 6'h33 == _T_352 ? _T_71 : _GEN_2098; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2100 = 6'h34 == _T_352 ? _T_72 : _GEN_2099; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2101 = 6'h35 == _T_352 ? _T_73 : _GEN_2100; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2102 = 6'h36 == _T_352 ? _T_74 : _GEN_2101; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2103 = 6'h37 == _T_352 ? _T_75 : _GEN_2102; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2104 = 6'h38 == _T_352 ? _T_76 : _GEN_2103; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2105 = 6'h39 == _T_352 ? _T_77 : _GEN_2104; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2106 = 6'h3a == _T_352 ? _T_78 : _GEN_2105; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2107 = 6'h3b == _T_352 ? _T_79 : _GEN_2106; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2108 = 6'h3c == _T_352 ? _T_80 : _GEN_2107; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2109 = 6'h3d == _T_352 ? _T_81 : _GEN_2108; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2110 = 6'h3e == _T_352 ? _T_82 : _GEN_2109; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2111 = 6'h3f == _T_352 ? _T_83 : _GEN_2110; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2113 = 6'h1 == _T_356 ? _T_21 : _T_20; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2114 = 6'h2 == _T_356 ? _T_22 : _GEN_2113; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2115 = 6'h3 == _T_356 ? _T_23 : _GEN_2114; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2116 = 6'h4 == _T_356 ? _T_24 : _GEN_2115; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2117 = 6'h5 == _T_356 ? _T_25 : _GEN_2116; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2118 = 6'h6 == _T_356 ? _T_26 : _GEN_2117; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2119 = 6'h7 == _T_356 ? _T_27 : _GEN_2118; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2120 = 6'h8 == _T_356 ? _T_28 : _GEN_2119; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2121 = 6'h9 == _T_356 ? _T_29 : _GEN_2120; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2122 = 6'ha == _T_356 ? _T_30 : _GEN_2121; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2123 = 6'hb == _T_356 ? _T_31 : _GEN_2122; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2124 = 6'hc == _T_356 ? _T_32 : _GEN_2123; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2125 = 6'hd == _T_356 ? _T_33 : _GEN_2124; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2126 = 6'he == _T_356 ? _T_34 : _GEN_2125; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2127 = 6'hf == _T_356 ? _T_35 : _GEN_2126; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2128 = 6'h10 == _T_356 ? _T_36 : _GEN_2127; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2129 = 6'h11 == _T_356 ? _T_37 : _GEN_2128; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2130 = 6'h12 == _T_356 ? _T_38 : _GEN_2129; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2131 = 6'h13 == _T_356 ? _T_39 : _GEN_2130; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2132 = 6'h14 == _T_356 ? _T_40 : _GEN_2131; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2133 = 6'h15 == _T_356 ? _T_41 : _GEN_2132; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2134 = 6'h16 == _T_356 ? _T_42 : _GEN_2133; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2135 = 6'h17 == _T_356 ? _T_43 : _GEN_2134; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2136 = 6'h18 == _T_356 ? _T_44 : _GEN_2135; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2137 = 6'h19 == _T_356 ? _T_45 : _GEN_2136; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2138 = 6'h1a == _T_356 ? _T_46 : _GEN_2137; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2139 = 6'h1b == _T_356 ? _T_47 : _GEN_2138; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2140 = 6'h1c == _T_356 ? _T_48 : _GEN_2139; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2141 = 6'h1d == _T_356 ? _T_49 : _GEN_2140; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2142 = 6'h1e == _T_356 ? _T_50 : _GEN_2141; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2143 = 6'h1f == _T_356 ? _T_51 : _GEN_2142; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2144 = 6'h20 == _T_356 ? _T_52 : _GEN_2143; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2145 = 6'h21 == _T_356 ? _T_53 : _GEN_2144; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2146 = 6'h22 == _T_356 ? _T_54 : _GEN_2145; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2147 = 6'h23 == _T_356 ? _T_55 : _GEN_2146; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2148 = 6'h24 == _T_356 ? _T_56 : _GEN_2147; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2149 = 6'h25 == _T_356 ? _T_57 : _GEN_2148; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2150 = 6'h26 == _T_356 ? _T_58 : _GEN_2149; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2151 = 6'h27 == _T_356 ? _T_59 : _GEN_2150; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2152 = 6'h28 == _T_356 ? _T_60 : _GEN_2151; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2153 = 6'h29 == _T_356 ? _T_61 : _GEN_2152; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2154 = 6'h2a == _T_356 ? _T_62 : _GEN_2153; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2155 = 6'h2b == _T_356 ? _T_63 : _GEN_2154; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2156 = 6'h2c == _T_356 ? _T_64 : _GEN_2155; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2157 = 6'h2d == _T_356 ? _T_65 : _GEN_2156; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2158 = 6'h2e == _T_356 ? _T_66 : _GEN_2157; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2159 = 6'h2f == _T_356 ? _T_67 : _GEN_2158; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2160 = 6'h30 == _T_356 ? _T_68 : _GEN_2159; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2161 = 6'h31 == _T_356 ? _T_69 : _GEN_2160; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2162 = 6'h32 == _T_356 ? _T_70 : _GEN_2161; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2163 = 6'h33 == _T_356 ? _T_71 : _GEN_2162; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2164 = 6'h34 == _T_356 ? _T_72 : _GEN_2163; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2165 = 6'h35 == _T_356 ? _T_73 : _GEN_2164; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2166 = 6'h36 == _T_356 ? _T_74 : _GEN_2165; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2167 = 6'h37 == _T_356 ? _T_75 : _GEN_2166; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2168 = 6'h38 == _T_356 ? _T_76 : _GEN_2167; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2169 = 6'h39 == _T_356 ? _T_77 : _GEN_2168; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2170 = 6'h3a == _T_356 ? _T_78 : _GEN_2169; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2171 = 6'h3b == _T_356 ? _T_79 : _GEN_2170; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2172 = 6'h3c == _T_356 ? _T_80 : _GEN_2171; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2173 = 6'h3d == _T_356 ? _T_81 : _GEN_2172; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2174 = 6'h3e == _T_356 ? _T_82 : _GEN_2173; // @[execute.scala 79:10:@1969.4]
  assign _GEN_2175 = 6'h3f == _T_356 ? _T_83 : _GEN_2174; // @[execute.scala 79:10:@1969.4]
  assign _T_358 = _T_348 ? _GEN_2111 : _GEN_2175; // @[execute.scala 79:10:@1969.4]
  assign _T_360 = io_amount < 6'h2f; // @[execute.scala 79:15:@1970.4]
  assign _T_362 = io_amount - 6'h2f; // @[execute.scala 79:37:@1971.4]
  assign _T_363 = $unsigned(_T_362); // @[execute.scala 79:37:@1972.4]
  assign _T_364 = _T_363[5:0]; // @[execute.scala 79:37:@1973.4]
  assign _T_367 = 6'h11 + io_amount; // @[execute.scala 79:60:@1974.4]
  assign _T_368 = 6'h11 + io_amount; // @[execute.scala 79:60:@1975.4]
  assign _GEN_2177 = 6'h1 == _T_364 ? _T_21 : _T_20; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2178 = 6'h2 == _T_364 ? _T_22 : _GEN_2177; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2179 = 6'h3 == _T_364 ? _T_23 : _GEN_2178; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2180 = 6'h4 == _T_364 ? _T_24 : _GEN_2179; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2181 = 6'h5 == _T_364 ? _T_25 : _GEN_2180; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2182 = 6'h6 == _T_364 ? _T_26 : _GEN_2181; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2183 = 6'h7 == _T_364 ? _T_27 : _GEN_2182; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2184 = 6'h8 == _T_364 ? _T_28 : _GEN_2183; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2185 = 6'h9 == _T_364 ? _T_29 : _GEN_2184; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2186 = 6'ha == _T_364 ? _T_30 : _GEN_2185; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2187 = 6'hb == _T_364 ? _T_31 : _GEN_2186; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2188 = 6'hc == _T_364 ? _T_32 : _GEN_2187; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2189 = 6'hd == _T_364 ? _T_33 : _GEN_2188; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2190 = 6'he == _T_364 ? _T_34 : _GEN_2189; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2191 = 6'hf == _T_364 ? _T_35 : _GEN_2190; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2192 = 6'h10 == _T_364 ? _T_36 : _GEN_2191; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2193 = 6'h11 == _T_364 ? _T_37 : _GEN_2192; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2194 = 6'h12 == _T_364 ? _T_38 : _GEN_2193; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2195 = 6'h13 == _T_364 ? _T_39 : _GEN_2194; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2196 = 6'h14 == _T_364 ? _T_40 : _GEN_2195; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2197 = 6'h15 == _T_364 ? _T_41 : _GEN_2196; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2198 = 6'h16 == _T_364 ? _T_42 : _GEN_2197; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2199 = 6'h17 == _T_364 ? _T_43 : _GEN_2198; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2200 = 6'h18 == _T_364 ? _T_44 : _GEN_2199; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2201 = 6'h19 == _T_364 ? _T_45 : _GEN_2200; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2202 = 6'h1a == _T_364 ? _T_46 : _GEN_2201; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2203 = 6'h1b == _T_364 ? _T_47 : _GEN_2202; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2204 = 6'h1c == _T_364 ? _T_48 : _GEN_2203; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2205 = 6'h1d == _T_364 ? _T_49 : _GEN_2204; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2206 = 6'h1e == _T_364 ? _T_50 : _GEN_2205; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2207 = 6'h1f == _T_364 ? _T_51 : _GEN_2206; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2208 = 6'h20 == _T_364 ? _T_52 : _GEN_2207; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2209 = 6'h21 == _T_364 ? _T_53 : _GEN_2208; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2210 = 6'h22 == _T_364 ? _T_54 : _GEN_2209; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2211 = 6'h23 == _T_364 ? _T_55 : _GEN_2210; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2212 = 6'h24 == _T_364 ? _T_56 : _GEN_2211; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2213 = 6'h25 == _T_364 ? _T_57 : _GEN_2212; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2214 = 6'h26 == _T_364 ? _T_58 : _GEN_2213; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2215 = 6'h27 == _T_364 ? _T_59 : _GEN_2214; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2216 = 6'h28 == _T_364 ? _T_60 : _GEN_2215; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2217 = 6'h29 == _T_364 ? _T_61 : _GEN_2216; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2218 = 6'h2a == _T_364 ? _T_62 : _GEN_2217; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2219 = 6'h2b == _T_364 ? _T_63 : _GEN_2218; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2220 = 6'h2c == _T_364 ? _T_64 : _GEN_2219; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2221 = 6'h2d == _T_364 ? _T_65 : _GEN_2220; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2222 = 6'h2e == _T_364 ? _T_66 : _GEN_2221; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2223 = 6'h2f == _T_364 ? _T_67 : _GEN_2222; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2224 = 6'h30 == _T_364 ? _T_68 : _GEN_2223; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2225 = 6'h31 == _T_364 ? _T_69 : _GEN_2224; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2226 = 6'h32 == _T_364 ? _T_70 : _GEN_2225; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2227 = 6'h33 == _T_364 ? _T_71 : _GEN_2226; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2228 = 6'h34 == _T_364 ? _T_72 : _GEN_2227; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2229 = 6'h35 == _T_364 ? _T_73 : _GEN_2228; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2230 = 6'h36 == _T_364 ? _T_74 : _GEN_2229; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2231 = 6'h37 == _T_364 ? _T_75 : _GEN_2230; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2232 = 6'h38 == _T_364 ? _T_76 : _GEN_2231; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2233 = 6'h39 == _T_364 ? _T_77 : _GEN_2232; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2234 = 6'h3a == _T_364 ? _T_78 : _GEN_2233; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2235 = 6'h3b == _T_364 ? _T_79 : _GEN_2234; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2236 = 6'h3c == _T_364 ? _T_80 : _GEN_2235; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2237 = 6'h3d == _T_364 ? _T_81 : _GEN_2236; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2238 = 6'h3e == _T_364 ? _T_82 : _GEN_2237; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2239 = 6'h3f == _T_364 ? _T_83 : _GEN_2238; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2241 = 6'h1 == _T_368 ? _T_21 : _T_20; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2242 = 6'h2 == _T_368 ? _T_22 : _GEN_2241; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2243 = 6'h3 == _T_368 ? _T_23 : _GEN_2242; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2244 = 6'h4 == _T_368 ? _T_24 : _GEN_2243; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2245 = 6'h5 == _T_368 ? _T_25 : _GEN_2244; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2246 = 6'h6 == _T_368 ? _T_26 : _GEN_2245; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2247 = 6'h7 == _T_368 ? _T_27 : _GEN_2246; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2248 = 6'h8 == _T_368 ? _T_28 : _GEN_2247; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2249 = 6'h9 == _T_368 ? _T_29 : _GEN_2248; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2250 = 6'ha == _T_368 ? _T_30 : _GEN_2249; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2251 = 6'hb == _T_368 ? _T_31 : _GEN_2250; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2252 = 6'hc == _T_368 ? _T_32 : _GEN_2251; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2253 = 6'hd == _T_368 ? _T_33 : _GEN_2252; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2254 = 6'he == _T_368 ? _T_34 : _GEN_2253; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2255 = 6'hf == _T_368 ? _T_35 : _GEN_2254; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2256 = 6'h10 == _T_368 ? _T_36 : _GEN_2255; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2257 = 6'h11 == _T_368 ? _T_37 : _GEN_2256; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2258 = 6'h12 == _T_368 ? _T_38 : _GEN_2257; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2259 = 6'h13 == _T_368 ? _T_39 : _GEN_2258; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2260 = 6'h14 == _T_368 ? _T_40 : _GEN_2259; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2261 = 6'h15 == _T_368 ? _T_41 : _GEN_2260; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2262 = 6'h16 == _T_368 ? _T_42 : _GEN_2261; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2263 = 6'h17 == _T_368 ? _T_43 : _GEN_2262; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2264 = 6'h18 == _T_368 ? _T_44 : _GEN_2263; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2265 = 6'h19 == _T_368 ? _T_45 : _GEN_2264; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2266 = 6'h1a == _T_368 ? _T_46 : _GEN_2265; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2267 = 6'h1b == _T_368 ? _T_47 : _GEN_2266; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2268 = 6'h1c == _T_368 ? _T_48 : _GEN_2267; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2269 = 6'h1d == _T_368 ? _T_49 : _GEN_2268; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2270 = 6'h1e == _T_368 ? _T_50 : _GEN_2269; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2271 = 6'h1f == _T_368 ? _T_51 : _GEN_2270; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2272 = 6'h20 == _T_368 ? _T_52 : _GEN_2271; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2273 = 6'h21 == _T_368 ? _T_53 : _GEN_2272; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2274 = 6'h22 == _T_368 ? _T_54 : _GEN_2273; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2275 = 6'h23 == _T_368 ? _T_55 : _GEN_2274; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2276 = 6'h24 == _T_368 ? _T_56 : _GEN_2275; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2277 = 6'h25 == _T_368 ? _T_57 : _GEN_2276; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2278 = 6'h26 == _T_368 ? _T_58 : _GEN_2277; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2279 = 6'h27 == _T_368 ? _T_59 : _GEN_2278; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2280 = 6'h28 == _T_368 ? _T_60 : _GEN_2279; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2281 = 6'h29 == _T_368 ? _T_61 : _GEN_2280; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2282 = 6'h2a == _T_368 ? _T_62 : _GEN_2281; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2283 = 6'h2b == _T_368 ? _T_63 : _GEN_2282; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2284 = 6'h2c == _T_368 ? _T_64 : _GEN_2283; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2285 = 6'h2d == _T_368 ? _T_65 : _GEN_2284; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2286 = 6'h2e == _T_368 ? _T_66 : _GEN_2285; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2287 = 6'h2f == _T_368 ? _T_67 : _GEN_2286; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2288 = 6'h30 == _T_368 ? _T_68 : _GEN_2287; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2289 = 6'h31 == _T_368 ? _T_69 : _GEN_2288; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2290 = 6'h32 == _T_368 ? _T_70 : _GEN_2289; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2291 = 6'h33 == _T_368 ? _T_71 : _GEN_2290; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2292 = 6'h34 == _T_368 ? _T_72 : _GEN_2291; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2293 = 6'h35 == _T_368 ? _T_73 : _GEN_2292; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2294 = 6'h36 == _T_368 ? _T_74 : _GEN_2293; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2295 = 6'h37 == _T_368 ? _T_75 : _GEN_2294; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2296 = 6'h38 == _T_368 ? _T_76 : _GEN_2295; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2297 = 6'h39 == _T_368 ? _T_77 : _GEN_2296; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2298 = 6'h3a == _T_368 ? _T_78 : _GEN_2297; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2299 = 6'h3b == _T_368 ? _T_79 : _GEN_2298; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2300 = 6'h3c == _T_368 ? _T_80 : _GEN_2299; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2301 = 6'h3d == _T_368 ? _T_81 : _GEN_2300; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2302 = 6'h3e == _T_368 ? _T_82 : _GEN_2301; // @[execute.scala 79:10:@1976.4]
  assign _GEN_2303 = 6'h3f == _T_368 ? _T_83 : _GEN_2302; // @[execute.scala 79:10:@1976.4]
  assign _T_370 = _T_360 ? _GEN_2239 : _GEN_2303; // @[execute.scala 79:10:@1976.4]
  assign _T_372 = io_amount < 6'h2e; // @[execute.scala 79:15:@1977.4]
  assign _T_374 = io_amount - 6'h2e; // @[execute.scala 79:37:@1978.4]
  assign _T_375 = $unsigned(_T_374); // @[execute.scala 79:37:@1979.4]
  assign _T_376 = _T_375[5:0]; // @[execute.scala 79:37:@1980.4]
  assign _T_379 = 6'h12 + io_amount; // @[execute.scala 79:60:@1981.4]
  assign _T_380 = 6'h12 + io_amount; // @[execute.scala 79:60:@1982.4]
  assign _GEN_2305 = 6'h1 == _T_376 ? _T_21 : _T_20; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2306 = 6'h2 == _T_376 ? _T_22 : _GEN_2305; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2307 = 6'h3 == _T_376 ? _T_23 : _GEN_2306; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2308 = 6'h4 == _T_376 ? _T_24 : _GEN_2307; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2309 = 6'h5 == _T_376 ? _T_25 : _GEN_2308; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2310 = 6'h6 == _T_376 ? _T_26 : _GEN_2309; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2311 = 6'h7 == _T_376 ? _T_27 : _GEN_2310; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2312 = 6'h8 == _T_376 ? _T_28 : _GEN_2311; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2313 = 6'h9 == _T_376 ? _T_29 : _GEN_2312; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2314 = 6'ha == _T_376 ? _T_30 : _GEN_2313; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2315 = 6'hb == _T_376 ? _T_31 : _GEN_2314; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2316 = 6'hc == _T_376 ? _T_32 : _GEN_2315; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2317 = 6'hd == _T_376 ? _T_33 : _GEN_2316; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2318 = 6'he == _T_376 ? _T_34 : _GEN_2317; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2319 = 6'hf == _T_376 ? _T_35 : _GEN_2318; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2320 = 6'h10 == _T_376 ? _T_36 : _GEN_2319; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2321 = 6'h11 == _T_376 ? _T_37 : _GEN_2320; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2322 = 6'h12 == _T_376 ? _T_38 : _GEN_2321; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2323 = 6'h13 == _T_376 ? _T_39 : _GEN_2322; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2324 = 6'h14 == _T_376 ? _T_40 : _GEN_2323; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2325 = 6'h15 == _T_376 ? _T_41 : _GEN_2324; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2326 = 6'h16 == _T_376 ? _T_42 : _GEN_2325; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2327 = 6'h17 == _T_376 ? _T_43 : _GEN_2326; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2328 = 6'h18 == _T_376 ? _T_44 : _GEN_2327; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2329 = 6'h19 == _T_376 ? _T_45 : _GEN_2328; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2330 = 6'h1a == _T_376 ? _T_46 : _GEN_2329; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2331 = 6'h1b == _T_376 ? _T_47 : _GEN_2330; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2332 = 6'h1c == _T_376 ? _T_48 : _GEN_2331; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2333 = 6'h1d == _T_376 ? _T_49 : _GEN_2332; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2334 = 6'h1e == _T_376 ? _T_50 : _GEN_2333; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2335 = 6'h1f == _T_376 ? _T_51 : _GEN_2334; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2336 = 6'h20 == _T_376 ? _T_52 : _GEN_2335; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2337 = 6'h21 == _T_376 ? _T_53 : _GEN_2336; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2338 = 6'h22 == _T_376 ? _T_54 : _GEN_2337; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2339 = 6'h23 == _T_376 ? _T_55 : _GEN_2338; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2340 = 6'h24 == _T_376 ? _T_56 : _GEN_2339; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2341 = 6'h25 == _T_376 ? _T_57 : _GEN_2340; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2342 = 6'h26 == _T_376 ? _T_58 : _GEN_2341; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2343 = 6'h27 == _T_376 ? _T_59 : _GEN_2342; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2344 = 6'h28 == _T_376 ? _T_60 : _GEN_2343; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2345 = 6'h29 == _T_376 ? _T_61 : _GEN_2344; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2346 = 6'h2a == _T_376 ? _T_62 : _GEN_2345; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2347 = 6'h2b == _T_376 ? _T_63 : _GEN_2346; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2348 = 6'h2c == _T_376 ? _T_64 : _GEN_2347; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2349 = 6'h2d == _T_376 ? _T_65 : _GEN_2348; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2350 = 6'h2e == _T_376 ? _T_66 : _GEN_2349; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2351 = 6'h2f == _T_376 ? _T_67 : _GEN_2350; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2352 = 6'h30 == _T_376 ? _T_68 : _GEN_2351; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2353 = 6'h31 == _T_376 ? _T_69 : _GEN_2352; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2354 = 6'h32 == _T_376 ? _T_70 : _GEN_2353; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2355 = 6'h33 == _T_376 ? _T_71 : _GEN_2354; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2356 = 6'h34 == _T_376 ? _T_72 : _GEN_2355; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2357 = 6'h35 == _T_376 ? _T_73 : _GEN_2356; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2358 = 6'h36 == _T_376 ? _T_74 : _GEN_2357; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2359 = 6'h37 == _T_376 ? _T_75 : _GEN_2358; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2360 = 6'h38 == _T_376 ? _T_76 : _GEN_2359; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2361 = 6'h39 == _T_376 ? _T_77 : _GEN_2360; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2362 = 6'h3a == _T_376 ? _T_78 : _GEN_2361; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2363 = 6'h3b == _T_376 ? _T_79 : _GEN_2362; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2364 = 6'h3c == _T_376 ? _T_80 : _GEN_2363; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2365 = 6'h3d == _T_376 ? _T_81 : _GEN_2364; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2366 = 6'h3e == _T_376 ? _T_82 : _GEN_2365; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2367 = 6'h3f == _T_376 ? _T_83 : _GEN_2366; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2369 = 6'h1 == _T_380 ? _T_21 : _T_20; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2370 = 6'h2 == _T_380 ? _T_22 : _GEN_2369; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2371 = 6'h3 == _T_380 ? _T_23 : _GEN_2370; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2372 = 6'h4 == _T_380 ? _T_24 : _GEN_2371; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2373 = 6'h5 == _T_380 ? _T_25 : _GEN_2372; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2374 = 6'h6 == _T_380 ? _T_26 : _GEN_2373; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2375 = 6'h7 == _T_380 ? _T_27 : _GEN_2374; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2376 = 6'h8 == _T_380 ? _T_28 : _GEN_2375; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2377 = 6'h9 == _T_380 ? _T_29 : _GEN_2376; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2378 = 6'ha == _T_380 ? _T_30 : _GEN_2377; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2379 = 6'hb == _T_380 ? _T_31 : _GEN_2378; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2380 = 6'hc == _T_380 ? _T_32 : _GEN_2379; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2381 = 6'hd == _T_380 ? _T_33 : _GEN_2380; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2382 = 6'he == _T_380 ? _T_34 : _GEN_2381; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2383 = 6'hf == _T_380 ? _T_35 : _GEN_2382; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2384 = 6'h10 == _T_380 ? _T_36 : _GEN_2383; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2385 = 6'h11 == _T_380 ? _T_37 : _GEN_2384; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2386 = 6'h12 == _T_380 ? _T_38 : _GEN_2385; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2387 = 6'h13 == _T_380 ? _T_39 : _GEN_2386; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2388 = 6'h14 == _T_380 ? _T_40 : _GEN_2387; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2389 = 6'h15 == _T_380 ? _T_41 : _GEN_2388; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2390 = 6'h16 == _T_380 ? _T_42 : _GEN_2389; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2391 = 6'h17 == _T_380 ? _T_43 : _GEN_2390; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2392 = 6'h18 == _T_380 ? _T_44 : _GEN_2391; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2393 = 6'h19 == _T_380 ? _T_45 : _GEN_2392; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2394 = 6'h1a == _T_380 ? _T_46 : _GEN_2393; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2395 = 6'h1b == _T_380 ? _T_47 : _GEN_2394; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2396 = 6'h1c == _T_380 ? _T_48 : _GEN_2395; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2397 = 6'h1d == _T_380 ? _T_49 : _GEN_2396; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2398 = 6'h1e == _T_380 ? _T_50 : _GEN_2397; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2399 = 6'h1f == _T_380 ? _T_51 : _GEN_2398; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2400 = 6'h20 == _T_380 ? _T_52 : _GEN_2399; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2401 = 6'h21 == _T_380 ? _T_53 : _GEN_2400; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2402 = 6'h22 == _T_380 ? _T_54 : _GEN_2401; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2403 = 6'h23 == _T_380 ? _T_55 : _GEN_2402; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2404 = 6'h24 == _T_380 ? _T_56 : _GEN_2403; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2405 = 6'h25 == _T_380 ? _T_57 : _GEN_2404; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2406 = 6'h26 == _T_380 ? _T_58 : _GEN_2405; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2407 = 6'h27 == _T_380 ? _T_59 : _GEN_2406; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2408 = 6'h28 == _T_380 ? _T_60 : _GEN_2407; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2409 = 6'h29 == _T_380 ? _T_61 : _GEN_2408; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2410 = 6'h2a == _T_380 ? _T_62 : _GEN_2409; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2411 = 6'h2b == _T_380 ? _T_63 : _GEN_2410; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2412 = 6'h2c == _T_380 ? _T_64 : _GEN_2411; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2413 = 6'h2d == _T_380 ? _T_65 : _GEN_2412; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2414 = 6'h2e == _T_380 ? _T_66 : _GEN_2413; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2415 = 6'h2f == _T_380 ? _T_67 : _GEN_2414; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2416 = 6'h30 == _T_380 ? _T_68 : _GEN_2415; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2417 = 6'h31 == _T_380 ? _T_69 : _GEN_2416; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2418 = 6'h32 == _T_380 ? _T_70 : _GEN_2417; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2419 = 6'h33 == _T_380 ? _T_71 : _GEN_2418; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2420 = 6'h34 == _T_380 ? _T_72 : _GEN_2419; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2421 = 6'h35 == _T_380 ? _T_73 : _GEN_2420; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2422 = 6'h36 == _T_380 ? _T_74 : _GEN_2421; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2423 = 6'h37 == _T_380 ? _T_75 : _GEN_2422; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2424 = 6'h38 == _T_380 ? _T_76 : _GEN_2423; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2425 = 6'h39 == _T_380 ? _T_77 : _GEN_2424; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2426 = 6'h3a == _T_380 ? _T_78 : _GEN_2425; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2427 = 6'h3b == _T_380 ? _T_79 : _GEN_2426; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2428 = 6'h3c == _T_380 ? _T_80 : _GEN_2427; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2429 = 6'h3d == _T_380 ? _T_81 : _GEN_2428; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2430 = 6'h3e == _T_380 ? _T_82 : _GEN_2429; // @[execute.scala 79:10:@1983.4]
  assign _GEN_2431 = 6'h3f == _T_380 ? _T_83 : _GEN_2430; // @[execute.scala 79:10:@1983.4]
  assign _T_382 = _T_372 ? _GEN_2367 : _GEN_2431; // @[execute.scala 79:10:@1983.4]
  assign _T_384 = io_amount < 6'h2d; // @[execute.scala 79:15:@1984.4]
  assign _T_386 = io_amount - 6'h2d; // @[execute.scala 79:37:@1985.4]
  assign _T_387 = $unsigned(_T_386); // @[execute.scala 79:37:@1986.4]
  assign _T_388 = _T_387[5:0]; // @[execute.scala 79:37:@1987.4]
  assign _T_391 = 6'h13 + io_amount; // @[execute.scala 79:60:@1988.4]
  assign _T_392 = 6'h13 + io_amount; // @[execute.scala 79:60:@1989.4]
  assign _GEN_2433 = 6'h1 == _T_388 ? _T_21 : _T_20; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2434 = 6'h2 == _T_388 ? _T_22 : _GEN_2433; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2435 = 6'h3 == _T_388 ? _T_23 : _GEN_2434; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2436 = 6'h4 == _T_388 ? _T_24 : _GEN_2435; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2437 = 6'h5 == _T_388 ? _T_25 : _GEN_2436; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2438 = 6'h6 == _T_388 ? _T_26 : _GEN_2437; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2439 = 6'h7 == _T_388 ? _T_27 : _GEN_2438; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2440 = 6'h8 == _T_388 ? _T_28 : _GEN_2439; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2441 = 6'h9 == _T_388 ? _T_29 : _GEN_2440; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2442 = 6'ha == _T_388 ? _T_30 : _GEN_2441; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2443 = 6'hb == _T_388 ? _T_31 : _GEN_2442; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2444 = 6'hc == _T_388 ? _T_32 : _GEN_2443; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2445 = 6'hd == _T_388 ? _T_33 : _GEN_2444; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2446 = 6'he == _T_388 ? _T_34 : _GEN_2445; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2447 = 6'hf == _T_388 ? _T_35 : _GEN_2446; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2448 = 6'h10 == _T_388 ? _T_36 : _GEN_2447; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2449 = 6'h11 == _T_388 ? _T_37 : _GEN_2448; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2450 = 6'h12 == _T_388 ? _T_38 : _GEN_2449; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2451 = 6'h13 == _T_388 ? _T_39 : _GEN_2450; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2452 = 6'h14 == _T_388 ? _T_40 : _GEN_2451; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2453 = 6'h15 == _T_388 ? _T_41 : _GEN_2452; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2454 = 6'h16 == _T_388 ? _T_42 : _GEN_2453; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2455 = 6'h17 == _T_388 ? _T_43 : _GEN_2454; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2456 = 6'h18 == _T_388 ? _T_44 : _GEN_2455; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2457 = 6'h19 == _T_388 ? _T_45 : _GEN_2456; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2458 = 6'h1a == _T_388 ? _T_46 : _GEN_2457; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2459 = 6'h1b == _T_388 ? _T_47 : _GEN_2458; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2460 = 6'h1c == _T_388 ? _T_48 : _GEN_2459; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2461 = 6'h1d == _T_388 ? _T_49 : _GEN_2460; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2462 = 6'h1e == _T_388 ? _T_50 : _GEN_2461; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2463 = 6'h1f == _T_388 ? _T_51 : _GEN_2462; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2464 = 6'h20 == _T_388 ? _T_52 : _GEN_2463; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2465 = 6'h21 == _T_388 ? _T_53 : _GEN_2464; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2466 = 6'h22 == _T_388 ? _T_54 : _GEN_2465; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2467 = 6'h23 == _T_388 ? _T_55 : _GEN_2466; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2468 = 6'h24 == _T_388 ? _T_56 : _GEN_2467; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2469 = 6'h25 == _T_388 ? _T_57 : _GEN_2468; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2470 = 6'h26 == _T_388 ? _T_58 : _GEN_2469; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2471 = 6'h27 == _T_388 ? _T_59 : _GEN_2470; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2472 = 6'h28 == _T_388 ? _T_60 : _GEN_2471; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2473 = 6'h29 == _T_388 ? _T_61 : _GEN_2472; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2474 = 6'h2a == _T_388 ? _T_62 : _GEN_2473; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2475 = 6'h2b == _T_388 ? _T_63 : _GEN_2474; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2476 = 6'h2c == _T_388 ? _T_64 : _GEN_2475; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2477 = 6'h2d == _T_388 ? _T_65 : _GEN_2476; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2478 = 6'h2e == _T_388 ? _T_66 : _GEN_2477; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2479 = 6'h2f == _T_388 ? _T_67 : _GEN_2478; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2480 = 6'h30 == _T_388 ? _T_68 : _GEN_2479; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2481 = 6'h31 == _T_388 ? _T_69 : _GEN_2480; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2482 = 6'h32 == _T_388 ? _T_70 : _GEN_2481; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2483 = 6'h33 == _T_388 ? _T_71 : _GEN_2482; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2484 = 6'h34 == _T_388 ? _T_72 : _GEN_2483; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2485 = 6'h35 == _T_388 ? _T_73 : _GEN_2484; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2486 = 6'h36 == _T_388 ? _T_74 : _GEN_2485; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2487 = 6'h37 == _T_388 ? _T_75 : _GEN_2486; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2488 = 6'h38 == _T_388 ? _T_76 : _GEN_2487; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2489 = 6'h39 == _T_388 ? _T_77 : _GEN_2488; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2490 = 6'h3a == _T_388 ? _T_78 : _GEN_2489; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2491 = 6'h3b == _T_388 ? _T_79 : _GEN_2490; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2492 = 6'h3c == _T_388 ? _T_80 : _GEN_2491; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2493 = 6'h3d == _T_388 ? _T_81 : _GEN_2492; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2494 = 6'h3e == _T_388 ? _T_82 : _GEN_2493; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2495 = 6'h3f == _T_388 ? _T_83 : _GEN_2494; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2497 = 6'h1 == _T_392 ? _T_21 : _T_20; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2498 = 6'h2 == _T_392 ? _T_22 : _GEN_2497; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2499 = 6'h3 == _T_392 ? _T_23 : _GEN_2498; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2500 = 6'h4 == _T_392 ? _T_24 : _GEN_2499; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2501 = 6'h5 == _T_392 ? _T_25 : _GEN_2500; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2502 = 6'h6 == _T_392 ? _T_26 : _GEN_2501; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2503 = 6'h7 == _T_392 ? _T_27 : _GEN_2502; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2504 = 6'h8 == _T_392 ? _T_28 : _GEN_2503; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2505 = 6'h9 == _T_392 ? _T_29 : _GEN_2504; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2506 = 6'ha == _T_392 ? _T_30 : _GEN_2505; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2507 = 6'hb == _T_392 ? _T_31 : _GEN_2506; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2508 = 6'hc == _T_392 ? _T_32 : _GEN_2507; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2509 = 6'hd == _T_392 ? _T_33 : _GEN_2508; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2510 = 6'he == _T_392 ? _T_34 : _GEN_2509; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2511 = 6'hf == _T_392 ? _T_35 : _GEN_2510; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2512 = 6'h10 == _T_392 ? _T_36 : _GEN_2511; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2513 = 6'h11 == _T_392 ? _T_37 : _GEN_2512; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2514 = 6'h12 == _T_392 ? _T_38 : _GEN_2513; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2515 = 6'h13 == _T_392 ? _T_39 : _GEN_2514; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2516 = 6'h14 == _T_392 ? _T_40 : _GEN_2515; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2517 = 6'h15 == _T_392 ? _T_41 : _GEN_2516; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2518 = 6'h16 == _T_392 ? _T_42 : _GEN_2517; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2519 = 6'h17 == _T_392 ? _T_43 : _GEN_2518; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2520 = 6'h18 == _T_392 ? _T_44 : _GEN_2519; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2521 = 6'h19 == _T_392 ? _T_45 : _GEN_2520; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2522 = 6'h1a == _T_392 ? _T_46 : _GEN_2521; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2523 = 6'h1b == _T_392 ? _T_47 : _GEN_2522; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2524 = 6'h1c == _T_392 ? _T_48 : _GEN_2523; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2525 = 6'h1d == _T_392 ? _T_49 : _GEN_2524; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2526 = 6'h1e == _T_392 ? _T_50 : _GEN_2525; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2527 = 6'h1f == _T_392 ? _T_51 : _GEN_2526; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2528 = 6'h20 == _T_392 ? _T_52 : _GEN_2527; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2529 = 6'h21 == _T_392 ? _T_53 : _GEN_2528; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2530 = 6'h22 == _T_392 ? _T_54 : _GEN_2529; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2531 = 6'h23 == _T_392 ? _T_55 : _GEN_2530; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2532 = 6'h24 == _T_392 ? _T_56 : _GEN_2531; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2533 = 6'h25 == _T_392 ? _T_57 : _GEN_2532; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2534 = 6'h26 == _T_392 ? _T_58 : _GEN_2533; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2535 = 6'h27 == _T_392 ? _T_59 : _GEN_2534; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2536 = 6'h28 == _T_392 ? _T_60 : _GEN_2535; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2537 = 6'h29 == _T_392 ? _T_61 : _GEN_2536; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2538 = 6'h2a == _T_392 ? _T_62 : _GEN_2537; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2539 = 6'h2b == _T_392 ? _T_63 : _GEN_2538; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2540 = 6'h2c == _T_392 ? _T_64 : _GEN_2539; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2541 = 6'h2d == _T_392 ? _T_65 : _GEN_2540; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2542 = 6'h2e == _T_392 ? _T_66 : _GEN_2541; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2543 = 6'h2f == _T_392 ? _T_67 : _GEN_2542; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2544 = 6'h30 == _T_392 ? _T_68 : _GEN_2543; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2545 = 6'h31 == _T_392 ? _T_69 : _GEN_2544; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2546 = 6'h32 == _T_392 ? _T_70 : _GEN_2545; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2547 = 6'h33 == _T_392 ? _T_71 : _GEN_2546; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2548 = 6'h34 == _T_392 ? _T_72 : _GEN_2547; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2549 = 6'h35 == _T_392 ? _T_73 : _GEN_2548; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2550 = 6'h36 == _T_392 ? _T_74 : _GEN_2549; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2551 = 6'h37 == _T_392 ? _T_75 : _GEN_2550; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2552 = 6'h38 == _T_392 ? _T_76 : _GEN_2551; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2553 = 6'h39 == _T_392 ? _T_77 : _GEN_2552; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2554 = 6'h3a == _T_392 ? _T_78 : _GEN_2553; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2555 = 6'h3b == _T_392 ? _T_79 : _GEN_2554; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2556 = 6'h3c == _T_392 ? _T_80 : _GEN_2555; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2557 = 6'h3d == _T_392 ? _T_81 : _GEN_2556; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2558 = 6'h3e == _T_392 ? _T_82 : _GEN_2557; // @[execute.scala 79:10:@1990.4]
  assign _GEN_2559 = 6'h3f == _T_392 ? _T_83 : _GEN_2558; // @[execute.scala 79:10:@1990.4]
  assign _T_394 = _T_384 ? _GEN_2495 : _GEN_2559; // @[execute.scala 79:10:@1990.4]
  assign _T_396 = io_amount < 6'h2c; // @[execute.scala 79:15:@1991.4]
  assign _T_398 = io_amount - 6'h2c; // @[execute.scala 79:37:@1992.4]
  assign _T_399 = $unsigned(_T_398); // @[execute.scala 79:37:@1993.4]
  assign _T_400 = _T_399[5:0]; // @[execute.scala 79:37:@1994.4]
  assign _T_403 = 6'h14 + io_amount; // @[execute.scala 79:60:@1995.4]
  assign _T_404 = 6'h14 + io_amount; // @[execute.scala 79:60:@1996.4]
  assign _GEN_2561 = 6'h1 == _T_400 ? _T_21 : _T_20; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2562 = 6'h2 == _T_400 ? _T_22 : _GEN_2561; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2563 = 6'h3 == _T_400 ? _T_23 : _GEN_2562; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2564 = 6'h4 == _T_400 ? _T_24 : _GEN_2563; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2565 = 6'h5 == _T_400 ? _T_25 : _GEN_2564; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2566 = 6'h6 == _T_400 ? _T_26 : _GEN_2565; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2567 = 6'h7 == _T_400 ? _T_27 : _GEN_2566; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2568 = 6'h8 == _T_400 ? _T_28 : _GEN_2567; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2569 = 6'h9 == _T_400 ? _T_29 : _GEN_2568; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2570 = 6'ha == _T_400 ? _T_30 : _GEN_2569; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2571 = 6'hb == _T_400 ? _T_31 : _GEN_2570; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2572 = 6'hc == _T_400 ? _T_32 : _GEN_2571; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2573 = 6'hd == _T_400 ? _T_33 : _GEN_2572; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2574 = 6'he == _T_400 ? _T_34 : _GEN_2573; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2575 = 6'hf == _T_400 ? _T_35 : _GEN_2574; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2576 = 6'h10 == _T_400 ? _T_36 : _GEN_2575; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2577 = 6'h11 == _T_400 ? _T_37 : _GEN_2576; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2578 = 6'h12 == _T_400 ? _T_38 : _GEN_2577; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2579 = 6'h13 == _T_400 ? _T_39 : _GEN_2578; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2580 = 6'h14 == _T_400 ? _T_40 : _GEN_2579; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2581 = 6'h15 == _T_400 ? _T_41 : _GEN_2580; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2582 = 6'h16 == _T_400 ? _T_42 : _GEN_2581; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2583 = 6'h17 == _T_400 ? _T_43 : _GEN_2582; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2584 = 6'h18 == _T_400 ? _T_44 : _GEN_2583; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2585 = 6'h19 == _T_400 ? _T_45 : _GEN_2584; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2586 = 6'h1a == _T_400 ? _T_46 : _GEN_2585; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2587 = 6'h1b == _T_400 ? _T_47 : _GEN_2586; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2588 = 6'h1c == _T_400 ? _T_48 : _GEN_2587; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2589 = 6'h1d == _T_400 ? _T_49 : _GEN_2588; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2590 = 6'h1e == _T_400 ? _T_50 : _GEN_2589; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2591 = 6'h1f == _T_400 ? _T_51 : _GEN_2590; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2592 = 6'h20 == _T_400 ? _T_52 : _GEN_2591; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2593 = 6'h21 == _T_400 ? _T_53 : _GEN_2592; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2594 = 6'h22 == _T_400 ? _T_54 : _GEN_2593; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2595 = 6'h23 == _T_400 ? _T_55 : _GEN_2594; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2596 = 6'h24 == _T_400 ? _T_56 : _GEN_2595; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2597 = 6'h25 == _T_400 ? _T_57 : _GEN_2596; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2598 = 6'h26 == _T_400 ? _T_58 : _GEN_2597; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2599 = 6'h27 == _T_400 ? _T_59 : _GEN_2598; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2600 = 6'h28 == _T_400 ? _T_60 : _GEN_2599; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2601 = 6'h29 == _T_400 ? _T_61 : _GEN_2600; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2602 = 6'h2a == _T_400 ? _T_62 : _GEN_2601; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2603 = 6'h2b == _T_400 ? _T_63 : _GEN_2602; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2604 = 6'h2c == _T_400 ? _T_64 : _GEN_2603; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2605 = 6'h2d == _T_400 ? _T_65 : _GEN_2604; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2606 = 6'h2e == _T_400 ? _T_66 : _GEN_2605; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2607 = 6'h2f == _T_400 ? _T_67 : _GEN_2606; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2608 = 6'h30 == _T_400 ? _T_68 : _GEN_2607; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2609 = 6'h31 == _T_400 ? _T_69 : _GEN_2608; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2610 = 6'h32 == _T_400 ? _T_70 : _GEN_2609; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2611 = 6'h33 == _T_400 ? _T_71 : _GEN_2610; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2612 = 6'h34 == _T_400 ? _T_72 : _GEN_2611; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2613 = 6'h35 == _T_400 ? _T_73 : _GEN_2612; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2614 = 6'h36 == _T_400 ? _T_74 : _GEN_2613; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2615 = 6'h37 == _T_400 ? _T_75 : _GEN_2614; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2616 = 6'h38 == _T_400 ? _T_76 : _GEN_2615; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2617 = 6'h39 == _T_400 ? _T_77 : _GEN_2616; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2618 = 6'h3a == _T_400 ? _T_78 : _GEN_2617; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2619 = 6'h3b == _T_400 ? _T_79 : _GEN_2618; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2620 = 6'h3c == _T_400 ? _T_80 : _GEN_2619; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2621 = 6'h3d == _T_400 ? _T_81 : _GEN_2620; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2622 = 6'h3e == _T_400 ? _T_82 : _GEN_2621; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2623 = 6'h3f == _T_400 ? _T_83 : _GEN_2622; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2625 = 6'h1 == _T_404 ? _T_21 : _T_20; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2626 = 6'h2 == _T_404 ? _T_22 : _GEN_2625; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2627 = 6'h3 == _T_404 ? _T_23 : _GEN_2626; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2628 = 6'h4 == _T_404 ? _T_24 : _GEN_2627; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2629 = 6'h5 == _T_404 ? _T_25 : _GEN_2628; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2630 = 6'h6 == _T_404 ? _T_26 : _GEN_2629; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2631 = 6'h7 == _T_404 ? _T_27 : _GEN_2630; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2632 = 6'h8 == _T_404 ? _T_28 : _GEN_2631; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2633 = 6'h9 == _T_404 ? _T_29 : _GEN_2632; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2634 = 6'ha == _T_404 ? _T_30 : _GEN_2633; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2635 = 6'hb == _T_404 ? _T_31 : _GEN_2634; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2636 = 6'hc == _T_404 ? _T_32 : _GEN_2635; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2637 = 6'hd == _T_404 ? _T_33 : _GEN_2636; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2638 = 6'he == _T_404 ? _T_34 : _GEN_2637; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2639 = 6'hf == _T_404 ? _T_35 : _GEN_2638; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2640 = 6'h10 == _T_404 ? _T_36 : _GEN_2639; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2641 = 6'h11 == _T_404 ? _T_37 : _GEN_2640; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2642 = 6'h12 == _T_404 ? _T_38 : _GEN_2641; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2643 = 6'h13 == _T_404 ? _T_39 : _GEN_2642; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2644 = 6'h14 == _T_404 ? _T_40 : _GEN_2643; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2645 = 6'h15 == _T_404 ? _T_41 : _GEN_2644; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2646 = 6'h16 == _T_404 ? _T_42 : _GEN_2645; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2647 = 6'h17 == _T_404 ? _T_43 : _GEN_2646; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2648 = 6'h18 == _T_404 ? _T_44 : _GEN_2647; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2649 = 6'h19 == _T_404 ? _T_45 : _GEN_2648; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2650 = 6'h1a == _T_404 ? _T_46 : _GEN_2649; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2651 = 6'h1b == _T_404 ? _T_47 : _GEN_2650; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2652 = 6'h1c == _T_404 ? _T_48 : _GEN_2651; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2653 = 6'h1d == _T_404 ? _T_49 : _GEN_2652; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2654 = 6'h1e == _T_404 ? _T_50 : _GEN_2653; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2655 = 6'h1f == _T_404 ? _T_51 : _GEN_2654; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2656 = 6'h20 == _T_404 ? _T_52 : _GEN_2655; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2657 = 6'h21 == _T_404 ? _T_53 : _GEN_2656; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2658 = 6'h22 == _T_404 ? _T_54 : _GEN_2657; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2659 = 6'h23 == _T_404 ? _T_55 : _GEN_2658; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2660 = 6'h24 == _T_404 ? _T_56 : _GEN_2659; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2661 = 6'h25 == _T_404 ? _T_57 : _GEN_2660; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2662 = 6'h26 == _T_404 ? _T_58 : _GEN_2661; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2663 = 6'h27 == _T_404 ? _T_59 : _GEN_2662; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2664 = 6'h28 == _T_404 ? _T_60 : _GEN_2663; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2665 = 6'h29 == _T_404 ? _T_61 : _GEN_2664; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2666 = 6'h2a == _T_404 ? _T_62 : _GEN_2665; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2667 = 6'h2b == _T_404 ? _T_63 : _GEN_2666; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2668 = 6'h2c == _T_404 ? _T_64 : _GEN_2667; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2669 = 6'h2d == _T_404 ? _T_65 : _GEN_2668; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2670 = 6'h2e == _T_404 ? _T_66 : _GEN_2669; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2671 = 6'h2f == _T_404 ? _T_67 : _GEN_2670; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2672 = 6'h30 == _T_404 ? _T_68 : _GEN_2671; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2673 = 6'h31 == _T_404 ? _T_69 : _GEN_2672; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2674 = 6'h32 == _T_404 ? _T_70 : _GEN_2673; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2675 = 6'h33 == _T_404 ? _T_71 : _GEN_2674; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2676 = 6'h34 == _T_404 ? _T_72 : _GEN_2675; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2677 = 6'h35 == _T_404 ? _T_73 : _GEN_2676; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2678 = 6'h36 == _T_404 ? _T_74 : _GEN_2677; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2679 = 6'h37 == _T_404 ? _T_75 : _GEN_2678; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2680 = 6'h38 == _T_404 ? _T_76 : _GEN_2679; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2681 = 6'h39 == _T_404 ? _T_77 : _GEN_2680; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2682 = 6'h3a == _T_404 ? _T_78 : _GEN_2681; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2683 = 6'h3b == _T_404 ? _T_79 : _GEN_2682; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2684 = 6'h3c == _T_404 ? _T_80 : _GEN_2683; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2685 = 6'h3d == _T_404 ? _T_81 : _GEN_2684; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2686 = 6'h3e == _T_404 ? _T_82 : _GEN_2685; // @[execute.scala 79:10:@1997.4]
  assign _GEN_2687 = 6'h3f == _T_404 ? _T_83 : _GEN_2686; // @[execute.scala 79:10:@1997.4]
  assign _T_406 = _T_396 ? _GEN_2623 : _GEN_2687; // @[execute.scala 79:10:@1997.4]
  assign _T_408 = io_amount < 6'h2b; // @[execute.scala 79:15:@1998.4]
  assign _T_410 = io_amount - 6'h2b; // @[execute.scala 79:37:@1999.4]
  assign _T_411 = $unsigned(_T_410); // @[execute.scala 79:37:@2000.4]
  assign _T_412 = _T_411[5:0]; // @[execute.scala 79:37:@2001.4]
  assign _T_415 = 6'h15 + io_amount; // @[execute.scala 79:60:@2002.4]
  assign _T_416 = 6'h15 + io_amount; // @[execute.scala 79:60:@2003.4]
  assign _GEN_2689 = 6'h1 == _T_412 ? _T_21 : _T_20; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2690 = 6'h2 == _T_412 ? _T_22 : _GEN_2689; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2691 = 6'h3 == _T_412 ? _T_23 : _GEN_2690; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2692 = 6'h4 == _T_412 ? _T_24 : _GEN_2691; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2693 = 6'h5 == _T_412 ? _T_25 : _GEN_2692; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2694 = 6'h6 == _T_412 ? _T_26 : _GEN_2693; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2695 = 6'h7 == _T_412 ? _T_27 : _GEN_2694; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2696 = 6'h8 == _T_412 ? _T_28 : _GEN_2695; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2697 = 6'h9 == _T_412 ? _T_29 : _GEN_2696; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2698 = 6'ha == _T_412 ? _T_30 : _GEN_2697; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2699 = 6'hb == _T_412 ? _T_31 : _GEN_2698; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2700 = 6'hc == _T_412 ? _T_32 : _GEN_2699; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2701 = 6'hd == _T_412 ? _T_33 : _GEN_2700; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2702 = 6'he == _T_412 ? _T_34 : _GEN_2701; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2703 = 6'hf == _T_412 ? _T_35 : _GEN_2702; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2704 = 6'h10 == _T_412 ? _T_36 : _GEN_2703; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2705 = 6'h11 == _T_412 ? _T_37 : _GEN_2704; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2706 = 6'h12 == _T_412 ? _T_38 : _GEN_2705; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2707 = 6'h13 == _T_412 ? _T_39 : _GEN_2706; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2708 = 6'h14 == _T_412 ? _T_40 : _GEN_2707; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2709 = 6'h15 == _T_412 ? _T_41 : _GEN_2708; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2710 = 6'h16 == _T_412 ? _T_42 : _GEN_2709; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2711 = 6'h17 == _T_412 ? _T_43 : _GEN_2710; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2712 = 6'h18 == _T_412 ? _T_44 : _GEN_2711; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2713 = 6'h19 == _T_412 ? _T_45 : _GEN_2712; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2714 = 6'h1a == _T_412 ? _T_46 : _GEN_2713; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2715 = 6'h1b == _T_412 ? _T_47 : _GEN_2714; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2716 = 6'h1c == _T_412 ? _T_48 : _GEN_2715; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2717 = 6'h1d == _T_412 ? _T_49 : _GEN_2716; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2718 = 6'h1e == _T_412 ? _T_50 : _GEN_2717; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2719 = 6'h1f == _T_412 ? _T_51 : _GEN_2718; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2720 = 6'h20 == _T_412 ? _T_52 : _GEN_2719; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2721 = 6'h21 == _T_412 ? _T_53 : _GEN_2720; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2722 = 6'h22 == _T_412 ? _T_54 : _GEN_2721; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2723 = 6'h23 == _T_412 ? _T_55 : _GEN_2722; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2724 = 6'h24 == _T_412 ? _T_56 : _GEN_2723; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2725 = 6'h25 == _T_412 ? _T_57 : _GEN_2724; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2726 = 6'h26 == _T_412 ? _T_58 : _GEN_2725; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2727 = 6'h27 == _T_412 ? _T_59 : _GEN_2726; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2728 = 6'h28 == _T_412 ? _T_60 : _GEN_2727; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2729 = 6'h29 == _T_412 ? _T_61 : _GEN_2728; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2730 = 6'h2a == _T_412 ? _T_62 : _GEN_2729; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2731 = 6'h2b == _T_412 ? _T_63 : _GEN_2730; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2732 = 6'h2c == _T_412 ? _T_64 : _GEN_2731; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2733 = 6'h2d == _T_412 ? _T_65 : _GEN_2732; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2734 = 6'h2e == _T_412 ? _T_66 : _GEN_2733; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2735 = 6'h2f == _T_412 ? _T_67 : _GEN_2734; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2736 = 6'h30 == _T_412 ? _T_68 : _GEN_2735; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2737 = 6'h31 == _T_412 ? _T_69 : _GEN_2736; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2738 = 6'h32 == _T_412 ? _T_70 : _GEN_2737; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2739 = 6'h33 == _T_412 ? _T_71 : _GEN_2738; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2740 = 6'h34 == _T_412 ? _T_72 : _GEN_2739; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2741 = 6'h35 == _T_412 ? _T_73 : _GEN_2740; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2742 = 6'h36 == _T_412 ? _T_74 : _GEN_2741; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2743 = 6'h37 == _T_412 ? _T_75 : _GEN_2742; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2744 = 6'h38 == _T_412 ? _T_76 : _GEN_2743; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2745 = 6'h39 == _T_412 ? _T_77 : _GEN_2744; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2746 = 6'h3a == _T_412 ? _T_78 : _GEN_2745; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2747 = 6'h3b == _T_412 ? _T_79 : _GEN_2746; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2748 = 6'h3c == _T_412 ? _T_80 : _GEN_2747; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2749 = 6'h3d == _T_412 ? _T_81 : _GEN_2748; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2750 = 6'h3e == _T_412 ? _T_82 : _GEN_2749; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2751 = 6'h3f == _T_412 ? _T_83 : _GEN_2750; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2753 = 6'h1 == _T_416 ? _T_21 : _T_20; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2754 = 6'h2 == _T_416 ? _T_22 : _GEN_2753; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2755 = 6'h3 == _T_416 ? _T_23 : _GEN_2754; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2756 = 6'h4 == _T_416 ? _T_24 : _GEN_2755; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2757 = 6'h5 == _T_416 ? _T_25 : _GEN_2756; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2758 = 6'h6 == _T_416 ? _T_26 : _GEN_2757; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2759 = 6'h7 == _T_416 ? _T_27 : _GEN_2758; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2760 = 6'h8 == _T_416 ? _T_28 : _GEN_2759; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2761 = 6'h9 == _T_416 ? _T_29 : _GEN_2760; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2762 = 6'ha == _T_416 ? _T_30 : _GEN_2761; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2763 = 6'hb == _T_416 ? _T_31 : _GEN_2762; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2764 = 6'hc == _T_416 ? _T_32 : _GEN_2763; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2765 = 6'hd == _T_416 ? _T_33 : _GEN_2764; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2766 = 6'he == _T_416 ? _T_34 : _GEN_2765; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2767 = 6'hf == _T_416 ? _T_35 : _GEN_2766; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2768 = 6'h10 == _T_416 ? _T_36 : _GEN_2767; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2769 = 6'h11 == _T_416 ? _T_37 : _GEN_2768; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2770 = 6'h12 == _T_416 ? _T_38 : _GEN_2769; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2771 = 6'h13 == _T_416 ? _T_39 : _GEN_2770; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2772 = 6'h14 == _T_416 ? _T_40 : _GEN_2771; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2773 = 6'h15 == _T_416 ? _T_41 : _GEN_2772; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2774 = 6'h16 == _T_416 ? _T_42 : _GEN_2773; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2775 = 6'h17 == _T_416 ? _T_43 : _GEN_2774; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2776 = 6'h18 == _T_416 ? _T_44 : _GEN_2775; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2777 = 6'h19 == _T_416 ? _T_45 : _GEN_2776; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2778 = 6'h1a == _T_416 ? _T_46 : _GEN_2777; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2779 = 6'h1b == _T_416 ? _T_47 : _GEN_2778; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2780 = 6'h1c == _T_416 ? _T_48 : _GEN_2779; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2781 = 6'h1d == _T_416 ? _T_49 : _GEN_2780; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2782 = 6'h1e == _T_416 ? _T_50 : _GEN_2781; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2783 = 6'h1f == _T_416 ? _T_51 : _GEN_2782; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2784 = 6'h20 == _T_416 ? _T_52 : _GEN_2783; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2785 = 6'h21 == _T_416 ? _T_53 : _GEN_2784; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2786 = 6'h22 == _T_416 ? _T_54 : _GEN_2785; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2787 = 6'h23 == _T_416 ? _T_55 : _GEN_2786; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2788 = 6'h24 == _T_416 ? _T_56 : _GEN_2787; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2789 = 6'h25 == _T_416 ? _T_57 : _GEN_2788; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2790 = 6'h26 == _T_416 ? _T_58 : _GEN_2789; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2791 = 6'h27 == _T_416 ? _T_59 : _GEN_2790; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2792 = 6'h28 == _T_416 ? _T_60 : _GEN_2791; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2793 = 6'h29 == _T_416 ? _T_61 : _GEN_2792; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2794 = 6'h2a == _T_416 ? _T_62 : _GEN_2793; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2795 = 6'h2b == _T_416 ? _T_63 : _GEN_2794; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2796 = 6'h2c == _T_416 ? _T_64 : _GEN_2795; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2797 = 6'h2d == _T_416 ? _T_65 : _GEN_2796; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2798 = 6'h2e == _T_416 ? _T_66 : _GEN_2797; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2799 = 6'h2f == _T_416 ? _T_67 : _GEN_2798; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2800 = 6'h30 == _T_416 ? _T_68 : _GEN_2799; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2801 = 6'h31 == _T_416 ? _T_69 : _GEN_2800; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2802 = 6'h32 == _T_416 ? _T_70 : _GEN_2801; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2803 = 6'h33 == _T_416 ? _T_71 : _GEN_2802; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2804 = 6'h34 == _T_416 ? _T_72 : _GEN_2803; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2805 = 6'h35 == _T_416 ? _T_73 : _GEN_2804; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2806 = 6'h36 == _T_416 ? _T_74 : _GEN_2805; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2807 = 6'h37 == _T_416 ? _T_75 : _GEN_2806; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2808 = 6'h38 == _T_416 ? _T_76 : _GEN_2807; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2809 = 6'h39 == _T_416 ? _T_77 : _GEN_2808; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2810 = 6'h3a == _T_416 ? _T_78 : _GEN_2809; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2811 = 6'h3b == _T_416 ? _T_79 : _GEN_2810; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2812 = 6'h3c == _T_416 ? _T_80 : _GEN_2811; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2813 = 6'h3d == _T_416 ? _T_81 : _GEN_2812; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2814 = 6'h3e == _T_416 ? _T_82 : _GEN_2813; // @[execute.scala 79:10:@2004.4]
  assign _GEN_2815 = 6'h3f == _T_416 ? _T_83 : _GEN_2814; // @[execute.scala 79:10:@2004.4]
  assign _T_418 = _T_408 ? _GEN_2751 : _GEN_2815; // @[execute.scala 79:10:@2004.4]
  assign _T_420 = io_amount < 6'h2a; // @[execute.scala 79:15:@2005.4]
  assign _T_422 = io_amount - 6'h2a; // @[execute.scala 79:37:@2006.4]
  assign _T_423 = $unsigned(_T_422); // @[execute.scala 79:37:@2007.4]
  assign _T_424 = _T_423[5:0]; // @[execute.scala 79:37:@2008.4]
  assign _T_427 = 6'h16 + io_amount; // @[execute.scala 79:60:@2009.4]
  assign _T_428 = 6'h16 + io_amount; // @[execute.scala 79:60:@2010.4]
  assign _GEN_2817 = 6'h1 == _T_424 ? _T_21 : _T_20; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2818 = 6'h2 == _T_424 ? _T_22 : _GEN_2817; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2819 = 6'h3 == _T_424 ? _T_23 : _GEN_2818; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2820 = 6'h4 == _T_424 ? _T_24 : _GEN_2819; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2821 = 6'h5 == _T_424 ? _T_25 : _GEN_2820; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2822 = 6'h6 == _T_424 ? _T_26 : _GEN_2821; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2823 = 6'h7 == _T_424 ? _T_27 : _GEN_2822; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2824 = 6'h8 == _T_424 ? _T_28 : _GEN_2823; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2825 = 6'h9 == _T_424 ? _T_29 : _GEN_2824; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2826 = 6'ha == _T_424 ? _T_30 : _GEN_2825; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2827 = 6'hb == _T_424 ? _T_31 : _GEN_2826; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2828 = 6'hc == _T_424 ? _T_32 : _GEN_2827; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2829 = 6'hd == _T_424 ? _T_33 : _GEN_2828; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2830 = 6'he == _T_424 ? _T_34 : _GEN_2829; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2831 = 6'hf == _T_424 ? _T_35 : _GEN_2830; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2832 = 6'h10 == _T_424 ? _T_36 : _GEN_2831; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2833 = 6'h11 == _T_424 ? _T_37 : _GEN_2832; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2834 = 6'h12 == _T_424 ? _T_38 : _GEN_2833; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2835 = 6'h13 == _T_424 ? _T_39 : _GEN_2834; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2836 = 6'h14 == _T_424 ? _T_40 : _GEN_2835; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2837 = 6'h15 == _T_424 ? _T_41 : _GEN_2836; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2838 = 6'h16 == _T_424 ? _T_42 : _GEN_2837; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2839 = 6'h17 == _T_424 ? _T_43 : _GEN_2838; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2840 = 6'h18 == _T_424 ? _T_44 : _GEN_2839; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2841 = 6'h19 == _T_424 ? _T_45 : _GEN_2840; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2842 = 6'h1a == _T_424 ? _T_46 : _GEN_2841; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2843 = 6'h1b == _T_424 ? _T_47 : _GEN_2842; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2844 = 6'h1c == _T_424 ? _T_48 : _GEN_2843; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2845 = 6'h1d == _T_424 ? _T_49 : _GEN_2844; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2846 = 6'h1e == _T_424 ? _T_50 : _GEN_2845; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2847 = 6'h1f == _T_424 ? _T_51 : _GEN_2846; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2848 = 6'h20 == _T_424 ? _T_52 : _GEN_2847; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2849 = 6'h21 == _T_424 ? _T_53 : _GEN_2848; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2850 = 6'h22 == _T_424 ? _T_54 : _GEN_2849; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2851 = 6'h23 == _T_424 ? _T_55 : _GEN_2850; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2852 = 6'h24 == _T_424 ? _T_56 : _GEN_2851; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2853 = 6'h25 == _T_424 ? _T_57 : _GEN_2852; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2854 = 6'h26 == _T_424 ? _T_58 : _GEN_2853; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2855 = 6'h27 == _T_424 ? _T_59 : _GEN_2854; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2856 = 6'h28 == _T_424 ? _T_60 : _GEN_2855; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2857 = 6'h29 == _T_424 ? _T_61 : _GEN_2856; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2858 = 6'h2a == _T_424 ? _T_62 : _GEN_2857; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2859 = 6'h2b == _T_424 ? _T_63 : _GEN_2858; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2860 = 6'h2c == _T_424 ? _T_64 : _GEN_2859; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2861 = 6'h2d == _T_424 ? _T_65 : _GEN_2860; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2862 = 6'h2e == _T_424 ? _T_66 : _GEN_2861; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2863 = 6'h2f == _T_424 ? _T_67 : _GEN_2862; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2864 = 6'h30 == _T_424 ? _T_68 : _GEN_2863; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2865 = 6'h31 == _T_424 ? _T_69 : _GEN_2864; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2866 = 6'h32 == _T_424 ? _T_70 : _GEN_2865; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2867 = 6'h33 == _T_424 ? _T_71 : _GEN_2866; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2868 = 6'h34 == _T_424 ? _T_72 : _GEN_2867; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2869 = 6'h35 == _T_424 ? _T_73 : _GEN_2868; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2870 = 6'h36 == _T_424 ? _T_74 : _GEN_2869; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2871 = 6'h37 == _T_424 ? _T_75 : _GEN_2870; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2872 = 6'h38 == _T_424 ? _T_76 : _GEN_2871; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2873 = 6'h39 == _T_424 ? _T_77 : _GEN_2872; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2874 = 6'h3a == _T_424 ? _T_78 : _GEN_2873; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2875 = 6'h3b == _T_424 ? _T_79 : _GEN_2874; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2876 = 6'h3c == _T_424 ? _T_80 : _GEN_2875; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2877 = 6'h3d == _T_424 ? _T_81 : _GEN_2876; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2878 = 6'h3e == _T_424 ? _T_82 : _GEN_2877; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2879 = 6'h3f == _T_424 ? _T_83 : _GEN_2878; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2881 = 6'h1 == _T_428 ? _T_21 : _T_20; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2882 = 6'h2 == _T_428 ? _T_22 : _GEN_2881; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2883 = 6'h3 == _T_428 ? _T_23 : _GEN_2882; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2884 = 6'h4 == _T_428 ? _T_24 : _GEN_2883; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2885 = 6'h5 == _T_428 ? _T_25 : _GEN_2884; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2886 = 6'h6 == _T_428 ? _T_26 : _GEN_2885; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2887 = 6'h7 == _T_428 ? _T_27 : _GEN_2886; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2888 = 6'h8 == _T_428 ? _T_28 : _GEN_2887; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2889 = 6'h9 == _T_428 ? _T_29 : _GEN_2888; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2890 = 6'ha == _T_428 ? _T_30 : _GEN_2889; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2891 = 6'hb == _T_428 ? _T_31 : _GEN_2890; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2892 = 6'hc == _T_428 ? _T_32 : _GEN_2891; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2893 = 6'hd == _T_428 ? _T_33 : _GEN_2892; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2894 = 6'he == _T_428 ? _T_34 : _GEN_2893; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2895 = 6'hf == _T_428 ? _T_35 : _GEN_2894; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2896 = 6'h10 == _T_428 ? _T_36 : _GEN_2895; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2897 = 6'h11 == _T_428 ? _T_37 : _GEN_2896; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2898 = 6'h12 == _T_428 ? _T_38 : _GEN_2897; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2899 = 6'h13 == _T_428 ? _T_39 : _GEN_2898; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2900 = 6'h14 == _T_428 ? _T_40 : _GEN_2899; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2901 = 6'h15 == _T_428 ? _T_41 : _GEN_2900; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2902 = 6'h16 == _T_428 ? _T_42 : _GEN_2901; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2903 = 6'h17 == _T_428 ? _T_43 : _GEN_2902; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2904 = 6'h18 == _T_428 ? _T_44 : _GEN_2903; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2905 = 6'h19 == _T_428 ? _T_45 : _GEN_2904; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2906 = 6'h1a == _T_428 ? _T_46 : _GEN_2905; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2907 = 6'h1b == _T_428 ? _T_47 : _GEN_2906; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2908 = 6'h1c == _T_428 ? _T_48 : _GEN_2907; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2909 = 6'h1d == _T_428 ? _T_49 : _GEN_2908; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2910 = 6'h1e == _T_428 ? _T_50 : _GEN_2909; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2911 = 6'h1f == _T_428 ? _T_51 : _GEN_2910; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2912 = 6'h20 == _T_428 ? _T_52 : _GEN_2911; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2913 = 6'h21 == _T_428 ? _T_53 : _GEN_2912; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2914 = 6'h22 == _T_428 ? _T_54 : _GEN_2913; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2915 = 6'h23 == _T_428 ? _T_55 : _GEN_2914; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2916 = 6'h24 == _T_428 ? _T_56 : _GEN_2915; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2917 = 6'h25 == _T_428 ? _T_57 : _GEN_2916; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2918 = 6'h26 == _T_428 ? _T_58 : _GEN_2917; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2919 = 6'h27 == _T_428 ? _T_59 : _GEN_2918; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2920 = 6'h28 == _T_428 ? _T_60 : _GEN_2919; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2921 = 6'h29 == _T_428 ? _T_61 : _GEN_2920; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2922 = 6'h2a == _T_428 ? _T_62 : _GEN_2921; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2923 = 6'h2b == _T_428 ? _T_63 : _GEN_2922; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2924 = 6'h2c == _T_428 ? _T_64 : _GEN_2923; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2925 = 6'h2d == _T_428 ? _T_65 : _GEN_2924; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2926 = 6'h2e == _T_428 ? _T_66 : _GEN_2925; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2927 = 6'h2f == _T_428 ? _T_67 : _GEN_2926; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2928 = 6'h30 == _T_428 ? _T_68 : _GEN_2927; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2929 = 6'h31 == _T_428 ? _T_69 : _GEN_2928; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2930 = 6'h32 == _T_428 ? _T_70 : _GEN_2929; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2931 = 6'h33 == _T_428 ? _T_71 : _GEN_2930; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2932 = 6'h34 == _T_428 ? _T_72 : _GEN_2931; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2933 = 6'h35 == _T_428 ? _T_73 : _GEN_2932; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2934 = 6'h36 == _T_428 ? _T_74 : _GEN_2933; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2935 = 6'h37 == _T_428 ? _T_75 : _GEN_2934; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2936 = 6'h38 == _T_428 ? _T_76 : _GEN_2935; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2937 = 6'h39 == _T_428 ? _T_77 : _GEN_2936; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2938 = 6'h3a == _T_428 ? _T_78 : _GEN_2937; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2939 = 6'h3b == _T_428 ? _T_79 : _GEN_2938; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2940 = 6'h3c == _T_428 ? _T_80 : _GEN_2939; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2941 = 6'h3d == _T_428 ? _T_81 : _GEN_2940; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2942 = 6'h3e == _T_428 ? _T_82 : _GEN_2941; // @[execute.scala 79:10:@2011.4]
  assign _GEN_2943 = 6'h3f == _T_428 ? _T_83 : _GEN_2942; // @[execute.scala 79:10:@2011.4]
  assign _T_430 = _T_420 ? _GEN_2879 : _GEN_2943; // @[execute.scala 79:10:@2011.4]
  assign _T_432 = io_amount < 6'h29; // @[execute.scala 79:15:@2012.4]
  assign _T_434 = io_amount - 6'h29; // @[execute.scala 79:37:@2013.4]
  assign _T_435 = $unsigned(_T_434); // @[execute.scala 79:37:@2014.4]
  assign _T_436 = _T_435[5:0]; // @[execute.scala 79:37:@2015.4]
  assign _T_439 = 6'h17 + io_amount; // @[execute.scala 79:60:@2016.4]
  assign _T_440 = 6'h17 + io_amount; // @[execute.scala 79:60:@2017.4]
  assign _GEN_2945 = 6'h1 == _T_436 ? _T_21 : _T_20; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2946 = 6'h2 == _T_436 ? _T_22 : _GEN_2945; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2947 = 6'h3 == _T_436 ? _T_23 : _GEN_2946; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2948 = 6'h4 == _T_436 ? _T_24 : _GEN_2947; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2949 = 6'h5 == _T_436 ? _T_25 : _GEN_2948; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2950 = 6'h6 == _T_436 ? _T_26 : _GEN_2949; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2951 = 6'h7 == _T_436 ? _T_27 : _GEN_2950; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2952 = 6'h8 == _T_436 ? _T_28 : _GEN_2951; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2953 = 6'h9 == _T_436 ? _T_29 : _GEN_2952; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2954 = 6'ha == _T_436 ? _T_30 : _GEN_2953; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2955 = 6'hb == _T_436 ? _T_31 : _GEN_2954; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2956 = 6'hc == _T_436 ? _T_32 : _GEN_2955; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2957 = 6'hd == _T_436 ? _T_33 : _GEN_2956; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2958 = 6'he == _T_436 ? _T_34 : _GEN_2957; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2959 = 6'hf == _T_436 ? _T_35 : _GEN_2958; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2960 = 6'h10 == _T_436 ? _T_36 : _GEN_2959; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2961 = 6'h11 == _T_436 ? _T_37 : _GEN_2960; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2962 = 6'h12 == _T_436 ? _T_38 : _GEN_2961; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2963 = 6'h13 == _T_436 ? _T_39 : _GEN_2962; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2964 = 6'h14 == _T_436 ? _T_40 : _GEN_2963; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2965 = 6'h15 == _T_436 ? _T_41 : _GEN_2964; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2966 = 6'h16 == _T_436 ? _T_42 : _GEN_2965; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2967 = 6'h17 == _T_436 ? _T_43 : _GEN_2966; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2968 = 6'h18 == _T_436 ? _T_44 : _GEN_2967; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2969 = 6'h19 == _T_436 ? _T_45 : _GEN_2968; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2970 = 6'h1a == _T_436 ? _T_46 : _GEN_2969; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2971 = 6'h1b == _T_436 ? _T_47 : _GEN_2970; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2972 = 6'h1c == _T_436 ? _T_48 : _GEN_2971; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2973 = 6'h1d == _T_436 ? _T_49 : _GEN_2972; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2974 = 6'h1e == _T_436 ? _T_50 : _GEN_2973; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2975 = 6'h1f == _T_436 ? _T_51 : _GEN_2974; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2976 = 6'h20 == _T_436 ? _T_52 : _GEN_2975; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2977 = 6'h21 == _T_436 ? _T_53 : _GEN_2976; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2978 = 6'h22 == _T_436 ? _T_54 : _GEN_2977; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2979 = 6'h23 == _T_436 ? _T_55 : _GEN_2978; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2980 = 6'h24 == _T_436 ? _T_56 : _GEN_2979; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2981 = 6'h25 == _T_436 ? _T_57 : _GEN_2980; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2982 = 6'h26 == _T_436 ? _T_58 : _GEN_2981; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2983 = 6'h27 == _T_436 ? _T_59 : _GEN_2982; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2984 = 6'h28 == _T_436 ? _T_60 : _GEN_2983; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2985 = 6'h29 == _T_436 ? _T_61 : _GEN_2984; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2986 = 6'h2a == _T_436 ? _T_62 : _GEN_2985; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2987 = 6'h2b == _T_436 ? _T_63 : _GEN_2986; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2988 = 6'h2c == _T_436 ? _T_64 : _GEN_2987; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2989 = 6'h2d == _T_436 ? _T_65 : _GEN_2988; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2990 = 6'h2e == _T_436 ? _T_66 : _GEN_2989; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2991 = 6'h2f == _T_436 ? _T_67 : _GEN_2990; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2992 = 6'h30 == _T_436 ? _T_68 : _GEN_2991; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2993 = 6'h31 == _T_436 ? _T_69 : _GEN_2992; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2994 = 6'h32 == _T_436 ? _T_70 : _GEN_2993; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2995 = 6'h33 == _T_436 ? _T_71 : _GEN_2994; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2996 = 6'h34 == _T_436 ? _T_72 : _GEN_2995; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2997 = 6'h35 == _T_436 ? _T_73 : _GEN_2996; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2998 = 6'h36 == _T_436 ? _T_74 : _GEN_2997; // @[execute.scala 79:10:@2018.4]
  assign _GEN_2999 = 6'h37 == _T_436 ? _T_75 : _GEN_2998; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3000 = 6'h38 == _T_436 ? _T_76 : _GEN_2999; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3001 = 6'h39 == _T_436 ? _T_77 : _GEN_3000; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3002 = 6'h3a == _T_436 ? _T_78 : _GEN_3001; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3003 = 6'h3b == _T_436 ? _T_79 : _GEN_3002; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3004 = 6'h3c == _T_436 ? _T_80 : _GEN_3003; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3005 = 6'h3d == _T_436 ? _T_81 : _GEN_3004; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3006 = 6'h3e == _T_436 ? _T_82 : _GEN_3005; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3007 = 6'h3f == _T_436 ? _T_83 : _GEN_3006; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3009 = 6'h1 == _T_440 ? _T_21 : _T_20; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3010 = 6'h2 == _T_440 ? _T_22 : _GEN_3009; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3011 = 6'h3 == _T_440 ? _T_23 : _GEN_3010; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3012 = 6'h4 == _T_440 ? _T_24 : _GEN_3011; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3013 = 6'h5 == _T_440 ? _T_25 : _GEN_3012; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3014 = 6'h6 == _T_440 ? _T_26 : _GEN_3013; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3015 = 6'h7 == _T_440 ? _T_27 : _GEN_3014; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3016 = 6'h8 == _T_440 ? _T_28 : _GEN_3015; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3017 = 6'h9 == _T_440 ? _T_29 : _GEN_3016; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3018 = 6'ha == _T_440 ? _T_30 : _GEN_3017; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3019 = 6'hb == _T_440 ? _T_31 : _GEN_3018; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3020 = 6'hc == _T_440 ? _T_32 : _GEN_3019; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3021 = 6'hd == _T_440 ? _T_33 : _GEN_3020; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3022 = 6'he == _T_440 ? _T_34 : _GEN_3021; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3023 = 6'hf == _T_440 ? _T_35 : _GEN_3022; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3024 = 6'h10 == _T_440 ? _T_36 : _GEN_3023; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3025 = 6'h11 == _T_440 ? _T_37 : _GEN_3024; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3026 = 6'h12 == _T_440 ? _T_38 : _GEN_3025; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3027 = 6'h13 == _T_440 ? _T_39 : _GEN_3026; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3028 = 6'h14 == _T_440 ? _T_40 : _GEN_3027; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3029 = 6'h15 == _T_440 ? _T_41 : _GEN_3028; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3030 = 6'h16 == _T_440 ? _T_42 : _GEN_3029; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3031 = 6'h17 == _T_440 ? _T_43 : _GEN_3030; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3032 = 6'h18 == _T_440 ? _T_44 : _GEN_3031; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3033 = 6'h19 == _T_440 ? _T_45 : _GEN_3032; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3034 = 6'h1a == _T_440 ? _T_46 : _GEN_3033; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3035 = 6'h1b == _T_440 ? _T_47 : _GEN_3034; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3036 = 6'h1c == _T_440 ? _T_48 : _GEN_3035; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3037 = 6'h1d == _T_440 ? _T_49 : _GEN_3036; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3038 = 6'h1e == _T_440 ? _T_50 : _GEN_3037; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3039 = 6'h1f == _T_440 ? _T_51 : _GEN_3038; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3040 = 6'h20 == _T_440 ? _T_52 : _GEN_3039; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3041 = 6'h21 == _T_440 ? _T_53 : _GEN_3040; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3042 = 6'h22 == _T_440 ? _T_54 : _GEN_3041; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3043 = 6'h23 == _T_440 ? _T_55 : _GEN_3042; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3044 = 6'h24 == _T_440 ? _T_56 : _GEN_3043; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3045 = 6'h25 == _T_440 ? _T_57 : _GEN_3044; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3046 = 6'h26 == _T_440 ? _T_58 : _GEN_3045; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3047 = 6'h27 == _T_440 ? _T_59 : _GEN_3046; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3048 = 6'h28 == _T_440 ? _T_60 : _GEN_3047; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3049 = 6'h29 == _T_440 ? _T_61 : _GEN_3048; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3050 = 6'h2a == _T_440 ? _T_62 : _GEN_3049; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3051 = 6'h2b == _T_440 ? _T_63 : _GEN_3050; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3052 = 6'h2c == _T_440 ? _T_64 : _GEN_3051; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3053 = 6'h2d == _T_440 ? _T_65 : _GEN_3052; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3054 = 6'h2e == _T_440 ? _T_66 : _GEN_3053; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3055 = 6'h2f == _T_440 ? _T_67 : _GEN_3054; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3056 = 6'h30 == _T_440 ? _T_68 : _GEN_3055; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3057 = 6'h31 == _T_440 ? _T_69 : _GEN_3056; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3058 = 6'h32 == _T_440 ? _T_70 : _GEN_3057; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3059 = 6'h33 == _T_440 ? _T_71 : _GEN_3058; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3060 = 6'h34 == _T_440 ? _T_72 : _GEN_3059; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3061 = 6'h35 == _T_440 ? _T_73 : _GEN_3060; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3062 = 6'h36 == _T_440 ? _T_74 : _GEN_3061; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3063 = 6'h37 == _T_440 ? _T_75 : _GEN_3062; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3064 = 6'h38 == _T_440 ? _T_76 : _GEN_3063; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3065 = 6'h39 == _T_440 ? _T_77 : _GEN_3064; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3066 = 6'h3a == _T_440 ? _T_78 : _GEN_3065; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3067 = 6'h3b == _T_440 ? _T_79 : _GEN_3066; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3068 = 6'h3c == _T_440 ? _T_80 : _GEN_3067; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3069 = 6'h3d == _T_440 ? _T_81 : _GEN_3068; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3070 = 6'h3e == _T_440 ? _T_82 : _GEN_3069; // @[execute.scala 79:10:@2018.4]
  assign _GEN_3071 = 6'h3f == _T_440 ? _T_83 : _GEN_3070; // @[execute.scala 79:10:@2018.4]
  assign _T_442 = _T_432 ? _GEN_3007 : _GEN_3071; // @[execute.scala 79:10:@2018.4]
  assign _T_444 = io_amount < 6'h28; // @[execute.scala 79:15:@2019.4]
  assign _T_446 = io_amount - 6'h28; // @[execute.scala 79:37:@2020.4]
  assign _T_447 = $unsigned(_T_446); // @[execute.scala 79:37:@2021.4]
  assign _T_448 = _T_447[5:0]; // @[execute.scala 79:37:@2022.4]
  assign _T_451 = 6'h18 + io_amount; // @[execute.scala 79:60:@2023.4]
  assign _T_452 = 6'h18 + io_amount; // @[execute.scala 79:60:@2024.4]
  assign _GEN_3073 = 6'h1 == _T_448 ? _T_21 : _T_20; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3074 = 6'h2 == _T_448 ? _T_22 : _GEN_3073; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3075 = 6'h3 == _T_448 ? _T_23 : _GEN_3074; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3076 = 6'h4 == _T_448 ? _T_24 : _GEN_3075; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3077 = 6'h5 == _T_448 ? _T_25 : _GEN_3076; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3078 = 6'h6 == _T_448 ? _T_26 : _GEN_3077; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3079 = 6'h7 == _T_448 ? _T_27 : _GEN_3078; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3080 = 6'h8 == _T_448 ? _T_28 : _GEN_3079; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3081 = 6'h9 == _T_448 ? _T_29 : _GEN_3080; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3082 = 6'ha == _T_448 ? _T_30 : _GEN_3081; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3083 = 6'hb == _T_448 ? _T_31 : _GEN_3082; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3084 = 6'hc == _T_448 ? _T_32 : _GEN_3083; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3085 = 6'hd == _T_448 ? _T_33 : _GEN_3084; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3086 = 6'he == _T_448 ? _T_34 : _GEN_3085; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3087 = 6'hf == _T_448 ? _T_35 : _GEN_3086; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3088 = 6'h10 == _T_448 ? _T_36 : _GEN_3087; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3089 = 6'h11 == _T_448 ? _T_37 : _GEN_3088; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3090 = 6'h12 == _T_448 ? _T_38 : _GEN_3089; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3091 = 6'h13 == _T_448 ? _T_39 : _GEN_3090; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3092 = 6'h14 == _T_448 ? _T_40 : _GEN_3091; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3093 = 6'h15 == _T_448 ? _T_41 : _GEN_3092; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3094 = 6'h16 == _T_448 ? _T_42 : _GEN_3093; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3095 = 6'h17 == _T_448 ? _T_43 : _GEN_3094; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3096 = 6'h18 == _T_448 ? _T_44 : _GEN_3095; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3097 = 6'h19 == _T_448 ? _T_45 : _GEN_3096; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3098 = 6'h1a == _T_448 ? _T_46 : _GEN_3097; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3099 = 6'h1b == _T_448 ? _T_47 : _GEN_3098; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3100 = 6'h1c == _T_448 ? _T_48 : _GEN_3099; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3101 = 6'h1d == _T_448 ? _T_49 : _GEN_3100; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3102 = 6'h1e == _T_448 ? _T_50 : _GEN_3101; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3103 = 6'h1f == _T_448 ? _T_51 : _GEN_3102; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3104 = 6'h20 == _T_448 ? _T_52 : _GEN_3103; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3105 = 6'h21 == _T_448 ? _T_53 : _GEN_3104; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3106 = 6'h22 == _T_448 ? _T_54 : _GEN_3105; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3107 = 6'h23 == _T_448 ? _T_55 : _GEN_3106; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3108 = 6'h24 == _T_448 ? _T_56 : _GEN_3107; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3109 = 6'h25 == _T_448 ? _T_57 : _GEN_3108; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3110 = 6'h26 == _T_448 ? _T_58 : _GEN_3109; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3111 = 6'h27 == _T_448 ? _T_59 : _GEN_3110; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3112 = 6'h28 == _T_448 ? _T_60 : _GEN_3111; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3113 = 6'h29 == _T_448 ? _T_61 : _GEN_3112; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3114 = 6'h2a == _T_448 ? _T_62 : _GEN_3113; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3115 = 6'h2b == _T_448 ? _T_63 : _GEN_3114; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3116 = 6'h2c == _T_448 ? _T_64 : _GEN_3115; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3117 = 6'h2d == _T_448 ? _T_65 : _GEN_3116; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3118 = 6'h2e == _T_448 ? _T_66 : _GEN_3117; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3119 = 6'h2f == _T_448 ? _T_67 : _GEN_3118; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3120 = 6'h30 == _T_448 ? _T_68 : _GEN_3119; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3121 = 6'h31 == _T_448 ? _T_69 : _GEN_3120; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3122 = 6'h32 == _T_448 ? _T_70 : _GEN_3121; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3123 = 6'h33 == _T_448 ? _T_71 : _GEN_3122; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3124 = 6'h34 == _T_448 ? _T_72 : _GEN_3123; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3125 = 6'h35 == _T_448 ? _T_73 : _GEN_3124; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3126 = 6'h36 == _T_448 ? _T_74 : _GEN_3125; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3127 = 6'h37 == _T_448 ? _T_75 : _GEN_3126; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3128 = 6'h38 == _T_448 ? _T_76 : _GEN_3127; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3129 = 6'h39 == _T_448 ? _T_77 : _GEN_3128; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3130 = 6'h3a == _T_448 ? _T_78 : _GEN_3129; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3131 = 6'h3b == _T_448 ? _T_79 : _GEN_3130; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3132 = 6'h3c == _T_448 ? _T_80 : _GEN_3131; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3133 = 6'h3d == _T_448 ? _T_81 : _GEN_3132; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3134 = 6'h3e == _T_448 ? _T_82 : _GEN_3133; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3135 = 6'h3f == _T_448 ? _T_83 : _GEN_3134; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3137 = 6'h1 == _T_452 ? _T_21 : _T_20; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3138 = 6'h2 == _T_452 ? _T_22 : _GEN_3137; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3139 = 6'h3 == _T_452 ? _T_23 : _GEN_3138; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3140 = 6'h4 == _T_452 ? _T_24 : _GEN_3139; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3141 = 6'h5 == _T_452 ? _T_25 : _GEN_3140; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3142 = 6'h6 == _T_452 ? _T_26 : _GEN_3141; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3143 = 6'h7 == _T_452 ? _T_27 : _GEN_3142; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3144 = 6'h8 == _T_452 ? _T_28 : _GEN_3143; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3145 = 6'h9 == _T_452 ? _T_29 : _GEN_3144; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3146 = 6'ha == _T_452 ? _T_30 : _GEN_3145; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3147 = 6'hb == _T_452 ? _T_31 : _GEN_3146; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3148 = 6'hc == _T_452 ? _T_32 : _GEN_3147; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3149 = 6'hd == _T_452 ? _T_33 : _GEN_3148; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3150 = 6'he == _T_452 ? _T_34 : _GEN_3149; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3151 = 6'hf == _T_452 ? _T_35 : _GEN_3150; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3152 = 6'h10 == _T_452 ? _T_36 : _GEN_3151; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3153 = 6'h11 == _T_452 ? _T_37 : _GEN_3152; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3154 = 6'h12 == _T_452 ? _T_38 : _GEN_3153; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3155 = 6'h13 == _T_452 ? _T_39 : _GEN_3154; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3156 = 6'h14 == _T_452 ? _T_40 : _GEN_3155; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3157 = 6'h15 == _T_452 ? _T_41 : _GEN_3156; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3158 = 6'h16 == _T_452 ? _T_42 : _GEN_3157; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3159 = 6'h17 == _T_452 ? _T_43 : _GEN_3158; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3160 = 6'h18 == _T_452 ? _T_44 : _GEN_3159; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3161 = 6'h19 == _T_452 ? _T_45 : _GEN_3160; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3162 = 6'h1a == _T_452 ? _T_46 : _GEN_3161; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3163 = 6'h1b == _T_452 ? _T_47 : _GEN_3162; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3164 = 6'h1c == _T_452 ? _T_48 : _GEN_3163; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3165 = 6'h1d == _T_452 ? _T_49 : _GEN_3164; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3166 = 6'h1e == _T_452 ? _T_50 : _GEN_3165; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3167 = 6'h1f == _T_452 ? _T_51 : _GEN_3166; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3168 = 6'h20 == _T_452 ? _T_52 : _GEN_3167; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3169 = 6'h21 == _T_452 ? _T_53 : _GEN_3168; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3170 = 6'h22 == _T_452 ? _T_54 : _GEN_3169; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3171 = 6'h23 == _T_452 ? _T_55 : _GEN_3170; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3172 = 6'h24 == _T_452 ? _T_56 : _GEN_3171; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3173 = 6'h25 == _T_452 ? _T_57 : _GEN_3172; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3174 = 6'h26 == _T_452 ? _T_58 : _GEN_3173; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3175 = 6'h27 == _T_452 ? _T_59 : _GEN_3174; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3176 = 6'h28 == _T_452 ? _T_60 : _GEN_3175; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3177 = 6'h29 == _T_452 ? _T_61 : _GEN_3176; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3178 = 6'h2a == _T_452 ? _T_62 : _GEN_3177; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3179 = 6'h2b == _T_452 ? _T_63 : _GEN_3178; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3180 = 6'h2c == _T_452 ? _T_64 : _GEN_3179; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3181 = 6'h2d == _T_452 ? _T_65 : _GEN_3180; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3182 = 6'h2e == _T_452 ? _T_66 : _GEN_3181; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3183 = 6'h2f == _T_452 ? _T_67 : _GEN_3182; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3184 = 6'h30 == _T_452 ? _T_68 : _GEN_3183; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3185 = 6'h31 == _T_452 ? _T_69 : _GEN_3184; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3186 = 6'h32 == _T_452 ? _T_70 : _GEN_3185; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3187 = 6'h33 == _T_452 ? _T_71 : _GEN_3186; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3188 = 6'h34 == _T_452 ? _T_72 : _GEN_3187; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3189 = 6'h35 == _T_452 ? _T_73 : _GEN_3188; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3190 = 6'h36 == _T_452 ? _T_74 : _GEN_3189; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3191 = 6'h37 == _T_452 ? _T_75 : _GEN_3190; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3192 = 6'h38 == _T_452 ? _T_76 : _GEN_3191; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3193 = 6'h39 == _T_452 ? _T_77 : _GEN_3192; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3194 = 6'h3a == _T_452 ? _T_78 : _GEN_3193; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3195 = 6'h3b == _T_452 ? _T_79 : _GEN_3194; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3196 = 6'h3c == _T_452 ? _T_80 : _GEN_3195; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3197 = 6'h3d == _T_452 ? _T_81 : _GEN_3196; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3198 = 6'h3e == _T_452 ? _T_82 : _GEN_3197; // @[execute.scala 79:10:@2025.4]
  assign _GEN_3199 = 6'h3f == _T_452 ? _T_83 : _GEN_3198; // @[execute.scala 79:10:@2025.4]
  assign _T_454 = _T_444 ? _GEN_3135 : _GEN_3199; // @[execute.scala 79:10:@2025.4]
  assign _T_456 = io_amount < 6'h27; // @[execute.scala 79:15:@2026.4]
  assign _T_458 = io_amount - 6'h27; // @[execute.scala 79:37:@2027.4]
  assign _T_459 = $unsigned(_T_458); // @[execute.scala 79:37:@2028.4]
  assign _T_460 = _T_459[5:0]; // @[execute.scala 79:37:@2029.4]
  assign _T_463 = 6'h19 + io_amount; // @[execute.scala 79:60:@2030.4]
  assign _T_464 = 6'h19 + io_amount; // @[execute.scala 79:60:@2031.4]
  assign _GEN_3201 = 6'h1 == _T_460 ? _T_21 : _T_20; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3202 = 6'h2 == _T_460 ? _T_22 : _GEN_3201; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3203 = 6'h3 == _T_460 ? _T_23 : _GEN_3202; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3204 = 6'h4 == _T_460 ? _T_24 : _GEN_3203; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3205 = 6'h5 == _T_460 ? _T_25 : _GEN_3204; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3206 = 6'h6 == _T_460 ? _T_26 : _GEN_3205; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3207 = 6'h7 == _T_460 ? _T_27 : _GEN_3206; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3208 = 6'h8 == _T_460 ? _T_28 : _GEN_3207; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3209 = 6'h9 == _T_460 ? _T_29 : _GEN_3208; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3210 = 6'ha == _T_460 ? _T_30 : _GEN_3209; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3211 = 6'hb == _T_460 ? _T_31 : _GEN_3210; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3212 = 6'hc == _T_460 ? _T_32 : _GEN_3211; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3213 = 6'hd == _T_460 ? _T_33 : _GEN_3212; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3214 = 6'he == _T_460 ? _T_34 : _GEN_3213; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3215 = 6'hf == _T_460 ? _T_35 : _GEN_3214; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3216 = 6'h10 == _T_460 ? _T_36 : _GEN_3215; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3217 = 6'h11 == _T_460 ? _T_37 : _GEN_3216; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3218 = 6'h12 == _T_460 ? _T_38 : _GEN_3217; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3219 = 6'h13 == _T_460 ? _T_39 : _GEN_3218; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3220 = 6'h14 == _T_460 ? _T_40 : _GEN_3219; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3221 = 6'h15 == _T_460 ? _T_41 : _GEN_3220; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3222 = 6'h16 == _T_460 ? _T_42 : _GEN_3221; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3223 = 6'h17 == _T_460 ? _T_43 : _GEN_3222; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3224 = 6'h18 == _T_460 ? _T_44 : _GEN_3223; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3225 = 6'h19 == _T_460 ? _T_45 : _GEN_3224; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3226 = 6'h1a == _T_460 ? _T_46 : _GEN_3225; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3227 = 6'h1b == _T_460 ? _T_47 : _GEN_3226; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3228 = 6'h1c == _T_460 ? _T_48 : _GEN_3227; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3229 = 6'h1d == _T_460 ? _T_49 : _GEN_3228; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3230 = 6'h1e == _T_460 ? _T_50 : _GEN_3229; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3231 = 6'h1f == _T_460 ? _T_51 : _GEN_3230; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3232 = 6'h20 == _T_460 ? _T_52 : _GEN_3231; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3233 = 6'h21 == _T_460 ? _T_53 : _GEN_3232; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3234 = 6'h22 == _T_460 ? _T_54 : _GEN_3233; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3235 = 6'h23 == _T_460 ? _T_55 : _GEN_3234; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3236 = 6'h24 == _T_460 ? _T_56 : _GEN_3235; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3237 = 6'h25 == _T_460 ? _T_57 : _GEN_3236; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3238 = 6'h26 == _T_460 ? _T_58 : _GEN_3237; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3239 = 6'h27 == _T_460 ? _T_59 : _GEN_3238; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3240 = 6'h28 == _T_460 ? _T_60 : _GEN_3239; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3241 = 6'h29 == _T_460 ? _T_61 : _GEN_3240; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3242 = 6'h2a == _T_460 ? _T_62 : _GEN_3241; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3243 = 6'h2b == _T_460 ? _T_63 : _GEN_3242; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3244 = 6'h2c == _T_460 ? _T_64 : _GEN_3243; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3245 = 6'h2d == _T_460 ? _T_65 : _GEN_3244; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3246 = 6'h2e == _T_460 ? _T_66 : _GEN_3245; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3247 = 6'h2f == _T_460 ? _T_67 : _GEN_3246; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3248 = 6'h30 == _T_460 ? _T_68 : _GEN_3247; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3249 = 6'h31 == _T_460 ? _T_69 : _GEN_3248; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3250 = 6'h32 == _T_460 ? _T_70 : _GEN_3249; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3251 = 6'h33 == _T_460 ? _T_71 : _GEN_3250; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3252 = 6'h34 == _T_460 ? _T_72 : _GEN_3251; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3253 = 6'h35 == _T_460 ? _T_73 : _GEN_3252; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3254 = 6'h36 == _T_460 ? _T_74 : _GEN_3253; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3255 = 6'h37 == _T_460 ? _T_75 : _GEN_3254; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3256 = 6'h38 == _T_460 ? _T_76 : _GEN_3255; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3257 = 6'h39 == _T_460 ? _T_77 : _GEN_3256; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3258 = 6'h3a == _T_460 ? _T_78 : _GEN_3257; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3259 = 6'h3b == _T_460 ? _T_79 : _GEN_3258; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3260 = 6'h3c == _T_460 ? _T_80 : _GEN_3259; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3261 = 6'h3d == _T_460 ? _T_81 : _GEN_3260; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3262 = 6'h3e == _T_460 ? _T_82 : _GEN_3261; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3263 = 6'h3f == _T_460 ? _T_83 : _GEN_3262; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3265 = 6'h1 == _T_464 ? _T_21 : _T_20; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3266 = 6'h2 == _T_464 ? _T_22 : _GEN_3265; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3267 = 6'h3 == _T_464 ? _T_23 : _GEN_3266; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3268 = 6'h4 == _T_464 ? _T_24 : _GEN_3267; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3269 = 6'h5 == _T_464 ? _T_25 : _GEN_3268; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3270 = 6'h6 == _T_464 ? _T_26 : _GEN_3269; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3271 = 6'h7 == _T_464 ? _T_27 : _GEN_3270; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3272 = 6'h8 == _T_464 ? _T_28 : _GEN_3271; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3273 = 6'h9 == _T_464 ? _T_29 : _GEN_3272; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3274 = 6'ha == _T_464 ? _T_30 : _GEN_3273; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3275 = 6'hb == _T_464 ? _T_31 : _GEN_3274; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3276 = 6'hc == _T_464 ? _T_32 : _GEN_3275; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3277 = 6'hd == _T_464 ? _T_33 : _GEN_3276; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3278 = 6'he == _T_464 ? _T_34 : _GEN_3277; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3279 = 6'hf == _T_464 ? _T_35 : _GEN_3278; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3280 = 6'h10 == _T_464 ? _T_36 : _GEN_3279; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3281 = 6'h11 == _T_464 ? _T_37 : _GEN_3280; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3282 = 6'h12 == _T_464 ? _T_38 : _GEN_3281; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3283 = 6'h13 == _T_464 ? _T_39 : _GEN_3282; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3284 = 6'h14 == _T_464 ? _T_40 : _GEN_3283; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3285 = 6'h15 == _T_464 ? _T_41 : _GEN_3284; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3286 = 6'h16 == _T_464 ? _T_42 : _GEN_3285; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3287 = 6'h17 == _T_464 ? _T_43 : _GEN_3286; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3288 = 6'h18 == _T_464 ? _T_44 : _GEN_3287; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3289 = 6'h19 == _T_464 ? _T_45 : _GEN_3288; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3290 = 6'h1a == _T_464 ? _T_46 : _GEN_3289; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3291 = 6'h1b == _T_464 ? _T_47 : _GEN_3290; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3292 = 6'h1c == _T_464 ? _T_48 : _GEN_3291; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3293 = 6'h1d == _T_464 ? _T_49 : _GEN_3292; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3294 = 6'h1e == _T_464 ? _T_50 : _GEN_3293; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3295 = 6'h1f == _T_464 ? _T_51 : _GEN_3294; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3296 = 6'h20 == _T_464 ? _T_52 : _GEN_3295; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3297 = 6'h21 == _T_464 ? _T_53 : _GEN_3296; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3298 = 6'h22 == _T_464 ? _T_54 : _GEN_3297; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3299 = 6'h23 == _T_464 ? _T_55 : _GEN_3298; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3300 = 6'h24 == _T_464 ? _T_56 : _GEN_3299; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3301 = 6'h25 == _T_464 ? _T_57 : _GEN_3300; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3302 = 6'h26 == _T_464 ? _T_58 : _GEN_3301; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3303 = 6'h27 == _T_464 ? _T_59 : _GEN_3302; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3304 = 6'h28 == _T_464 ? _T_60 : _GEN_3303; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3305 = 6'h29 == _T_464 ? _T_61 : _GEN_3304; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3306 = 6'h2a == _T_464 ? _T_62 : _GEN_3305; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3307 = 6'h2b == _T_464 ? _T_63 : _GEN_3306; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3308 = 6'h2c == _T_464 ? _T_64 : _GEN_3307; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3309 = 6'h2d == _T_464 ? _T_65 : _GEN_3308; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3310 = 6'h2e == _T_464 ? _T_66 : _GEN_3309; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3311 = 6'h2f == _T_464 ? _T_67 : _GEN_3310; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3312 = 6'h30 == _T_464 ? _T_68 : _GEN_3311; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3313 = 6'h31 == _T_464 ? _T_69 : _GEN_3312; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3314 = 6'h32 == _T_464 ? _T_70 : _GEN_3313; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3315 = 6'h33 == _T_464 ? _T_71 : _GEN_3314; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3316 = 6'h34 == _T_464 ? _T_72 : _GEN_3315; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3317 = 6'h35 == _T_464 ? _T_73 : _GEN_3316; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3318 = 6'h36 == _T_464 ? _T_74 : _GEN_3317; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3319 = 6'h37 == _T_464 ? _T_75 : _GEN_3318; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3320 = 6'h38 == _T_464 ? _T_76 : _GEN_3319; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3321 = 6'h39 == _T_464 ? _T_77 : _GEN_3320; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3322 = 6'h3a == _T_464 ? _T_78 : _GEN_3321; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3323 = 6'h3b == _T_464 ? _T_79 : _GEN_3322; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3324 = 6'h3c == _T_464 ? _T_80 : _GEN_3323; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3325 = 6'h3d == _T_464 ? _T_81 : _GEN_3324; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3326 = 6'h3e == _T_464 ? _T_82 : _GEN_3325; // @[execute.scala 79:10:@2032.4]
  assign _GEN_3327 = 6'h3f == _T_464 ? _T_83 : _GEN_3326; // @[execute.scala 79:10:@2032.4]
  assign _T_466 = _T_456 ? _GEN_3263 : _GEN_3327; // @[execute.scala 79:10:@2032.4]
  assign _T_468 = io_amount < 6'h26; // @[execute.scala 79:15:@2033.4]
  assign _T_470 = io_amount - 6'h26; // @[execute.scala 79:37:@2034.4]
  assign _T_471 = $unsigned(_T_470); // @[execute.scala 79:37:@2035.4]
  assign _T_472 = _T_471[5:0]; // @[execute.scala 79:37:@2036.4]
  assign _T_475 = 6'h1a + io_amount; // @[execute.scala 79:60:@2037.4]
  assign _T_476 = 6'h1a + io_amount; // @[execute.scala 79:60:@2038.4]
  assign _GEN_3329 = 6'h1 == _T_472 ? _T_21 : _T_20; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3330 = 6'h2 == _T_472 ? _T_22 : _GEN_3329; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3331 = 6'h3 == _T_472 ? _T_23 : _GEN_3330; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3332 = 6'h4 == _T_472 ? _T_24 : _GEN_3331; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3333 = 6'h5 == _T_472 ? _T_25 : _GEN_3332; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3334 = 6'h6 == _T_472 ? _T_26 : _GEN_3333; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3335 = 6'h7 == _T_472 ? _T_27 : _GEN_3334; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3336 = 6'h8 == _T_472 ? _T_28 : _GEN_3335; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3337 = 6'h9 == _T_472 ? _T_29 : _GEN_3336; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3338 = 6'ha == _T_472 ? _T_30 : _GEN_3337; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3339 = 6'hb == _T_472 ? _T_31 : _GEN_3338; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3340 = 6'hc == _T_472 ? _T_32 : _GEN_3339; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3341 = 6'hd == _T_472 ? _T_33 : _GEN_3340; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3342 = 6'he == _T_472 ? _T_34 : _GEN_3341; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3343 = 6'hf == _T_472 ? _T_35 : _GEN_3342; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3344 = 6'h10 == _T_472 ? _T_36 : _GEN_3343; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3345 = 6'h11 == _T_472 ? _T_37 : _GEN_3344; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3346 = 6'h12 == _T_472 ? _T_38 : _GEN_3345; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3347 = 6'h13 == _T_472 ? _T_39 : _GEN_3346; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3348 = 6'h14 == _T_472 ? _T_40 : _GEN_3347; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3349 = 6'h15 == _T_472 ? _T_41 : _GEN_3348; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3350 = 6'h16 == _T_472 ? _T_42 : _GEN_3349; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3351 = 6'h17 == _T_472 ? _T_43 : _GEN_3350; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3352 = 6'h18 == _T_472 ? _T_44 : _GEN_3351; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3353 = 6'h19 == _T_472 ? _T_45 : _GEN_3352; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3354 = 6'h1a == _T_472 ? _T_46 : _GEN_3353; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3355 = 6'h1b == _T_472 ? _T_47 : _GEN_3354; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3356 = 6'h1c == _T_472 ? _T_48 : _GEN_3355; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3357 = 6'h1d == _T_472 ? _T_49 : _GEN_3356; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3358 = 6'h1e == _T_472 ? _T_50 : _GEN_3357; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3359 = 6'h1f == _T_472 ? _T_51 : _GEN_3358; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3360 = 6'h20 == _T_472 ? _T_52 : _GEN_3359; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3361 = 6'h21 == _T_472 ? _T_53 : _GEN_3360; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3362 = 6'h22 == _T_472 ? _T_54 : _GEN_3361; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3363 = 6'h23 == _T_472 ? _T_55 : _GEN_3362; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3364 = 6'h24 == _T_472 ? _T_56 : _GEN_3363; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3365 = 6'h25 == _T_472 ? _T_57 : _GEN_3364; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3366 = 6'h26 == _T_472 ? _T_58 : _GEN_3365; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3367 = 6'h27 == _T_472 ? _T_59 : _GEN_3366; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3368 = 6'h28 == _T_472 ? _T_60 : _GEN_3367; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3369 = 6'h29 == _T_472 ? _T_61 : _GEN_3368; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3370 = 6'h2a == _T_472 ? _T_62 : _GEN_3369; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3371 = 6'h2b == _T_472 ? _T_63 : _GEN_3370; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3372 = 6'h2c == _T_472 ? _T_64 : _GEN_3371; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3373 = 6'h2d == _T_472 ? _T_65 : _GEN_3372; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3374 = 6'h2e == _T_472 ? _T_66 : _GEN_3373; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3375 = 6'h2f == _T_472 ? _T_67 : _GEN_3374; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3376 = 6'h30 == _T_472 ? _T_68 : _GEN_3375; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3377 = 6'h31 == _T_472 ? _T_69 : _GEN_3376; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3378 = 6'h32 == _T_472 ? _T_70 : _GEN_3377; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3379 = 6'h33 == _T_472 ? _T_71 : _GEN_3378; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3380 = 6'h34 == _T_472 ? _T_72 : _GEN_3379; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3381 = 6'h35 == _T_472 ? _T_73 : _GEN_3380; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3382 = 6'h36 == _T_472 ? _T_74 : _GEN_3381; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3383 = 6'h37 == _T_472 ? _T_75 : _GEN_3382; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3384 = 6'h38 == _T_472 ? _T_76 : _GEN_3383; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3385 = 6'h39 == _T_472 ? _T_77 : _GEN_3384; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3386 = 6'h3a == _T_472 ? _T_78 : _GEN_3385; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3387 = 6'h3b == _T_472 ? _T_79 : _GEN_3386; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3388 = 6'h3c == _T_472 ? _T_80 : _GEN_3387; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3389 = 6'h3d == _T_472 ? _T_81 : _GEN_3388; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3390 = 6'h3e == _T_472 ? _T_82 : _GEN_3389; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3391 = 6'h3f == _T_472 ? _T_83 : _GEN_3390; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3393 = 6'h1 == _T_476 ? _T_21 : _T_20; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3394 = 6'h2 == _T_476 ? _T_22 : _GEN_3393; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3395 = 6'h3 == _T_476 ? _T_23 : _GEN_3394; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3396 = 6'h4 == _T_476 ? _T_24 : _GEN_3395; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3397 = 6'h5 == _T_476 ? _T_25 : _GEN_3396; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3398 = 6'h6 == _T_476 ? _T_26 : _GEN_3397; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3399 = 6'h7 == _T_476 ? _T_27 : _GEN_3398; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3400 = 6'h8 == _T_476 ? _T_28 : _GEN_3399; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3401 = 6'h9 == _T_476 ? _T_29 : _GEN_3400; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3402 = 6'ha == _T_476 ? _T_30 : _GEN_3401; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3403 = 6'hb == _T_476 ? _T_31 : _GEN_3402; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3404 = 6'hc == _T_476 ? _T_32 : _GEN_3403; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3405 = 6'hd == _T_476 ? _T_33 : _GEN_3404; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3406 = 6'he == _T_476 ? _T_34 : _GEN_3405; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3407 = 6'hf == _T_476 ? _T_35 : _GEN_3406; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3408 = 6'h10 == _T_476 ? _T_36 : _GEN_3407; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3409 = 6'h11 == _T_476 ? _T_37 : _GEN_3408; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3410 = 6'h12 == _T_476 ? _T_38 : _GEN_3409; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3411 = 6'h13 == _T_476 ? _T_39 : _GEN_3410; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3412 = 6'h14 == _T_476 ? _T_40 : _GEN_3411; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3413 = 6'h15 == _T_476 ? _T_41 : _GEN_3412; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3414 = 6'h16 == _T_476 ? _T_42 : _GEN_3413; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3415 = 6'h17 == _T_476 ? _T_43 : _GEN_3414; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3416 = 6'h18 == _T_476 ? _T_44 : _GEN_3415; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3417 = 6'h19 == _T_476 ? _T_45 : _GEN_3416; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3418 = 6'h1a == _T_476 ? _T_46 : _GEN_3417; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3419 = 6'h1b == _T_476 ? _T_47 : _GEN_3418; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3420 = 6'h1c == _T_476 ? _T_48 : _GEN_3419; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3421 = 6'h1d == _T_476 ? _T_49 : _GEN_3420; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3422 = 6'h1e == _T_476 ? _T_50 : _GEN_3421; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3423 = 6'h1f == _T_476 ? _T_51 : _GEN_3422; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3424 = 6'h20 == _T_476 ? _T_52 : _GEN_3423; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3425 = 6'h21 == _T_476 ? _T_53 : _GEN_3424; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3426 = 6'h22 == _T_476 ? _T_54 : _GEN_3425; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3427 = 6'h23 == _T_476 ? _T_55 : _GEN_3426; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3428 = 6'h24 == _T_476 ? _T_56 : _GEN_3427; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3429 = 6'h25 == _T_476 ? _T_57 : _GEN_3428; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3430 = 6'h26 == _T_476 ? _T_58 : _GEN_3429; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3431 = 6'h27 == _T_476 ? _T_59 : _GEN_3430; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3432 = 6'h28 == _T_476 ? _T_60 : _GEN_3431; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3433 = 6'h29 == _T_476 ? _T_61 : _GEN_3432; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3434 = 6'h2a == _T_476 ? _T_62 : _GEN_3433; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3435 = 6'h2b == _T_476 ? _T_63 : _GEN_3434; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3436 = 6'h2c == _T_476 ? _T_64 : _GEN_3435; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3437 = 6'h2d == _T_476 ? _T_65 : _GEN_3436; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3438 = 6'h2e == _T_476 ? _T_66 : _GEN_3437; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3439 = 6'h2f == _T_476 ? _T_67 : _GEN_3438; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3440 = 6'h30 == _T_476 ? _T_68 : _GEN_3439; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3441 = 6'h31 == _T_476 ? _T_69 : _GEN_3440; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3442 = 6'h32 == _T_476 ? _T_70 : _GEN_3441; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3443 = 6'h33 == _T_476 ? _T_71 : _GEN_3442; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3444 = 6'h34 == _T_476 ? _T_72 : _GEN_3443; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3445 = 6'h35 == _T_476 ? _T_73 : _GEN_3444; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3446 = 6'h36 == _T_476 ? _T_74 : _GEN_3445; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3447 = 6'h37 == _T_476 ? _T_75 : _GEN_3446; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3448 = 6'h38 == _T_476 ? _T_76 : _GEN_3447; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3449 = 6'h39 == _T_476 ? _T_77 : _GEN_3448; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3450 = 6'h3a == _T_476 ? _T_78 : _GEN_3449; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3451 = 6'h3b == _T_476 ? _T_79 : _GEN_3450; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3452 = 6'h3c == _T_476 ? _T_80 : _GEN_3451; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3453 = 6'h3d == _T_476 ? _T_81 : _GEN_3452; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3454 = 6'h3e == _T_476 ? _T_82 : _GEN_3453; // @[execute.scala 79:10:@2039.4]
  assign _GEN_3455 = 6'h3f == _T_476 ? _T_83 : _GEN_3454; // @[execute.scala 79:10:@2039.4]
  assign _T_478 = _T_468 ? _GEN_3391 : _GEN_3455; // @[execute.scala 79:10:@2039.4]
  assign _T_480 = io_amount < 6'h25; // @[execute.scala 79:15:@2040.4]
  assign _T_482 = io_amount - 6'h25; // @[execute.scala 79:37:@2041.4]
  assign _T_483 = $unsigned(_T_482); // @[execute.scala 79:37:@2042.4]
  assign _T_484 = _T_483[5:0]; // @[execute.scala 79:37:@2043.4]
  assign _T_487 = 6'h1b + io_amount; // @[execute.scala 79:60:@2044.4]
  assign _T_488 = 6'h1b + io_amount; // @[execute.scala 79:60:@2045.4]
  assign _GEN_3457 = 6'h1 == _T_484 ? _T_21 : _T_20; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3458 = 6'h2 == _T_484 ? _T_22 : _GEN_3457; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3459 = 6'h3 == _T_484 ? _T_23 : _GEN_3458; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3460 = 6'h4 == _T_484 ? _T_24 : _GEN_3459; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3461 = 6'h5 == _T_484 ? _T_25 : _GEN_3460; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3462 = 6'h6 == _T_484 ? _T_26 : _GEN_3461; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3463 = 6'h7 == _T_484 ? _T_27 : _GEN_3462; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3464 = 6'h8 == _T_484 ? _T_28 : _GEN_3463; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3465 = 6'h9 == _T_484 ? _T_29 : _GEN_3464; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3466 = 6'ha == _T_484 ? _T_30 : _GEN_3465; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3467 = 6'hb == _T_484 ? _T_31 : _GEN_3466; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3468 = 6'hc == _T_484 ? _T_32 : _GEN_3467; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3469 = 6'hd == _T_484 ? _T_33 : _GEN_3468; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3470 = 6'he == _T_484 ? _T_34 : _GEN_3469; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3471 = 6'hf == _T_484 ? _T_35 : _GEN_3470; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3472 = 6'h10 == _T_484 ? _T_36 : _GEN_3471; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3473 = 6'h11 == _T_484 ? _T_37 : _GEN_3472; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3474 = 6'h12 == _T_484 ? _T_38 : _GEN_3473; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3475 = 6'h13 == _T_484 ? _T_39 : _GEN_3474; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3476 = 6'h14 == _T_484 ? _T_40 : _GEN_3475; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3477 = 6'h15 == _T_484 ? _T_41 : _GEN_3476; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3478 = 6'h16 == _T_484 ? _T_42 : _GEN_3477; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3479 = 6'h17 == _T_484 ? _T_43 : _GEN_3478; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3480 = 6'h18 == _T_484 ? _T_44 : _GEN_3479; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3481 = 6'h19 == _T_484 ? _T_45 : _GEN_3480; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3482 = 6'h1a == _T_484 ? _T_46 : _GEN_3481; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3483 = 6'h1b == _T_484 ? _T_47 : _GEN_3482; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3484 = 6'h1c == _T_484 ? _T_48 : _GEN_3483; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3485 = 6'h1d == _T_484 ? _T_49 : _GEN_3484; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3486 = 6'h1e == _T_484 ? _T_50 : _GEN_3485; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3487 = 6'h1f == _T_484 ? _T_51 : _GEN_3486; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3488 = 6'h20 == _T_484 ? _T_52 : _GEN_3487; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3489 = 6'h21 == _T_484 ? _T_53 : _GEN_3488; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3490 = 6'h22 == _T_484 ? _T_54 : _GEN_3489; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3491 = 6'h23 == _T_484 ? _T_55 : _GEN_3490; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3492 = 6'h24 == _T_484 ? _T_56 : _GEN_3491; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3493 = 6'h25 == _T_484 ? _T_57 : _GEN_3492; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3494 = 6'h26 == _T_484 ? _T_58 : _GEN_3493; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3495 = 6'h27 == _T_484 ? _T_59 : _GEN_3494; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3496 = 6'h28 == _T_484 ? _T_60 : _GEN_3495; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3497 = 6'h29 == _T_484 ? _T_61 : _GEN_3496; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3498 = 6'h2a == _T_484 ? _T_62 : _GEN_3497; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3499 = 6'h2b == _T_484 ? _T_63 : _GEN_3498; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3500 = 6'h2c == _T_484 ? _T_64 : _GEN_3499; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3501 = 6'h2d == _T_484 ? _T_65 : _GEN_3500; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3502 = 6'h2e == _T_484 ? _T_66 : _GEN_3501; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3503 = 6'h2f == _T_484 ? _T_67 : _GEN_3502; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3504 = 6'h30 == _T_484 ? _T_68 : _GEN_3503; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3505 = 6'h31 == _T_484 ? _T_69 : _GEN_3504; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3506 = 6'h32 == _T_484 ? _T_70 : _GEN_3505; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3507 = 6'h33 == _T_484 ? _T_71 : _GEN_3506; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3508 = 6'h34 == _T_484 ? _T_72 : _GEN_3507; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3509 = 6'h35 == _T_484 ? _T_73 : _GEN_3508; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3510 = 6'h36 == _T_484 ? _T_74 : _GEN_3509; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3511 = 6'h37 == _T_484 ? _T_75 : _GEN_3510; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3512 = 6'h38 == _T_484 ? _T_76 : _GEN_3511; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3513 = 6'h39 == _T_484 ? _T_77 : _GEN_3512; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3514 = 6'h3a == _T_484 ? _T_78 : _GEN_3513; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3515 = 6'h3b == _T_484 ? _T_79 : _GEN_3514; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3516 = 6'h3c == _T_484 ? _T_80 : _GEN_3515; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3517 = 6'h3d == _T_484 ? _T_81 : _GEN_3516; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3518 = 6'h3e == _T_484 ? _T_82 : _GEN_3517; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3519 = 6'h3f == _T_484 ? _T_83 : _GEN_3518; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3521 = 6'h1 == _T_488 ? _T_21 : _T_20; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3522 = 6'h2 == _T_488 ? _T_22 : _GEN_3521; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3523 = 6'h3 == _T_488 ? _T_23 : _GEN_3522; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3524 = 6'h4 == _T_488 ? _T_24 : _GEN_3523; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3525 = 6'h5 == _T_488 ? _T_25 : _GEN_3524; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3526 = 6'h6 == _T_488 ? _T_26 : _GEN_3525; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3527 = 6'h7 == _T_488 ? _T_27 : _GEN_3526; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3528 = 6'h8 == _T_488 ? _T_28 : _GEN_3527; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3529 = 6'h9 == _T_488 ? _T_29 : _GEN_3528; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3530 = 6'ha == _T_488 ? _T_30 : _GEN_3529; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3531 = 6'hb == _T_488 ? _T_31 : _GEN_3530; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3532 = 6'hc == _T_488 ? _T_32 : _GEN_3531; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3533 = 6'hd == _T_488 ? _T_33 : _GEN_3532; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3534 = 6'he == _T_488 ? _T_34 : _GEN_3533; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3535 = 6'hf == _T_488 ? _T_35 : _GEN_3534; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3536 = 6'h10 == _T_488 ? _T_36 : _GEN_3535; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3537 = 6'h11 == _T_488 ? _T_37 : _GEN_3536; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3538 = 6'h12 == _T_488 ? _T_38 : _GEN_3537; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3539 = 6'h13 == _T_488 ? _T_39 : _GEN_3538; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3540 = 6'h14 == _T_488 ? _T_40 : _GEN_3539; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3541 = 6'h15 == _T_488 ? _T_41 : _GEN_3540; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3542 = 6'h16 == _T_488 ? _T_42 : _GEN_3541; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3543 = 6'h17 == _T_488 ? _T_43 : _GEN_3542; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3544 = 6'h18 == _T_488 ? _T_44 : _GEN_3543; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3545 = 6'h19 == _T_488 ? _T_45 : _GEN_3544; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3546 = 6'h1a == _T_488 ? _T_46 : _GEN_3545; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3547 = 6'h1b == _T_488 ? _T_47 : _GEN_3546; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3548 = 6'h1c == _T_488 ? _T_48 : _GEN_3547; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3549 = 6'h1d == _T_488 ? _T_49 : _GEN_3548; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3550 = 6'h1e == _T_488 ? _T_50 : _GEN_3549; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3551 = 6'h1f == _T_488 ? _T_51 : _GEN_3550; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3552 = 6'h20 == _T_488 ? _T_52 : _GEN_3551; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3553 = 6'h21 == _T_488 ? _T_53 : _GEN_3552; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3554 = 6'h22 == _T_488 ? _T_54 : _GEN_3553; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3555 = 6'h23 == _T_488 ? _T_55 : _GEN_3554; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3556 = 6'h24 == _T_488 ? _T_56 : _GEN_3555; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3557 = 6'h25 == _T_488 ? _T_57 : _GEN_3556; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3558 = 6'h26 == _T_488 ? _T_58 : _GEN_3557; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3559 = 6'h27 == _T_488 ? _T_59 : _GEN_3558; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3560 = 6'h28 == _T_488 ? _T_60 : _GEN_3559; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3561 = 6'h29 == _T_488 ? _T_61 : _GEN_3560; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3562 = 6'h2a == _T_488 ? _T_62 : _GEN_3561; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3563 = 6'h2b == _T_488 ? _T_63 : _GEN_3562; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3564 = 6'h2c == _T_488 ? _T_64 : _GEN_3563; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3565 = 6'h2d == _T_488 ? _T_65 : _GEN_3564; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3566 = 6'h2e == _T_488 ? _T_66 : _GEN_3565; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3567 = 6'h2f == _T_488 ? _T_67 : _GEN_3566; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3568 = 6'h30 == _T_488 ? _T_68 : _GEN_3567; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3569 = 6'h31 == _T_488 ? _T_69 : _GEN_3568; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3570 = 6'h32 == _T_488 ? _T_70 : _GEN_3569; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3571 = 6'h33 == _T_488 ? _T_71 : _GEN_3570; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3572 = 6'h34 == _T_488 ? _T_72 : _GEN_3571; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3573 = 6'h35 == _T_488 ? _T_73 : _GEN_3572; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3574 = 6'h36 == _T_488 ? _T_74 : _GEN_3573; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3575 = 6'h37 == _T_488 ? _T_75 : _GEN_3574; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3576 = 6'h38 == _T_488 ? _T_76 : _GEN_3575; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3577 = 6'h39 == _T_488 ? _T_77 : _GEN_3576; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3578 = 6'h3a == _T_488 ? _T_78 : _GEN_3577; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3579 = 6'h3b == _T_488 ? _T_79 : _GEN_3578; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3580 = 6'h3c == _T_488 ? _T_80 : _GEN_3579; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3581 = 6'h3d == _T_488 ? _T_81 : _GEN_3580; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3582 = 6'h3e == _T_488 ? _T_82 : _GEN_3581; // @[execute.scala 79:10:@2046.4]
  assign _GEN_3583 = 6'h3f == _T_488 ? _T_83 : _GEN_3582; // @[execute.scala 79:10:@2046.4]
  assign _T_490 = _T_480 ? _GEN_3519 : _GEN_3583; // @[execute.scala 79:10:@2046.4]
  assign _T_492 = io_amount < 6'h24; // @[execute.scala 79:15:@2047.4]
  assign _T_494 = io_amount - 6'h24; // @[execute.scala 79:37:@2048.4]
  assign _T_495 = $unsigned(_T_494); // @[execute.scala 79:37:@2049.4]
  assign _T_496 = _T_495[5:0]; // @[execute.scala 79:37:@2050.4]
  assign _T_499 = 6'h1c + io_amount; // @[execute.scala 79:60:@2051.4]
  assign _T_500 = 6'h1c + io_amount; // @[execute.scala 79:60:@2052.4]
  assign _GEN_3585 = 6'h1 == _T_496 ? _T_21 : _T_20; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3586 = 6'h2 == _T_496 ? _T_22 : _GEN_3585; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3587 = 6'h3 == _T_496 ? _T_23 : _GEN_3586; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3588 = 6'h4 == _T_496 ? _T_24 : _GEN_3587; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3589 = 6'h5 == _T_496 ? _T_25 : _GEN_3588; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3590 = 6'h6 == _T_496 ? _T_26 : _GEN_3589; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3591 = 6'h7 == _T_496 ? _T_27 : _GEN_3590; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3592 = 6'h8 == _T_496 ? _T_28 : _GEN_3591; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3593 = 6'h9 == _T_496 ? _T_29 : _GEN_3592; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3594 = 6'ha == _T_496 ? _T_30 : _GEN_3593; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3595 = 6'hb == _T_496 ? _T_31 : _GEN_3594; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3596 = 6'hc == _T_496 ? _T_32 : _GEN_3595; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3597 = 6'hd == _T_496 ? _T_33 : _GEN_3596; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3598 = 6'he == _T_496 ? _T_34 : _GEN_3597; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3599 = 6'hf == _T_496 ? _T_35 : _GEN_3598; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3600 = 6'h10 == _T_496 ? _T_36 : _GEN_3599; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3601 = 6'h11 == _T_496 ? _T_37 : _GEN_3600; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3602 = 6'h12 == _T_496 ? _T_38 : _GEN_3601; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3603 = 6'h13 == _T_496 ? _T_39 : _GEN_3602; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3604 = 6'h14 == _T_496 ? _T_40 : _GEN_3603; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3605 = 6'h15 == _T_496 ? _T_41 : _GEN_3604; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3606 = 6'h16 == _T_496 ? _T_42 : _GEN_3605; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3607 = 6'h17 == _T_496 ? _T_43 : _GEN_3606; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3608 = 6'h18 == _T_496 ? _T_44 : _GEN_3607; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3609 = 6'h19 == _T_496 ? _T_45 : _GEN_3608; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3610 = 6'h1a == _T_496 ? _T_46 : _GEN_3609; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3611 = 6'h1b == _T_496 ? _T_47 : _GEN_3610; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3612 = 6'h1c == _T_496 ? _T_48 : _GEN_3611; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3613 = 6'h1d == _T_496 ? _T_49 : _GEN_3612; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3614 = 6'h1e == _T_496 ? _T_50 : _GEN_3613; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3615 = 6'h1f == _T_496 ? _T_51 : _GEN_3614; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3616 = 6'h20 == _T_496 ? _T_52 : _GEN_3615; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3617 = 6'h21 == _T_496 ? _T_53 : _GEN_3616; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3618 = 6'h22 == _T_496 ? _T_54 : _GEN_3617; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3619 = 6'h23 == _T_496 ? _T_55 : _GEN_3618; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3620 = 6'h24 == _T_496 ? _T_56 : _GEN_3619; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3621 = 6'h25 == _T_496 ? _T_57 : _GEN_3620; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3622 = 6'h26 == _T_496 ? _T_58 : _GEN_3621; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3623 = 6'h27 == _T_496 ? _T_59 : _GEN_3622; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3624 = 6'h28 == _T_496 ? _T_60 : _GEN_3623; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3625 = 6'h29 == _T_496 ? _T_61 : _GEN_3624; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3626 = 6'h2a == _T_496 ? _T_62 : _GEN_3625; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3627 = 6'h2b == _T_496 ? _T_63 : _GEN_3626; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3628 = 6'h2c == _T_496 ? _T_64 : _GEN_3627; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3629 = 6'h2d == _T_496 ? _T_65 : _GEN_3628; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3630 = 6'h2e == _T_496 ? _T_66 : _GEN_3629; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3631 = 6'h2f == _T_496 ? _T_67 : _GEN_3630; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3632 = 6'h30 == _T_496 ? _T_68 : _GEN_3631; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3633 = 6'h31 == _T_496 ? _T_69 : _GEN_3632; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3634 = 6'h32 == _T_496 ? _T_70 : _GEN_3633; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3635 = 6'h33 == _T_496 ? _T_71 : _GEN_3634; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3636 = 6'h34 == _T_496 ? _T_72 : _GEN_3635; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3637 = 6'h35 == _T_496 ? _T_73 : _GEN_3636; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3638 = 6'h36 == _T_496 ? _T_74 : _GEN_3637; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3639 = 6'h37 == _T_496 ? _T_75 : _GEN_3638; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3640 = 6'h38 == _T_496 ? _T_76 : _GEN_3639; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3641 = 6'h39 == _T_496 ? _T_77 : _GEN_3640; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3642 = 6'h3a == _T_496 ? _T_78 : _GEN_3641; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3643 = 6'h3b == _T_496 ? _T_79 : _GEN_3642; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3644 = 6'h3c == _T_496 ? _T_80 : _GEN_3643; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3645 = 6'h3d == _T_496 ? _T_81 : _GEN_3644; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3646 = 6'h3e == _T_496 ? _T_82 : _GEN_3645; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3647 = 6'h3f == _T_496 ? _T_83 : _GEN_3646; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3649 = 6'h1 == _T_500 ? _T_21 : _T_20; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3650 = 6'h2 == _T_500 ? _T_22 : _GEN_3649; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3651 = 6'h3 == _T_500 ? _T_23 : _GEN_3650; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3652 = 6'h4 == _T_500 ? _T_24 : _GEN_3651; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3653 = 6'h5 == _T_500 ? _T_25 : _GEN_3652; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3654 = 6'h6 == _T_500 ? _T_26 : _GEN_3653; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3655 = 6'h7 == _T_500 ? _T_27 : _GEN_3654; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3656 = 6'h8 == _T_500 ? _T_28 : _GEN_3655; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3657 = 6'h9 == _T_500 ? _T_29 : _GEN_3656; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3658 = 6'ha == _T_500 ? _T_30 : _GEN_3657; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3659 = 6'hb == _T_500 ? _T_31 : _GEN_3658; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3660 = 6'hc == _T_500 ? _T_32 : _GEN_3659; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3661 = 6'hd == _T_500 ? _T_33 : _GEN_3660; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3662 = 6'he == _T_500 ? _T_34 : _GEN_3661; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3663 = 6'hf == _T_500 ? _T_35 : _GEN_3662; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3664 = 6'h10 == _T_500 ? _T_36 : _GEN_3663; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3665 = 6'h11 == _T_500 ? _T_37 : _GEN_3664; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3666 = 6'h12 == _T_500 ? _T_38 : _GEN_3665; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3667 = 6'h13 == _T_500 ? _T_39 : _GEN_3666; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3668 = 6'h14 == _T_500 ? _T_40 : _GEN_3667; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3669 = 6'h15 == _T_500 ? _T_41 : _GEN_3668; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3670 = 6'h16 == _T_500 ? _T_42 : _GEN_3669; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3671 = 6'h17 == _T_500 ? _T_43 : _GEN_3670; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3672 = 6'h18 == _T_500 ? _T_44 : _GEN_3671; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3673 = 6'h19 == _T_500 ? _T_45 : _GEN_3672; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3674 = 6'h1a == _T_500 ? _T_46 : _GEN_3673; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3675 = 6'h1b == _T_500 ? _T_47 : _GEN_3674; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3676 = 6'h1c == _T_500 ? _T_48 : _GEN_3675; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3677 = 6'h1d == _T_500 ? _T_49 : _GEN_3676; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3678 = 6'h1e == _T_500 ? _T_50 : _GEN_3677; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3679 = 6'h1f == _T_500 ? _T_51 : _GEN_3678; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3680 = 6'h20 == _T_500 ? _T_52 : _GEN_3679; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3681 = 6'h21 == _T_500 ? _T_53 : _GEN_3680; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3682 = 6'h22 == _T_500 ? _T_54 : _GEN_3681; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3683 = 6'h23 == _T_500 ? _T_55 : _GEN_3682; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3684 = 6'h24 == _T_500 ? _T_56 : _GEN_3683; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3685 = 6'h25 == _T_500 ? _T_57 : _GEN_3684; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3686 = 6'h26 == _T_500 ? _T_58 : _GEN_3685; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3687 = 6'h27 == _T_500 ? _T_59 : _GEN_3686; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3688 = 6'h28 == _T_500 ? _T_60 : _GEN_3687; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3689 = 6'h29 == _T_500 ? _T_61 : _GEN_3688; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3690 = 6'h2a == _T_500 ? _T_62 : _GEN_3689; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3691 = 6'h2b == _T_500 ? _T_63 : _GEN_3690; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3692 = 6'h2c == _T_500 ? _T_64 : _GEN_3691; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3693 = 6'h2d == _T_500 ? _T_65 : _GEN_3692; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3694 = 6'h2e == _T_500 ? _T_66 : _GEN_3693; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3695 = 6'h2f == _T_500 ? _T_67 : _GEN_3694; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3696 = 6'h30 == _T_500 ? _T_68 : _GEN_3695; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3697 = 6'h31 == _T_500 ? _T_69 : _GEN_3696; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3698 = 6'h32 == _T_500 ? _T_70 : _GEN_3697; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3699 = 6'h33 == _T_500 ? _T_71 : _GEN_3698; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3700 = 6'h34 == _T_500 ? _T_72 : _GEN_3699; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3701 = 6'h35 == _T_500 ? _T_73 : _GEN_3700; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3702 = 6'h36 == _T_500 ? _T_74 : _GEN_3701; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3703 = 6'h37 == _T_500 ? _T_75 : _GEN_3702; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3704 = 6'h38 == _T_500 ? _T_76 : _GEN_3703; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3705 = 6'h39 == _T_500 ? _T_77 : _GEN_3704; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3706 = 6'h3a == _T_500 ? _T_78 : _GEN_3705; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3707 = 6'h3b == _T_500 ? _T_79 : _GEN_3706; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3708 = 6'h3c == _T_500 ? _T_80 : _GEN_3707; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3709 = 6'h3d == _T_500 ? _T_81 : _GEN_3708; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3710 = 6'h3e == _T_500 ? _T_82 : _GEN_3709; // @[execute.scala 79:10:@2053.4]
  assign _GEN_3711 = 6'h3f == _T_500 ? _T_83 : _GEN_3710; // @[execute.scala 79:10:@2053.4]
  assign _T_502 = _T_492 ? _GEN_3647 : _GEN_3711; // @[execute.scala 79:10:@2053.4]
  assign _T_504 = io_amount < 6'h23; // @[execute.scala 79:15:@2054.4]
  assign _T_506 = io_amount - 6'h23; // @[execute.scala 79:37:@2055.4]
  assign _T_507 = $unsigned(_T_506); // @[execute.scala 79:37:@2056.4]
  assign _T_508 = _T_507[5:0]; // @[execute.scala 79:37:@2057.4]
  assign _T_511 = 6'h1d + io_amount; // @[execute.scala 79:60:@2058.4]
  assign _T_512 = 6'h1d + io_amount; // @[execute.scala 79:60:@2059.4]
  assign _GEN_3713 = 6'h1 == _T_508 ? _T_21 : _T_20; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3714 = 6'h2 == _T_508 ? _T_22 : _GEN_3713; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3715 = 6'h3 == _T_508 ? _T_23 : _GEN_3714; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3716 = 6'h4 == _T_508 ? _T_24 : _GEN_3715; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3717 = 6'h5 == _T_508 ? _T_25 : _GEN_3716; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3718 = 6'h6 == _T_508 ? _T_26 : _GEN_3717; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3719 = 6'h7 == _T_508 ? _T_27 : _GEN_3718; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3720 = 6'h8 == _T_508 ? _T_28 : _GEN_3719; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3721 = 6'h9 == _T_508 ? _T_29 : _GEN_3720; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3722 = 6'ha == _T_508 ? _T_30 : _GEN_3721; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3723 = 6'hb == _T_508 ? _T_31 : _GEN_3722; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3724 = 6'hc == _T_508 ? _T_32 : _GEN_3723; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3725 = 6'hd == _T_508 ? _T_33 : _GEN_3724; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3726 = 6'he == _T_508 ? _T_34 : _GEN_3725; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3727 = 6'hf == _T_508 ? _T_35 : _GEN_3726; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3728 = 6'h10 == _T_508 ? _T_36 : _GEN_3727; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3729 = 6'h11 == _T_508 ? _T_37 : _GEN_3728; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3730 = 6'h12 == _T_508 ? _T_38 : _GEN_3729; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3731 = 6'h13 == _T_508 ? _T_39 : _GEN_3730; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3732 = 6'h14 == _T_508 ? _T_40 : _GEN_3731; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3733 = 6'h15 == _T_508 ? _T_41 : _GEN_3732; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3734 = 6'h16 == _T_508 ? _T_42 : _GEN_3733; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3735 = 6'h17 == _T_508 ? _T_43 : _GEN_3734; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3736 = 6'h18 == _T_508 ? _T_44 : _GEN_3735; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3737 = 6'h19 == _T_508 ? _T_45 : _GEN_3736; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3738 = 6'h1a == _T_508 ? _T_46 : _GEN_3737; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3739 = 6'h1b == _T_508 ? _T_47 : _GEN_3738; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3740 = 6'h1c == _T_508 ? _T_48 : _GEN_3739; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3741 = 6'h1d == _T_508 ? _T_49 : _GEN_3740; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3742 = 6'h1e == _T_508 ? _T_50 : _GEN_3741; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3743 = 6'h1f == _T_508 ? _T_51 : _GEN_3742; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3744 = 6'h20 == _T_508 ? _T_52 : _GEN_3743; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3745 = 6'h21 == _T_508 ? _T_53 : _GEN_3744; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3746 = 6'h22 == _T_508 ? _T_54 : _GEN_3745; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3747 = 6'h23 == _T_508 ? _T_55 : _GEN_3746; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3748 = 6'h24 == _T_508 ? _T_56 : _GEN_3747; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3749 = 6'h25 == _T_508 ? _T_57 : _GEN_3748; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3750 = 6'h26 == _T_508 ? _T_58 : _GEN_3749; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3751 = 6'h27 == _T_508 ? _T_59 : _GEN_3750; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3752 = 6'h28 == _T_508 ? _T_60 : _GEN_3751; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3753 = 6'h29 == _T_508 ? _T_61 : _GEN_3752; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3754 = 6'h2a == _T_508 ? _T_62 : _GEN_3753; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3755 = 6'h2b == _T_508 ? _T_63 : _GEN_3754; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3756 = 6'h2c == _T_508 ? _T_64 : _GEN_3755; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3757 = 6'h2d == _T_508 ? _T_65 : _GEN_3756; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3758 = 6'h2e == _T_508 ? _T_66 : _GEN_3757; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3759 = 6'h2f == _T_508 ? _T_67 : _GEN_3758; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3760 = 6'h30 == _T_508 ? _T_68 : _GEN_3759; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3761 = 6'h31 == _T_508 ? _T_69 : _GEN_3760; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3762 = 6'h32 == _T_508 ? _T_70 : _GEN_3761; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3763 = 6'h33 == _T_508 ? _T_71 : _GEN_3762; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3764 = 6'h34 == _T_508 ? _T_72 : _GEN_3763; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3765 = 6'h35 == _T_508 ? _T_73 : _GEN_3764; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3766 = 6'h36 == _T_508 ? _T_74 : _GEN_3765; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3767 = 6'h37 == _T_508 ? _T_75 : _GEN_3766; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3768 = 6'h38 == _T_508 ? _T_76 : _GEN_3767; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3769 = 6'h39 == _T_508 ? _T_77 : _GEN_3768; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3770 = 6'h3a == _T_508 ? _T_78 : _GEN_3769; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3771 = 6'h3b == _T_508 ? _T_79 : _GEN_3770; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3772 = 6'h3c == _T_508 ? _T_80 : _GEN_3771; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3773 = 6'h3d == _T_508 ? _T_81 : _GEN_3772; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3774 = 6'h3e == _T_508 ? _T_82 : _GEN_3773; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3775 = 6'h3f == _T_508 ? _T_83 : _GEN_3774; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3777 = 6'h1 == _T_512 ? _T_21 : _T_20; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3778 = 6'h2 == _T_512 ? _T_22 : _GEN_3777; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3779 = 6'h3 == _T_512 ? _T_23 : _GEN_3778; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3780 = 6'h4 == _T_512 ? _T_24 : _GEN_3779; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3781 = 6'h5 == _T_512 ? _T_25 : _GEN_3780; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3782 = 6'h6 == _T_512 ? _T_26 : _GEN_3781; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3783 = 6'h7 == _T_512 ? _T_27 : _GEN_3782; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3784 = 6'h8 == _T_512 ? _T_28 : _GEN_3783; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3785 = 6'h9 == _T_512 ? _T_29 : _GEN_3784; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3786 = 6'ha == _T_512 ? _T_30 : _GEN_3785; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3787 = 6'hb == _T_512 ? _T_31 : _GEN_3786; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3788 = 6'hc == _T_512 ? _T_32 : _GEN_3787; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3789 = 6'hd == _T_512 ? _T_33 : _GEN_3788; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3790 = 6'he == _T_512 ? _T_34 : _GEN_3789; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3791 = 6'hf == _T_512 ? _T_35 : _GEN_3790; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3792 = 6'h10 == _T_512 ? _T_36 : _GEN_3791; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3793 = 6'h11 == _T_512 ? _T_37 : _GEN_3792; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3794 = 6'h12 == _T_512 ? _T_38 : _GEN_3793; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3795 = 6'h13 == _T_512 ? _T_39 : _GEN_3794; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3796 = 6'h14 == _T_512 ? _T_40 : _GEN_3795; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3797 = 6'h15 == _T_512 ? _T_41 : _GEN_3796; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3798 = 6'h16 == _T_512 ? _T_42 : _GEN_3797; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3799 = 6'h17 == _T_512 ? _T_43 : _GEN_3798; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3800 = 6'h18 == _T_512 ? _T_44 : _GEN_3799; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3801 = 6'h19 == _T_512 ? _T_45 : _GEN_3800; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3802 = 6'h1a == _T_512 ? _T_46 : _GEN_3801; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3803 = 6'h1b == _T_512 ? _T_47 : _GEN_3802; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3804 = 6'h1c == _T_512 ? _T_48 : _GEN_3803; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3805 = 6'h1d == _T_512 ? _T_49 : _GEN_3804; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3806 = 6'h1e == _T_512 ? _T_50 : _GEN_3805; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3807 = 6'h1f == _T_512 ? _T_51 : _GEN_3806; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3808 = 6'h20 == _T_512 ? _T_52 : _GEN_3807; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3809 = 6'h21 == _T_512 ? _T_53 : _GEN_3808; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3810 = 6'h22 == _T_512 ? _T_54 : _GEN_3809; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3811 = 6'h23 == _T_512 ? _T_55 : _GEN_3810; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3812 = 6'h24 == _T_512 ? _T_56 : _GEN_3811; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3813 = 6'h25 == _T_512 ? _T_57 : _GEN_3812; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3814 = 6'h26 == _T_512 ? _T_58 : _GEN_3813; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3815 = 6'h27 == _T_512 ? _T_59 : _GEN_3814; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3816 = 6'h28 == _T_512 ? _T_60 : _GEN_3815; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3817 = 6'h29 == _T_512 ? _T_61 : _GEN_3816; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3818 = 6'h2a == _T_512 ? _T_62 : _GEN_3817; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3819 = 6'h2b == _T_512 ? _T_63 : _GEN_3818; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3820 = 6'h2c == _T_512 ? _T_64 : _GEN_3819; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3821 = 6'h2d == _T_512 ? _T_65 : _GEN_3820; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3822 = 6'h2e == _T_512 ? _T_66 : _GEN_3821; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3823 = 6'h2f == _T_512 ? _T_67 : _GEN_3822; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3824 = 6'h30 == _T_512 ? _T_68 : _GEN_3823; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3825 = 6'h31 == _T_512 ? _T_69 : _GEN_3824; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3826 = 6'h32 == _T_512 ? _T_70 : _GEN_3825; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3827 = 6'h33 == _T_512 ? _T_71 : _GEN_3826; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3828 = 6'h34 == _T_512 ? _T_72 : _GEN_3827; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3829 = 6'h35 == _T_512 ? _T_73 : _GEN_3828; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3830 = 6'h36 == _T_512 ? _T_74 : _GEN_3829; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3831 = 6'h37 == _T_512 ? _T_75 : _GEN_3830; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3832 = 6'h38 == _T_512 ? _T_76 : _GEN_3831; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3833 = 6'h39 == _T_512 ? _T_77 : _GEN_3832; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3834 = 6'h3a == _T_512 ? _T_78 : _GEN_3833; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3835 = 6'h3b == _T_512 ? _T_79 : _GEN_3834; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3836 = 6'h3c == _T_512 ? _T_80 : _GEN_3835; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3837 = 6'h3d == _T_512 ? _T_81 : _GEN_3836; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3838 = 6'h3e == _T_512 ? _T_82 : _GEN_3837; // @[execute.scala 79:10:@2060.4]
  assign _GEN_3839 = 6'h3f == _T_512 ? _T_83 : _GEN_3838; // @[execute.scala 79:10:@2060.4]
  assign _T_514 = _T_504 ? _GEN_3775 : _GEN_3839; // @[execute.scala 79:10:@2060.4]
  assign _T_516 = io_amount < 6'h22; // @[execute.scala 79:15:@2061.4]
  assign _T_518 = io_amount - 6'h22; // @[execute.scala 79:37:@2062.4]
  assign _T_519 = $unsigned(_T_518); // @[execute.scala 79:37:@2063.4]
  assign _T_520 = _T_519[5:0]; // @[execute.scala 79:37:@2064.4]
  assign _T_523 = 6'h1e + io_amount; // @[execute.scala 79:60:@2065.4]
  assign _T_524 = 6'h1e + io_amount; // @[execute.scala 79:60:@2066.4]
  assign _GEN_3841 = 6'h1 == _T_520 ? _T_21 : _T_20; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3842 = 6'h2 == _T_520 ? _T_22 : _GEN_3841; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3843 = 6'h3 == _T_520 ? _T_23 : _GEN_3842; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3844 = 6'h4 == _T_520 ? _T_24 : _GEN_3843; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3845 = 6'h5 == _T_520 ? _T_25 : _GEN_3844; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3846 = 6'h6 == _T_520 ? _T_26 : _GEN_3845; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3847 = 6'h7 == _T_520 ? _T_27 : _GEN_3846; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3848 = 6'h8 == _T_520 ? _T_28 : _GEN_3847; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3849 = 6'h9 == _T_520 ? _T_29 : _GEN_3848; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3850 = 6'ha == _T_520 ? _T_30 : _GEN_3849; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3851 = 6'hb == _T_520 ? _T_31 : _GEN_3850; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3852 = 6'hc == _T_520 ? _T_32 : _GEN_3851; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3853 = 6'hd == _T_520 ? _T_33 : _GEN_3852; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3854 = 6'he == _T_520 ? _T_34 : _GEN_3853; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3855 = 6'hf == _T_520 ? _T_35 : _GEN_3854; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3856 = 6'h10 == _T_520 ? _T_36 : _GEN_3855; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3857 = 6'h11 == _T_520 ? _T_37 : _GEN_3856; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3858 = 6'h12 == _T_520 ? _T_38 : _GEN_3857; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3859 = 6'h13 == _T_520 ? _T_39 : _GEN_3858; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3860 = 6'h14 == _T_520 ? _T_40 : _GEN_3859; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3861 = 6'h15 == _T_520 ? _T_41 : _GEN_3860; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3862 = 6'h16 == _T_520 ? _T_42 : _GEN_3861; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3863 = 6'h17 == _T_520 ? _T_43 : _GEN_3862; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3864 = 6'h18 == _T_520 ? _T_44 : _GEN_3863; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3865 = 6'h19 == _T_520 ? _T_45 : _GEN_3864; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3866 = 6'h1a == _T_520 ? _T_46 : _GEN_3865; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3867 = 6'h1b == _T_520 ? _T_47 : _GEN_3866; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3868 = 6'h1c == _T_520 ? _T_48 : _GEN_3867; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3869 = 6'h1d == _T_520 ? _T_49 : _GEN_3868; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3870 = 6'h1e == _T_520 ? _T_50 : _GEN_3869; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3871 = 6'h1f == _T_520 ? _T_51 : _GEN_3870; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3872 = 6'h20 == _T_520 ? _T_52 : _GEN_3871; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3873 = 6'h21 == _T_520 ? _T_53 : _GEN_3872; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3874 = 6'h22 == _T_520 ? _T_54 : _GEN_3873; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3875 = 6'h23 == _T_520 ? _T_55 : _GEN_3874; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3876 = 6'h24 == _T_520 ? _T_56 : _GEN_3875; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3877 = 6'h25 == _T_520 ? _T_57 : _GEN_3876; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3878 = 6'h26 == _T_520 ? _T_58 : _GEN_3877; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3879 = 6'h27 == _T_520 ? _T_59 : _GEN_3878; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3880 = 6'h28 == _T_520 ? _T_60 : _GEN_3879; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3881 = 6'h29 == _T_520 ? _T_61 : _GEN_3880; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3882 = 6'h2a == _T_520 ? _T_62 : _GEN_3881; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3883 = 6'h2b == _T_520 ? _T_63 : _GEN_3882; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3884 = 6'h2c == _T_520 ? _T_64 : _GEN_3883; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3885 = 6'h2d == _T_520 ? _T_65 : _GEN_3884; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3886 = 6'h2e == _T_520 ? _T_66 : _GEN_3885; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3887 = 6'h2f == _T_520 ? _T_67 : _GEN_3886; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3888 = 6'h30 == _T_520 ? _T_68 : _GEN_3887; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3889 = 6'h31 == _T_520 ? _T_69 : _GEN_3888; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3890 = 6'h32 == _T_520 ? _T_70 : _GEN_3889; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3891 = 6'h33 == _T_520 ? _T_71 : _GEN_3890; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3892 = 6'h34 == _T_520 ? _T_72 : _GEN_3891; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3893 = 6'h35 == _T_520 ? _T_73 : _GEN_3892; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3894 = 6'h36 == _T_520 ? _T_74 : _GEN_3893; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3895 = 6'h37 == _T_520 ? _T_75 : _GEN_3894; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3896 = 6'h38 == _T_520 ? _T_76 : _GEN_3895; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3897 = 6'h39 == _T_520 ? _T_77 : _GEN_3896; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3898 = 6'h3a == _T_520 ? _T_78 : _GEN_3897; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3899 = 6'h3b == _T_520 ? _T_79 : _GEN_3898; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3900 = 6'h3c == _T_520 ? _T_80 : _GEN_3899; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3901 = 6'h3d == _T_520 ? _T_81 : _GEN_3900; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3902 = 6'h3e == _T_520 ? _T_82 : _GEN_3901; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3903 = 6'h3f == _T_520 ? _T_83 : _GEN_3902; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3905 = 6'h1 == _T_524 ? _T_21 : _T_20; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3906 = 6'h2 == _T_524 ? _T_22 : _GEN_3905; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3907 = 6'h3 == _T_524 ? _T_23 : _GEN_3906; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3908 = 6'h4 == _T_524 ? _T_24 : _GEN_3907; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3909 = 6'h5 == _T_524 ? _T_25 : _GEN_3908; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3910 = 6'h6 == _T_524 ? _T_26 : _GEN_3909; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3911 = 6'h7 == _T_524 ? _T_27 : _GEN_3910; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3912 = 6'h8 == _T_524 ? _T_28 : _GEN_3911; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3913 = 6'h9 == _T_524 ? _T_29 : _GEN_3912; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3914 = 6'ha == _T_524 ? _T_30 : _GEN_3913; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3915 = 6'hb == _T_524 ? _T_31 : _GEN_3914; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3916 = 6'hc == _T_524 ? _T_32 : _GEN_3915; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3917 = 6'hd == _T_524 ? _T_33 : _GEN_3916; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3918 = 6'he == _T_524 ? _T_34 : _GEN_3917; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3919 = 6'hf == _T_524 ? _T_35 : _GEN_3918; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3920 = 6'h10 == _T_524 ? _T_36 : _GEN_3919; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3921 = 6'h11 == _T_524 ? _T_37 : _GEN_3920; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3922 = 6'h12 == _T_524 ? _T_38 : _GEN_3921; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3923 = 6'h13 == _T_524 ? _T_39 : _GEN_3922; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3924 = 6'h14 == _T_524 ? _T_40 : _GEN_3923; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3925 = 6'h15 == _T_524 ? _T_41 : _GEN_3924; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3926 = 6'h16 == _T_524 ? _T_42 : _GEN_3925; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3927 = 6'h17 == _T_524 ? _T_43 : _GEN_3926; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3928 = 6'h18 == _T_524 ? _T_44 : _GEN_3927; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3929 = 6'h19 == _T_524 ? _T_45 : _GEN_3928; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3930 = 6'h1a == _T_524 ? _T_46 : _GEN_3929; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3931 = 6'h1b == _T_524 ? _T_47 : _GEN_3930; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3932 = 6'h1c == _T_524 ? _T_48 : _GEN_3931; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3933 = 6'h1d == _T_524 ? _T_49 : _GEN_3932; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3934 = 6'h1e == _T_524 ? _T_50 : _GEN_3933; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3935 = 6'h1f == _T_524 ? _T_51 : _GEN_3934; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3936 = 6'h20 == _T_524 ? _T_52 : _GEN_3935; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3937 = 6'h21 == _T_524 ? _T_53 : _GEN_3936; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3938 = 6'h22 == _T_524 ? _T_54 : _GEN_3937; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3939 = 6'h23 == _T_524 ? _T_55 : _GEN_3938; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3940 = 6'h24 == _T_524 ? _T_56 : _GEN_3939; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3941 = 6'h25 == _T_524 ? _T_57 : _GEN_3940; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3942 = 6'h26 == _T_524 ? _T_58 : _GEN_3941; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3943 = 6'h27 == _T_524 ? _T_59 : _GEN_3942; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3944 = 6'h28 == _T_524 ? _T_60 : _GEN_3943; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3945 = 6'h29 == _T_524 ? _T_61 : _GEN_3944; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3946 = 6'h2a == _T_524 ? _T_62 : _GEN_3945; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3947 = 6'h2b == _T_524 ? _T_63 : _GEN_3946; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3948 = 6'h2c == _T_524 ? _T_64 : _GEN_3947; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3949 = 6'h2d == _T_524 ? _T_65 : _GEN_3948; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3950 = 6'h2e == _T_524 ? _T_66 : _GEN_3949; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3951 = 6'h2f == _T_524 ? _T_67 : _GEN_3950; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3952 = 6'h30 == _T_524 ? _T_68 : _GEN_3951; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3953 = 6'h31 == _T_524 ? _T_69 : _GEN_3952; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3954 = 6'h32 == _T_524 ? _T_70 : _GEN_3953; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3955 = 6'h33 == _T_524 ? _T_71 : _GEN_3954; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3956 = 6'h34 == _T_524 ? _T_72 : _GEN_3955; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3957 = 6'h35 == _T_524 ? _T_73 : _GEN_3956; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3958 = 6'h36 == _T_524 ? _T_74 : _GEN_3957; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3959 = 6'h37 == _T_524 ? _T_75 : _GEN_3958; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3960 = 6'h38 == _T_524 ? _T_76 : _GEN_3959; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3961 = 6'h39 == _T_524 ? _T_77 : _GEN_3960; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3962 = 6'h3a == _T_524 ? _T_78 : _GEN_3961; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3963 = 6'h3b == _T_524 ? _T_79 : _GEN_3962; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3964 = 6'h3c == _T_524 ? _T_80 : _GEN_3963; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3965 = 6'h3d == _T_524 ? _T_81 : _GEN_3964; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3966 = 6'h3e == _T_524 ? _T_82 : _GEN_3965; // @[execute.scala 79:10:@2067.4]
  assign _GEN_3967 = 6'h3f == _T_524 ? _T_83 : _GEN_3966; // @[execute.scala 79:10:@2067.4]
  assign _T_526 = _T_516 ? _GEN_3903 : _GEN_3967; // @[execute.scala 79:10:@2067.4]
  assign _T_528 = io_amount < 6'h21; // @[execute.scala 79:15:@2068.4]
  assign _T_530 = io_amount - 6'h21; // @[execute.scala 79:37:@2069.4]
  assign _T_531 = $unsigned(_T_530); // @[execute.scala 79:37:@2070.4]
  assign _T_532 = _T_531[5:0]; // @[execute.scala 79:37:@2071.4]
  assign _T_535 = 6'h1f + io_amount; // @[execute.scala 79:60:@2072.4]
  assign _T_536 = 6'h1f + io_amount; // @[execute.scala 79:60:@2073.4]
  assign _GEN_3969 = 6'h1 == _T_532 ? _T_21 : _T_20; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3970 = 6'h2 == _T_532 ? _T_22 : _GEN_3969; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3971 = 6'h3 == _T_532 ? _T_23 : _GEN_3970; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3972 = 6'h4 == _T_532 ? _T_24 : _GEN_3971; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3973 = 6'h5 == _T_532 ? _T_25 : _GEN_3972; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3974 = 6'h6 == _T_532 ? _T_26 : _GEN_3973; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3975 = 6'h7 == _T_532 ? _T_27 : _GEN_3974; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3976 = 6'h8 == _T_532 ? _T_28 : _GEN_3975; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3977 = 6'h9 == _T_532 ? _T_29 : _GEN_3976; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3978 = 6'ha == _T_532 ? _T_30 : _GEN_3977; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3979 = 6'hb == _T_532 ? _T_31 : _GEN_3978; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3980 = 6'hc == _T_532 ? _T_32 : _GEN_3979; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3981 = 6'hd == _T_532 ? _T_33 : _GEN_3980; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3982 = 6'he == _T_532 ? _T_34 : _GEN_3981; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3983 = 6'hf == _T_532 ? _T_35 : _GEN_3982; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3984 = 6'h10 == _T_532 ? _T_36 : _GEN_3983; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3985 = 6'h11 == _T_532 ? _T_37 : _GEN_3984; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3986 = 6'h12 == _T_532 ? _T_38 : _GEN_3985; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3987 = 6'h13 == _T_532 ? _T_39 : _GEN_3986; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3988 = 6'h14 == _T_532 ? _T_40 : _GEN_3987; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3989 = 6'h15 == _T_532 ? _T_41 : _GEN_3988; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3990 = 6'h16 == _T_532 ? _T_42 : _GEN_3989; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3991 = 6'h17 == _T_532 ? _T_43 : _GEN_3990; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3992 = 6'h18 == _T_532 ? _T_44 : _GEN_3991; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3993 = 6'h19 == _T_532 ? _T_45 : _GEN_3992; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3994 = 6'h1a == _T_532 ? _T_46 : _GEN_3993; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3995 = 6'h1b == _T_532 ? _T_47 : _GEN_3994; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3996 = 6'h1c == _T_532 ? _T_48 : _GEN_3995; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3997 = 6'h1d == _T_532 ? _T_49 : _GEN_3996; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3998 = 6'h1e == _T_532 ? _T_50 : _GEN_3997; // @[execute.scala 79:10:@2074.4]
  assign _GEN_3999 = 6'h1f == _T_532 ? _T_51 : _GEN_3998; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4000 = 6'h20 == _T_532 ? _T_52 : _GEN_3999; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4001 = 6'h21 == _T_532 ? _T_53 : _GEN_4000; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4002 = 6'h22 == _T_532 ? _T_54 : _GEN_4001; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4003 = 6'h23 == _T_532 ? _T_55 : _GEN_4002; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4004 = 6'h24 == _T_532 ? _T_56 : _GEN_4003; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4005 = 6'h25 == _T_532 ? _T_57 : _GEN_4004; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4006 = 6'h26 == _T_532 ? _T_58 : _GEN_4005; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4007 = 6'h27 == _T_532 ? _T_59 : _GEN_4006; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4008 = 6'h28 == _T_532 ? _T_60 : _GEN_4007; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4009 = 6'h29 == _T_532 ? _T_61 : _GEN_4008; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4010 = 6'h2a == _T_532 ? _T_62 : _GEN_4009; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4011 = 6'h2b == _T_532 ? _T_63 : _GEN_4010; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4012 = 6'h2c == _T_532 ? _T_64 : _GEN_4011; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4013 = 6'h2d == _T_532 ? _T_65 : _GEN_4012; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4014 = 6'h2e == _T_532 ? _T_66 : _GEN_4013; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4015 = 6'h2f == _T_532 ? _T_67 : _GEN_4014; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4016 = 6'h30 == _T_532 ? _T_68 : _GEN_4015; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4017 = 6'h31 == _T_532 ? _T_69 : _GEN_4016; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4018 = 6'h32 == _T_532 ? _T_70 : _GEN_4017; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4019 = 6'h33 == _T_532 ? _T_71 : _GEN_4018; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4020 = 6'h34 == _T_532 ? _T_72 : _GEN_4019; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4021 = 6'h35 == _T_532 ? _T_73 : _GEN_4020; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4022 = 6'h36 == _T_532 ? _T_74 : _GEN_4021; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4023 = 6'h37 == _T_532 ? _T_75 : _GEN_4022; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4024 = 6'h38 == _T_532 ? _T_76 : _GEN_4023; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4025 = 6'h39 == _T_532 ? _T_77 : _GEN_4024; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4026 = 6'h3a == _T_532 ? _T_78 : _GEN_4025; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4027 = 6'h3b == _T_532 ? _T_79 : _GEN_4026; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4028 = 6'h3c == _T_532 ? _T_80 : _GEN_4027; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4029 = 6'h3d == _T_532 ? _T_81 : _GEN_4028; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4030 = 6'h3e == _T_532 ? _T_82 : _GEN_4029; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4031 = 6'h3f == _T_532 ? _T_83 : _GEN_4030; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4033 = 6'h1 == _T_536 ? _T_21 : _T_20; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4034 = 6'h2 == _T_536 ? _T_22 : _GEN_4033; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4035 = 6'h3 == _T_536 ? _T_23 : _GEN_4034; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4036 = 6'h4 == _T_536 ? _T_24 : _GEN_4035; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4037 = 6'h5 == _T_536 ? _T_25 : _GEN_4036; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4038 = 6'h6 == _T_536 ? _T_26 : _GEN_4037; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4039 = 6'h7 == _T_536 ? _T_27 : _GEN_4038; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4040 = 6'h8 == _T_536 ? _T_28 : _GEN_4039; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4041 = 6'h9 == _T_536 ? _T_29 : _GEN_4040; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4042 = 6'ha == _T_536 ? _T_30 : _GEN_4041; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4043 = 6'hb == _T_536 ? _T_31 : _GEN_4042; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4044 = 6'hc == _T_536 ? _T_32 : _GEN_4043; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4045 = 6'hd == _T_536 ? _T_33 : _GEN_4044; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4046 = 6'he == _T_536 ? _T_34 : _GEN_4045; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4047 = 6'hf == _T_536 ? _T_35 : _GEN_4046; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4048 = 6'h10 == _T_536 ? _T_36 : _GEN_4047; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4049 = 6'h11 == _T_536 ? _T_37 : _GEN_4048; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4050 = 6'h12 == _T_536 ? _T_38 : _GEN_4049; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4051 = 6'h13 == _T_536 ? _T_39 : _GEN_4050; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4052 = 6'h14 == _T_536 ? _T_40 : _GEN_4051; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4053 = 6'h15 == _T_536 ? _T_41 : _GEN_4052; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4054 = 6'h16 == _T_536 ? _T_42 : _GEN_4053; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4055 = 6'h17 == _T_536 ? _T_43 : _GEN_4054; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4056 = 6'h18 == _T_536 ? _T_44 : _GEN_4055; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4057 = 6'h19 == _T_536 ? _T_45 : _GEN_4056; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4058 = 6'h1a == _T_536 ? _T_46 : _GEN_4057; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4059 = 6'h1b == _T_536 ? _T_47 : _GEN_4058; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4060 = 6'h1c == _T_536 ? _T_48 : _GEN_4059; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4061 = 6'h1d == _T_536 ? _T_49 : _GEN_4060; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4062 = 6'h1e == _T_536 ? _T_50 : _GEN_4061; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4063 = 6'h1f == _T_536 ? _T_51 : _GEN_4062; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4064 = 6'h20 == _T_536 ? _T_52 : _GEN_4063; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4065 = 6'h21 == _T_536 ? _T_53 : _GEN_4064; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4066 = 6'h22 == _T_536 ? _T_54 : _GEN_4065; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4067 = 6'h23 == _T_536 ? _T_55 : _GEN_4066; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4068 = 6'h24 == _T_536 ? _T_56 : _GEN_4067; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4069 = 6'h25 == _T_536 ? _T_57 : _GEN_4068; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4070 = 6'h26 == _T_536 ? _T_58 : _GEN_4069; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4071 = 6'h27 == _T_536 ? _T_59 : _GEN_4070; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4072 = 6'h28 == _T_536 ? _T_60 : _GEN_4071; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4073 = 6'h29 == _T_536 ? _T_61 : _GEN_4072; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4074 = 6'h2a == _T_536 ? _T_62 : _GEN_4073; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4075 = 6'h2b == _T_536 ? _T_63 : _GEN_4074; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4076 = 6'h2c == _T_536 ? _T_64 : _GEN_4075; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4077 = 6'h2d == _T_536 ? _T_65 : _GEN_4076; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4078 = 6'h2e == _T_536 ? _T_66 : _GEN_4077; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4079 = 6'h2f == _T_536 ? _T_67 : _GEN_4078; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4080 = 6'h30 == _T_536 ? _T_68 : _GEN_4079; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4081 = 6'h31 == _T_536 ? _T_69 : _GEN_4080; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4082 = 6'h32 == _T_536 ? _T_70 : _GEN_4081; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4083 = 6'h33 == _T_536 ? _T_71 : _GEN_4082; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4084 = 6'h34 == _T_536 ? _T_72 : _GEN_4083; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4085 = 6'h35 == _T_536 ? _T_73 : _GEN_4084; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4086 = 6'h36 == _T_536 ? _T_74 : _GEN_4085; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4087 = 6'h37 == _T_536 ? _T_75 : _GEN_4086; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4088 = 6'h38 == _T_536 ? _T_76 : _GEN_4087; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4089 = 6'h39 == _T_536 ? _T_77 : _GEN_4088; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4090 = 6'h3a == _T_536 ? _T_78 : _GEN_4089; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4091 = 6'h3b == _T_536 ? _T_79 : _GEN_4090; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4092 = 6'h3c == _T_536 ? _T_80 : _GEN_4091; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4093 = 6'h3d == _T_536 ? _T_81 : _GEN_4092; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4094 = 6'h3e == _T_536 ? _T_82 : _GEN_4093; // @[execute.scala 79:10:@2074.4]
  assign _GEN_4095 = 6'h3f == _T_536 ? _T_83 : _GEN_4094; // @[execute.scala 79:10:@2074.4]
  assign _T_538 = _T_528 ? _GEN_4031 : _GEN_4095; // @[execute.scala 79:10:@2074.4]
  assign _T_540 = io_amount < 6'h20; // @[execute.scala 79:15:@2075.4]
  assign _T_542 = io_amount - 6'h20; // @[execute.scala 79:37:@2076.4]
  assign _T_543 = $unsigned(_T_542); // @[execute.scala 79:37:@2077.4]
  assign _T_544 = _T_543[5:0]; // @[execute.scala 79:37:@2078.4]
  assign _T_547 = 6'h20 + io_amount; // @[execute.scala 79:60:@2079.4]
  assign _T_548 = 6'h20 + io_amount; // @[execute.scala 79:60:@2080.4]
  assign _GEN_4097 = 6'h1 == _T_544 ? _T_21 : _T_20; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4098 = 6'h2 == _T_544 ? _T_22 : _GEN_4097; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4099 = 6'h3 == _T_544 ? _T_23 : _GEN_4098; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4100 = 6'h4 == _T_544 ? _T_24 : _GEN_4099; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4101 = 6'h5 == _T_544 ? _T_25 : _GEN_4100; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4102 = 6'h6 == _T_544 ? _T_26 : _GEN_4101; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4103 = 6'h7 == _T_544 ? _T_27 : _GEN_4102; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4104 = 6'h8 == _T_544 ? _T_28 : _GEN_4103; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4105 = 6'h9 == _T_544 ? _T_29 : _GEN_4104; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4106 = 6'ha == _T_544 ? _T_30 : _GEN_4105; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4107 = 6'hb == _T_544 ? _T_31 : _GEN_4106; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4108 = 6'hc == _T_544 ? _T_32 : _GEN_4107; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4109 = 6'hd == _T_544 ? _T_33 : _GEN_4108; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4110 = 6'he == _T_544 ? _T_34 : _GEN_4109; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4111 = 6'hf == _T_544 ? _T_35 : _GEN_4110; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4112 = 6'h10 == _T_544 ? _T_36 : _GEN_4111; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4113 = 6'h11 == _T_544 ? _T_37 : _GEN_4112; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4114 = 6'h12 == _T_544 ? _T_38 : _GEN_4113; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4115 = 6'h13 == _T_544 ? _T_39 : _GEN_4114; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4116 = 6'h14 == _T_544 ? _T_40 : _GEN_4115; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4117 = 6'h15 == _T_544 ? _T_41 : _GEN_4116; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4118 = 6'h16 == _T_544 ? _T_42 : _GEN_4117; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4119 = 6'h17 == _T_544 ? _T_43 : _GEN_4118; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4120 = 6'h18 == _T_544 ? _T_44 : _GEN_4119; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4121 = 6'h19 == _T_544 ? _T_45 : _GEN_4120; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4122 = 6'h1a == _T_544 ? _T_46 : _GEN_4121; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4123 = 6'h1b == _T_544 ? _T_47 : _GEN_4122; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4124 = 6'h1c == _T_544 ? _T_48 : _GEN_4123; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4125 = 6'h1d == _T_544 ? _T_49 : _GEN_4124; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4126 = 6'h1e == _T_544 ? _T_50 : _GEN_4125; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4127 = 6'h1f == _T_544 ? _T_51 : _GEN_4126; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4128 = 6'h20 == _T_544 ? _T_52 : _GEN_4127; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4129 = 6'h21 == _T_544 ? _T_53 : _GEN_4128; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4130 = 6'h22 == _T_544 ? _T_54 : _GEN_4129; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4131 = 6'h23 == _T_544 ? _T_55 : _GEN_4130; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4132 = 6'h24 == _T_544 ? _T_56 : _GEN_4131; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4133 = 6'h25 == _T_544 ? _T_57 : _GEN_4132; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4134 = 6'h26 == _T_544 ? _T_58 : _GEN_4133; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4135 = 6'h27 == _T_544 ? _T_59 : _GEN_4134; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4136 = 6'h28 == _T_544 ? _T_60 : _GEN_4135; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4137 = 6'h29 == _T_544 ? _T_61 : _GEN_4136; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4138 = 6'h2a == _T_544 ? _T_62 : _GEN_4137; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4139 = 6'h2b == _T_544 ? _T_63 : _GEN_4138; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4140 = 6'h2c == _T_544 ? _T_64 : _GEN_4139; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4141 = 6'h2d == _T_544 ? _T_65 : _GEN_4140; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4142 = 6'h2e == _T_544 ? _T_66 : _GEN_4141; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4143 = 6'h2f == _T_544 ? _T_67 : _GEN_4142; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4144 = 6'h30 == _T_544 ? _T_68 : _GEN_4143; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4145 = 6'h31 == _T_544 ? _T_69 : _GEN_4144; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4146 = 6'h32 == _T_544 ? _T_70 : _GEN_4145; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4147 = 6'h33 == _T_544 ? _T_71 : _GEN_4146; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4148 = 6'h34 == _T_544 ? _T_72 : _GEN_4147; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4149 = 6'h35 == _T_544 ? _T_73 : _GEN_4148; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4150 = 6'h36 == _T_544 ? _T_74 : _GEN_4149; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4151 = 6'h37 == _T_544 ? _T_75 : _GEN_4150; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4152 = 6'h38 == _T_544 ? _T_76 : _GEN_4151; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4153 = 6'h39 == _T_544 ? _T_77 : _GEN_4152; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4154 = 6'h3a == _T_544 ? _T_78 : _GEN_4153; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4155 = 6'h3b == _T_544 ? _T_79 : _GEN_4154; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4156 = 6'h3c == _T_544 ? _T_80 : _GEN_4155; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4157 = 6'h3d == _T_544 ? _T_81 : _GEN_4156; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4158 = 6'h3e == _T_544 ? _T_82 : _GEN_4157; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4159 = 6'h3f == _T_544 ? _T_83 : _GEN_4158; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4161 = 6'h1 == _T_548 ? _T_21 : _T_20; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4162 = 6'h2 == _T_548 ? _T_22 : _GEN_4161; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4163 = 6'h3 == _T_548 ? _T_23 : _GEN_4162; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4164 = 6'h4 == _T_548 ? _T_24 : _GEN_4163; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4165 = 6'h5 == _T_548 ? _T_25 : _GEN_4164; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4166 = 6'h6 == _T_548 ? _T_26 : _GEN_4165; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4167 = 6'h7 == _T_548 ? _T_27 : _GEN_4166; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4168 = 6'h8 == _T_548 ? _T_28 : _GEN_4167; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4169 = 6'h9 == _T_548 ? _T_29 : _GEN_4168; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4170 = 6'ha == _T_548 ? _T_30 : _GEN_4169; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4171 = 6'hb == _T_548 ? _T_31 : _GEN_4170; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4172 = 6'hc == _T_548 ? _T_32 : _GEN_4171; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4173 = 6'hd == _T_548 ? _T_33 : _GEN_4172; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4174 = 6'he == _T_548 ? _T_34 : _GEN_4173; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4175 = 6'hf == _T_548 ? _T_35 : _GEN_4174; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4176 = 6'h10 == _T_548 ? _T_36 : _GEN_4175; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4177 = 6'h11 == _T_548 ? _T_37 : _GEN_4176; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4178 = 6'h12 == _T_548 ? _T_38 : _GEN_4177; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4179 = 6'h13 == _T_548 ? _T_39 : _GEN_4178; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4180 = 6'h14 == _T_548 ? _T_40 : _GEN_4179; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4181 = 6'h15 == _T_548 ? _T_41 : _GEN_4180; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4182 = 6'h16 == _T_548 ? _T_42 : _GEN_4181; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4183 = 6'h17 == _T_548 ? _T_43 : _GEN_4182; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4184 = 6'h18 == _T_548 ? _T_44 : _GEN_4183; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4185 = 6'h19 == _T_548 ? _T_45 : _GEN_4184; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4186 = 6'h1a == _T_548 ? _T_46 : _GEN_4185; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4187 = 6'h1b == _T_548 ? _T_47 : _GEN_4186; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4188 = 6'h1c == _T_548 ? _T_48 : _GEN_4187; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4189 = 6'h1d == _T_548 ? _T_49 : _GEN_4188; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4190 = 6'h1e == _T_548 ? _T_50 : _GEN_4189; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4191 = 6'h1f == _T_548 ? _T_51 : _GEN_4190; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4192 = 6'h20 == _T_548 ? _T_52 : _GEN_4191; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4193 = 6'h21 == _T_548 ? _T_53 : _GEN_4192; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4194 = 6'h22 == _T_548 ? _T_54 : _GEN_4193; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4195 = 6'h23 == _T_548 ? _T_55 : _GEN_4194; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4196 = 6'h24 == _T_548 ? _T_56 : _GEN_4195; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4197 = 6'h25 == _T_548 ? _T_57 : _GEN_4196; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4198 = 6'h26 == _T_548 ? _T_58 : _GEN_4197; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4199 = 6'h27 == _T_548 ? _T_59 : _GEN_4198; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4200 = 6'h28 == _T_548 ? _T_60 : _GEN_4199; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4201 = 6'h29 == _T_548 ? _T_61 : _GEN_4200; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4202 = 6'h2a == _T_548 ? _T_62 : _GEN_4201; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4203 = 6'h2b == _T_548 ? _T_63 : _GEN_4202; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4204 = 6'h2c == _T_548 ? _T_64 : _GEN_4203; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4205 = 6'h2d == _T_548 ? _T_65 : _GEN_4204; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4206 = 6'h2e == _T_548 ? _T_66 : _GEN_4205; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4207 = 6'h2f == _T_548 ? _T_67 : _GEN_4206; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4208 = 6'h30 == _T_548 ? _T_68 : _GEN_4207; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4209 = 6'h31 == _T_548 ? _T_69 : _GEN_4208; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4210 = 6'h32 == _T_548 ? _T_70 : _GEN_4209; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4211 = 6'h33 == _T_548 ? _T_71 : _GEN_4210; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4212 = 6'h34 == _T_548 ? _T_72 : _GEN_4211; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4213 = 6'h35 == _T_548 ? _T_73 : _GEN_4212; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4214 = 6'h36 == _T_548 ? _T_74 : _GEN_4213; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4215 = 6'h37 == _T_548 ? _T_75 : _GEN_4214; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4216 = 6'h38 == _T_548 ? _T_76 : _GEN_4215; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4217 = 6'h39 == _T_548 ? _T_77 : _GEN_4216; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4218 = 6'h3a == _T_548 ? _T_78 : _GEN_4217; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4219 = 6'h3b == _T_548 ? _T_79 : _GEN_4218; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4220 = 6'h3c == _T_548 ? _T_80 : _GEN_4219; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4221 = 6'h3d == _T_548 ? _T_81 : _GEN_4220; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4222 = 6'h3e == _T_548 ? _T_82 : _GEN_4221; // @[execute.scala 79:10:@2081.4]
  assign _GEN_4223 = 6'h3f == _T_548 ? _T_83 : _GEN_4222; // @[execute.scala 79:10:@2081.4]
  assign _T_550 = _T_540 ? _GEN_4159 : _GEN_4223; // @[execute.scala 79:10:@2081.4]
  assign _T_552 = io_amount < 6'h1f; // @[execute.scala 79:15:@2082.4]
  assign _T_554 = io_amount - 6'h1f; // @[execute.scala 79:37:@2083.4]
  assign _T_555 = $unsigned(_T_554); // @[execute.scala 79:37:@2084.4]
  assign _T_556 = _T_555[5:0]; // @[execute.scala 79:37:@2085.4]
  assign _T_559 = 6'h21 + io_amount; // @[execute.scala 79:60:@2086.4]
  assign _T_560 = 6'h21 + io_amount; // @[execute.scala 79:60:@2087.4]
  assign _GEN_4225 = 6'h1 == _T_556 ? _T_21 : _T_20; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4226 = 6'h2 == _T_556 ? _T_22 : _GEN_4225; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4227 = 6'h3 == _T_556 ? _T_23 : _GEN_4226; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4228 = 6'h4 == _T_556 ? _T_24 : _GEN_4227; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4229 = 6'h5 == _T_556 ? _T_25 : _GEN_4228; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4230 = 6'h6 == _T_556 ? _T_26 : _GEN_4229; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4231 = 6'h7 == _T_556 ? _T_27 : _GEN_4230; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4232 = 6'h8 == _T_556 ? _T_28 : _GEN_4231; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4233 = 6'h9 == _T_556 ? _T_29 : _GEN_4232; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4234 = 6'ha == _T_556 ? _T_30 : _GEN_4233; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4235 = 6'hb == _T_556 ? _T_31 : _GEN_4234; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4236 = 6'hc == _T_556 ? _T_32 : _GEN_4235; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4237 = 6'hd == _T_556 ? _T_33 : _GEN_4236; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4238 = 6'he == _T_556 ? _T_34 : _GEN_4237; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4239 = 6'hf == _T_556 ? _T_35 : _GEN_4238; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4240 = 6'h10 == _T_556 ? _T_36 : _GEN_4239; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4241 = 6'h11 == _T_556 ? _T_37 : _GEN_4240; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4242 = 6'h12 == _T_556 ? _T_38 : _GEN_4241; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4243 = 6'h13 == _T_556 ? _T_39 : _GEN_4242; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4244 = 6'h14 == _T_556 ? _T_40 : _GEN_4243; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4245 = 6'h15 == _T_556 ? _T_41 : _GEN_4244; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4246 = 6'h16 == _T_556 ? _T_42 : _GEN_4245; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4247 = 6'h17 == _T_556 ? _T_43 : _GEN_4246; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4248 = 6'h18 == _T_556 ? _T_44 : _GEN_4247; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4249 = 6'h19 == _T_556 ? _T_45 : _GEN_4248; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4250 = 6'h1a == _T_556 ? _T_46 : _GEN_4249; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4251 = 6'h1b == _T_556 ? _T_47 : _GEN_4250; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4252 = 6'h1c == _T_556 ? _T_48 : _GEN_4251; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4253 = 6'h1d == _T_556 ? _T_49 : _GEN_4252; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4254 = 6'h1e == _T_556 ? _T_50 : _GEN_4253; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4255 = 6'h1f == _T_556 ? _T_51 : _GEN_4254; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4256 = 6'h20 == _T_556 ? _T_52 : _GEN_4255; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4257 = 6'h21 == _T_556 ? _T_53 : _GEN_4256; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4258 = 6'h22 == _T_556 ? _T_54 : _GEN_4257; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4259 = 6'h23 == _T_556 ? _T_55 : _GEN_4258; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4260 = 6'h24 == _T_556 ? _T_56 : _GEN_4259; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4261 = 6'h25 == _T_556 ? _T_57 : _GEN_4260; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4262 = 6'h26 == _T_556 ? _T_58 : _GEN_4261; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4263 = 6'h27 == _T_556 ? _T_59 : _GEN_4262; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4264 = 6'h28 == _T_556 ? _T_60 : _GEN_4263; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4265 = 6'h29 == _T_556 ? _T_61 : _GEN_4264; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4266 = 6'h2a == _T_556 ? _T_62 : _GEN_4265; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4267 = 6'h2b == _T_556 ? _T_63 : _GEN_4266; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4268 = 6'h2c == _T_556 ? _T_64 : _GEN_4267; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4269 = 6'h2d == _T_556 ? _T_65 : _GEN_4268; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4270 = 6'h2e == _T_556 ? _T_66 : _GEN_4269; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4271 = 6'h2f == _T_556 ? _T_67 : _GEN_4270; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4272 = 6'h30 == _T_556 ? _T_68 : _GEN_4271; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4273 = 6'h31 == _T_556 ? _T_69 : _GEN_4272; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4274 = 6'h32 == _T_556 ? _T_70 : _GEN_4273; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4275 = 6'h33 == _T_556 ? _T_71 : _GEN_4274; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4276 = 6'h34 == _T_556 ? _T_72 : _GEN_4275; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4277 = 6'h35 == _T_556 ? _T_73 : _GEN_4276; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4278 = 6'h36 == _T_556 ? _T_74 : _GEN_4277; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4279 = 6'h37 == _T_556 ? _T_75 : _GEN_4278; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4280 = 6'h38 == _T_556 ? _T_76 : _GEN_4279; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4281 = 6'h39 == _T_556 ? _T_77 : _GEN_4280; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4282 = 6'h3a == _T_556 ? _T_78 : _GEN_4281; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4283 = 6'h3b == _T_556 ? _T_79 : _GEN_4282; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4284 = 6'h3c == _T_556 ? _T_80 : _GEN_4283; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4285 = 6'h3d == _T_556 ? _T_81 : _GEN_4284; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4286 = 6'h3e == _T_556 ? _T_82 : _GEN_4285; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4287 = 6'h3f == _T_556 ? _T_83 : _GEN_4286; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4289 = 6'h1 == _T_560 ? _T_21 : _T_20; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4290 = 6'h2 == _T_560 ? _T_22 : _GEN_4289; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4291 = 6'h3 == _T_560 ? _T_23 : _GEN_4290; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4292 = 6'h4 == _T_560 ? _T_24 : _GEN_4291; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4293 = 6'h5 == _T_560 ? _T_25 : _GEN_4292; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4294 = 6'h6 == _T_560 ? _T_26 : _GEN_4293; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4295 = 6'h7 == _T_560 ? _T_27 : _GEN_4294; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4296 = 6'h8 == _T_560 ? _T_28 : _GEN_4295; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4297 = 6'h9 == _T_560 ? _T_29 : _GEN_4296; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4298 = 6'ha == _T_560 ? _T_30 : _GEN_4297; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4299 = 6'hb == _T_560 ? _T_31 : _GEN_4298; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4300 = 6'hc == _T_560 ? _T_32 : _GEN_4299; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4301 = 6'hd == _T_560 ? _T_33 : _GEN_4300; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4302 = 6'he == _T_560 ? _T_34 : _GEN_4301; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4303 = 6'hf == _T_560 ? _T_35 : _GEN_4302; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4304 = 6'h10 == _T_560 ? _T_36 : _GEN_4303; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4305 = 6'h11 == _T_560 ? _T_37 : _GEN_4304; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4306 = 6'h12 == _T_560 ? _T_38 : _GEN_4305; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4307 = 6'h13 == _T_560 ? _T_39 : _GEN_4306; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4308 = 6'h14 == _T_560 ? _T_40 : _GEN_4307; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4309 = 6'h15 == _T_560 ? _T_41 : _GEN_4308; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4310 = 6'h16 == _T_560 ? _T_42 : _GEN_4309; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4311 = 6'h17 == _T_560 ? _T_43 : _GEN_4310; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4312 = 6'h18 == _T_560 ? _T_44 : _GEN_4311; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4313 = 6'h19 == _T_560 ? _T_45 : _GEN_4312; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4314 = 6'h1a == _T_560 ? _T_46 : _GEN_4313; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4315 = 6'h1b == _T_560 ? _T_47 : _GEN_4314; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4316 = 6'h1c == _T_560 ? _T_48 : _GEN_4315; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4317 = 6'h1d == _T_560 ? _T_49 : _GEN_4316; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4318 = 6'h1e == _T_560 ? _T_50 : _GEN_4317; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4319 = 6'h1f == _T_560 ? _T_51 : _GEN_4318; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4320 = 6'h20 == _T_560 ? _T_52 : _GEN_4319; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4321 = 6'h21 == _T_560 ? _T_53 : _GEN_4320; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4322 = 6'h22 == _T_560 ? _T_54 : _GEN_4321; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4323 = 6'h23 == _T_560 ? _T_55 : _GEN_4322; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4324 = 6'h24 == _T_560 ? _T_56 : _GEN_4323; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4325 = 6'h25 == _T_560 ? _T_57 : _GEN_4324; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4326 = 6'h26 == _T_560 ? _T_58 : _GEN_4325; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4327 = 6'h27 == _T_560 ? _T_59 : _GEN_4326; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4328 = 6'h28 == _T_560 ? _T_60 : _GEN_4327; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4329 = 6'h29 == _T_560 ? _T_61 : _GEN_4328; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4330 = 6'h2a == _T_560 ? _T_62 : _GEN_4329; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4331 = 6'h2b == _T_560 ? _T_63 : _GEN_4330; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4332 = 6'h2c == _T_560 ? _T_64 : _GEN_4331; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4333 = 6'h2d == _T_560 ? _T_65 : _GEN_4332; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4334 = 6'h2e == _T_560 ? _T_66 : _GEN_4333; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4335 = 6'h2f == _T_560 ? _T_67 : _GEN_4334; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4336 = 6'h30 == _T_560 ? _T_68 : _GEN_4335; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4337 = 6'h31 == _T_560 ? _T_69 : _GEN_4336; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4338 = 6'h32 == _T_560 ? _T_70 : _GEN_4337; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4339 = 6'h33 == _T_560 ? _T_71 : _GEN_4338; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4340 = 6'h34 == _T_560 ? _T_72 : _GEN_4339; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4341 = 6'h35 == _T_560 ? _T_73 : _GEN_4340; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4342 = 6'h36 == _T_560 ? _T_74 : _GEN_4341; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4343 = 6'h37 == _T_560 ? _T_75 : _GEN_4342; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4344 = 6'h38 == _T_560 ? _T_76 : _GEN_4343; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4345 = 6'h39 == _T_560 ? _T_77 : _GEN_4344; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4346 = 6'h3a == _T_560 ? _T_78 : _GEN_4345; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4347 = 6'h3b == _T_560 ? _T_79 : _GEN_4346; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4348 = 6'h3c == _T_560 ? _T_80 : _GEN_4347; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4349 = 6'h3d == _T_560 ? _T_81 : _GEN_4348; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4350 = 6'h3e == _T_560 ? _T_82 : _GEN_4349; // @[execute.scala 79:10:@2088.4]
  assign _GEN_4351 = 6'h3f == _T_560 ? _T_83 : _GEN_4350; // @[execute.scala 79:10:@2088.4]
  assign _T_562 = _T_552 ? _GEN_4287 : _GEN_4351; // @[execute.scala 79:10:@2088.4]
  assign _T_564 = io_amount < 6'h1e; // @[execute.scala 79:15:@2089.4]
  assign _T_566 = io_amount - 6'h1e; // @[execute.scala 79:37:@2090.4]
  assign _T_567 = $unsigned(_T_566); // @[execute.scala 79:37:@2091.4]
  assign _T_568 = _T_567[5:0]; // @[execute.scala 79:37:@2092.4]
  assign _T_571 = 6'h22 + io_amount; // @[execute.scala 79:60:@2093.4]
  assign _T_572 = 6'h22 + io_amount; // @[execute.scala 79:60:@2094.4]
  assign _GEN_4353 = 6'h1 == _T_568 ? _T_21 : _T_20; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4354 = 6'h2 == _T_568 ? _T_22 : _GEN_4353; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4355 = 6'h3 == _T_568 ? _T_23 : _GEN_4354; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4356 = 6'h4 == _T_568 ? _T_24 : _GEN_4355; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4357 = 6'h5 == _T_568 ? _T_25 : _GEN_4356; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4358 = 6'h6 == _T_568 ? _T_26 : _GEN_4357; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4359 = 6'h7 == _T_568 ? _T_27 : _GEN_4358; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4360 = 6'h8 == _T_568 ? _T_28 : _GEN_4359; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4361 = 6'h9 == _T_568 ? _T_29 : _GEN_4360; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4362 = 6'ha == _T_568 ? _T_30 : _GEN_4361; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4363 = 6'hb == _T_568 ? _T_31 : _GEN_4362; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4364 = 6'hc == _T_568 ? _T_32 : _GEN_4363; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4365 = 6'hd == _T_568 ? _T_33 : _GEN_4364; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4366 = 6'he == _T_568 ? _T_34 : _GEN_4365; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4367 = 6'hf == _T_568 ? _T_35 : _GEN_4366; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4368 = 6'h10 == _T_568 ? _T_36 : _GEN_4367; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4369 = 6'h11 == _T_568 ? _T_37 : _GEN_4368; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4370 = 6'h12 == _T_568 ? _T_38 : _GEN_4369; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4371 = 6'h13 == _T_568 ? _T_39 : _GEN_4370; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4372 = 6'h14 == _T_568 ? _T_40 : _GEN_4371; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4373 = 6'h15 == _T_568 ? _T_41 : _GEN_4372; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4374 = 6'h16 == _T_568 ? _T_42 : _GEN_4373; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4375 = 6'h17 == _T_568 ? _T_43 : _GEN_4374; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4376 = 6'h18 == _T_568 ? _T_44 : _GEN_4375; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4377 = 6'h19 == _T_568 ? _T_45 : _GEN_4376; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4378 = 6'h1a == _T_568 ? _T_46 : _GEN_4377; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4379 = 6'h1b == _T_568 ? _T_47 : _GEN_4378; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4380 = 6'h1c == _T_568 ? _T_48 : _GEN_4379; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4381 = 6'h1d == _T_568 ? _T_49 : _GEN_4380; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4382 = 6'h1e == _T_568 ? _T_50 : _GEN_4381; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4383 = 6'h1f == _T_568 ? _T_51 : _GEN_4382; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4384 = 6'h20 == _T_568 ? _T_52 : _GEN_4383; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4385 = 6'h21 == _T_568 ? _T_53 : _GEN_4384; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4386 = 6'h22 == _T_568 ? _T_54 : _GEN_4385; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4387 = 6'h23 == _T_568 ? _T_55 : _GEN_4386; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4388 = 6'h24 == _T_568 ? _T_56 : _GEN_4387; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4389 = 6'h25 == _T_568 ? _T_57 : _GEN_4388; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4390 = 6'h26 == _T_568 ? _T_58 : _GEN_4389; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4391 = 6'h27 == _T_568 ? _T_59 : _GEN_4390; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4392 = 6'h28 == _T_568 ? _T_60 : _GEN_4391; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4393 = 6'h29 == _T_568 ? _T_61 : _GEN_4392; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4394 = 6'h2a == _T_568 ? _T_62 : _GEN_4393; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4395 = 6'h2b == _T_568 ? _T_63 : _GEN_4394; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4396 = 6'h2c == _T_568 ? _T_64 : _GEN_4395; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4397 = 6'h2d == _T_568 ? _T_65 : _GEN_4396; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4398 = 6'h2e == _T_568 ? _T_66 : _GEN_4397; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4399 = 6'h2f == _T_568 ? _T_67 : _GEN_4398; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4400 = 6'h30 == _T_568 ? _T_68 : _GEN_4399; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4401 = 6'h31 == _T_568 ? _T_69 : _GEN_4400; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4402 = 6'h32 == _T_568 ? _T_70 : _GEN_4401; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4403 = 6'h33 == _T_568 ? _T_71 : _GEN_4402; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4404 = 6'h34 == _T_568 ? _T_72 : _GEN_4403; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4405 = 6'h35 == _T_568 ? _T_73 : _GEN_4404; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4406 = 6'h36 == _T_568 ? _T_74 : _GEN_4405; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4407 = 6'h37 == _T_568 ? _T_75 : _GEN_4406; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4408 = 6'h38 == _T_568 ? _T_76 : _GEN_4407; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4409 = 6'h39 == _T_568 ? _T_77 : _GEN_4408; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4410 = 6'h3a == _T_568 ? _T_78 : _GEN_4409; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4411 = 6'h3b == _T_568 ? _T_79 : _GEN_4410; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4412 = 6'h3c == _T_568 ? _T_80 : _GEN_4411; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4413 = 6'h3d == _T_568 ? _T_81 : _GEN_4412; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4414 = 6'h3e == _T_568 ? _T_82 : _GEN_4413; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4415 = 6'h3f == _T_568 ? _T_83 : _GEN_4414; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4417 = 6'h1 == _T_572 ? _T_21 : _T_20; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4418 = 6'h2 == _T_572 ? _T_22 : _GEN_4417; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4419 = 6'h3 == _T_572 ? _T_23 : _GEN_4418; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4420 = 6'h4 == _T_572 ? _T_24 : _GEN_4419; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4421 = 6'h5 == _T_572 ? _T_25 : _GEN_4420; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4422 = 6'h6 == _T_572 ? _T_26 : _GEN_4421; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4423 = 6'h7 == _T_572 ? _T_27 : _GEN_4422; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4424 = 6'h8 == _T_572 ? _T_28 : _GEN_4423; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4425 = 6'h9 == _T_572 ? _T_29 : _GEN_4424; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4426 = 6'ha == _T_572 ? _T_30 : _GEN_4425; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4427 = 6'hb == _T_572 ? _T_31 : _GEN_4426; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4428 = 6'hc == _T_572 ? _T_32 : _GEN_4427; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4429 = 6'hd == _T_572 ? _T_33 : _GEN_4428; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4430 = 6'he == _T_572 ? _T_34 : _GEN_4429; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4431 = 6'hf == _T_572 ? _T_35 : _GEN_4430; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4432 = 6'h10 == _T_572 ? _T_36 : _GEN_4431; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4433 = 6'h11 == _T_572 ? _T_37 : _GEN_4432; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4434 = 6'h12 == _T_572 ? _T_38 : _GEN_4433; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4435 = 6'h13 == _T_572 ? _T_39 : _GEN_4434; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4436 = 6'h14 == _T_572 ? _T_40 : _GEN_4435; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4437 = 6'h15 == _T_572 ? _T_41 : _GEN_4436; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4438 = 6'h16 == _T_572 ? _T_42 : _GEN_4437; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4439 = 6'h17 == _T_572 ? _T_43 : _GEN_4438; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4440 = 6'h18 == _T_572 ? _T_44 : _GEN_4439; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4441 = 6'h19 == _T_572 ? _T_45 : _GEN_4440; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4442 = 6'h1a == _T_572 ? _T_46 : _GEN_4441; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4443 = 6'h1b == _T_572 ? _T_47 : _GEN_4442; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4444 = 6'h1c == _T_572 ? _T_48 : _GEN_4443; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4445 = 6'h1d == _T_572 ? _T_49 : _GEN_4444; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4446 = 6'h1e == _T_572 ? _T_50 : _GEN_4445; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4447 = 6'h1f == _T_572 ? _T_51 : _GEN_4446; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4448 = 6'h20 == _T_572 ? _T_52 : _GEN_4447; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4449 = 6'h21 == _T_572 ? _T_53 : _GEN_4448; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4450 = 6'h22 == _T_572 ? _T_54 : _GEN_4449; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4451 = 6'h23 == _T_572 ? _T_55 : _GEN_4450; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4452 = 6'h24 == _T_572 ? _T_56 : _GEN_4451; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4453 = 6'h25 == _T_572 ? _T_57 : _GEN_4452; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4454 = 6'h26 == _T_572 ? _T_58 : _GEN_4453; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4455 = 6'h27 == _T_572 ? _T_59 : _GEN_4454; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4456 = 6'h28 == _T_572 ? _T_60 : _GEN_4455; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4457 = 6'h29 == _T_572 ? _T_61 : _GEN_4456; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4458 = 6'h2a == _T_572 ? _T_62 : _GEN_4457; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4459 = 6'h2b == _T_572 ? _T_63 : _GEN_4458; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4460 = 6'h2c == _T_572 ? _T_64 : _GEN_4459; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4461 = 6'h2d == _T_572 ? _T_65 : _GEN_4460; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4462 = 6'h2e == _T_572 ? _T_66 : _GEN_4461; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4463 = 6'h2f == _T_572 ? _T_67 : _GEN_4462; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4464 = 6'h30 == _T_572 ? _T_68 : _GEN_4463; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4465 = 6'h31 == _T_572 ? _T_69 : _GEN_4464; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4466 = 6'h32 == _T_572 ? _T_70 : _GEN_4465; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4467 = 6'h33 == _T_572 ? _T_71 : _GEN_4466; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4468 = 6'h34 == _T_572 ? _T_72 : _GEN_4467; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4469 = 6'h35 == _T_572 ? _T_73 : _GEN_4468; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4470 = 6'h36 == _T_572 ? _T_74 : _GEN_4469; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4471 = 6'h37 == _T_572 ? _T_75 : _GEN_4470; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4472 = 6'h38 == _T_572 ? _T_76 : _GEN_4471; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4473 = 6'h39 == _T_572 ? _T_77 : _GEN_4472; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4474 = 6'h3a == _T_572 ? _T_78 : _GEN_4473; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4475 = 6'h3b == _T_572 ? _T_79 : _GEN_4474; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4476 = 6'h3c == _T_572 ? _T_80 : _GEN_4475; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4477 = 6'h3d == _T_572 ? _T_81 : _GEN_4476; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4478 = 6'h3e == _T_572 ? _T_82 : _GEN_4477; // @[execute.scala 79:10:@2095.4]
  assign _GEN_4479 = 6'h3f == _T_572 ? _T_83 : _GEN_4478; // @[execute.scala 79:10:@2095.4]
  assign _T_574 = _T_564 ? _GEN_4415 : _GEN_4479; // @[execute.scala 79:10:@2095.4]
  assign _T_576 = io_amount < 6'h1d; // @[execute.scala 79:15:@2096.4]
  assign _T_578 = io_amount - 6'h1d; // @[execute.scala 79:37:@2097.4]
  assign _T_579 = $unsigned(_T_578); // @[execute.scala 79:37:@2098.4]
  assign _T_580 = _T_579[5:0]; // @[execute.scala 79:37:@2099.4]
  assign _T_583 = 6'h23 + io_amount; // @[execute.scala 79:60:@2100.4]
  assign _T_584 = 6'h23 + io_amount; // @[execute.scala 79:60:@2101.4]
  assign _GEN_4481 = 6'h1 == _T_580 ? _T_21 : _T_20; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4482 = 6'h2 == _T_580 ? _T_22 : _GEN_4481; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4483 = 6'h3 == _T_580 ? _T_23 : _GEN_4482; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4484 = 6'h4 == _T_580 ? _T_24 : _GEN_4483; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4485 = 6'h5 == _T_580 ? _T_25 : _GEN_4484; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4486 = 6'h6 == _T_580 ? _T_26 : _GEN_4485; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4487 = 6'h7 == _T_580 ? _T_27 : _GEN_4486; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4488 = 6'h8 == _T_580 ? _T_28 : _GEN_4487; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4489 = 6'h9 == _T_580 ? _T_29 : _GEN_4488; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4490 = 6'ha == _T_580 ? _T_30 : _GEN_4489; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4491 = 6'hb == _T_580 ? _T_31 : _GEN_4490; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4492 = 6'hc == _T_580 ? _T_32 : _GEN_4491; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4493 = 6'hd == _T_580 ? _T_33 : _GEN_4492; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4494 = 6'he == _T_580 ? _T_34 : _GEN_4493; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4495 = 6'hf == _T_580 ? _T_35 : _GEN_4494; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4496 = 6'h10 == _T_580 ? _T_36 : _GEN_4495; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4497 = 6'h11 == _T_580 ? _T_37 : _GEN_4496; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4498 = 6'h12 == _T_580 ? _T_38 : _GEN_4497; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4499 = 6'h13 == _T_580 ? _T_39 : _GEN_4498; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4500 = 6'h14 == _T_580 ? _T_40 : _GEN_4499; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4501 = 6'h15 == _T_580 ? _T_41 : _GEN_4500; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4502 = 6'h16 == _T_580 ? _T_42 : _GEN_4501; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4503 = 6'h17 == _T_580 ? _T_43 : _GEN_4502; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4504 = 6'h18 == _T_580 ? _T_44 : _GEN_4503; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4505 = 6'h19 == _T_580 ? _T_45 : _GEN_4504; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4506 = 6'h1a == _T_580 ? _T_46 : _GEN_4505; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4507 = 6'h1b == _T_580 ? _T_47 : _GEN_4506; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4508 = 6'h1c == _T_580 ? _T_48 : _GEN_4507; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4509 = 6'h1d == _T_580 ? _T_49 : _GEN_4508; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4510 = 6'h1e == _T_580 ? _T_50 : _GEN_4509; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4511 = 6'h1f == _T_580 ? _T_51 : _GEN_4510; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4512 = 6'h20 == _T_580 ? _T_52 : _GEN_4511; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4513 = 6'h21 == _T_580 ? _T_53 : _GEN_4512; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4514 = 6'h22 == _T_580 ? _T_54 : _GEN_4513; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4515 = 6'h23 == _T_580 ? _T_55 : _GEN_4514; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4516 = 6'h24 == _T_580 ? _T_56 : _GEN_4515; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4517 = 6'h25 == _T_580 ? _T_57 : _GEN_4516; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4518 = 6'h26 == _T_580 ? _T_58 : _GEN_4517; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4519 = 6'h27 == _T_580 ? _T_59 : _GEN_4518; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4520 = 6'h28 == _T_580 ? _T_60 : _GEN_4519; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4521 = 6'h29 == _T_580 ? _T_61 : _GEN_4520; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4522 = 6'h2a == _T_580 ? _T_62 : _GEN_4521; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4523 = 6'h2b == _T_580 ? _T_63 : _GEN_4522; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4524 = 6'h2c == _T_580 ? _T_64 : _GEN_4523; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4525 = 6'h2d == _T_580 ? _T_65 : _GEN_4524; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4526 = 6'h2e == _T_580 ? _T_66 : _GEN_4525; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4527 = 6'h2f == _T_580 ? _T_67 : _GEN_4526; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4528 = 6'h30 == _T_580 ? _T_68 : _GEN_4527; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4529 = 6'h31 == _T_580 ? _T_69 : _GEN_4528; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4530 = 6'h32 == _T_580 ? _T_70 : _GEN_4529; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4531 = 6'h33 == _T_580 ? _T_71 : _GEN_4530; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4532 = 6'h34 == _T_580 ? _T_72 : _GEN_4531; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4533 = 6'h35 == _T_580 ? _T_73 : _GEN_4532; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4534 = 6'h36 == _T_580 ? _T_74 : _GEN_4533; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4535 = 6'h37 == _T_580 ? _T_75 : _GEN_4534; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4536 = 6'h38 == _T_580 ? _T_76 : _GEN_4535; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4537 = 6'h39 == _T_580 ? _T_77 : _GEN_4536; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4538 = 6'h3a == _T_580 ? _T_78 : _GEN_4537; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4539 = 6'h3b == _T_580 ? _T_79 : _GEN_4538; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4540 = 6'h3c == _T_580 ? _T_80 : _GEN_4539; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4541 = 6'h3d == _T_580 ? _T_81 : _GEN_4540; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4542 = 6'h3e == _T_580 ? _T_82 : _GEN_4541; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4543 = 6'h3f == _T_580 ? _T_83 : _GEN_4542; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4545 = 6'h1 == _T_584 ? _T_21 : _T_20; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4546 = 6'h2 == _T_584 ? _T_22 : _GEN_4545; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4547 = 6'h3 == _T_584 ? _T_23 : _GEN_4546; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4548 = 6'h4 == _T_584 ? _T_24 : _GEN_4547; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4549 = 6'h5 == _T_584 ? _T_25 : _GEN_4548; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4550 = 6'h6 == _T_584 ? _T_26 : _GEN_4549; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4551 = 6'h7 == _T_584 ? _T_27 : _GEN_4550; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4552 = 6'h8 == _T_584 ? _T_28 : _GEN_4551; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4553 = 6'h9 == _T_584 ? _T_29 : _GEN_4552; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4554 = 6'ha == _T_584 ? _T_30 : _GEN_4553; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4555 = 6'hb == _T_584 ? _T_31 : _GEN_4554; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4556 = 6'hc == _T_584 ? _T_32 : _GEN_4555; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4557 = 6'hd == _T_584 ? _T_33 : _GEN_4556; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4558 = 6'he == _T_584 ? _T_34 : _GEN_4557; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4559 = 6'hf == _T_584 ? _T_35 : _GEN_4558; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4560 = 6'h10 == _T_584 ? _T_36 : _GEN_4559; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4561 = 6'h11 == _T_584 ? _T_37 : _GEN_4560; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4562 = 6'h12 == _T_584 ? _T_38 : _GEN_4561; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4563 = 6'h13 == _T_584 ? _T_39 : _GEN_4562; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4564 = 6'h14 == _T_584 ? _T_40 : _GEN_4563; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4565 = 6'h15 == _T_584 ? _T_41 : _GEN_4564; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4566 = 6'h16 == _T_584 ? _T_42 : _GEN_4565; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4567 = 6'h17 == _T_584 ? _T_43 : _GEN_4566; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4568 = 6'h18 == _T_584 ? _T_44 : _GEN_4567; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4569 = 6'h19 == _T_584 ? _T_45 : _GEN_4568; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4570 = 6'h1a == _T_584 ? _T_46 : _GEN_4569; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4571 = 6'h1b == _T_584 ? _T_47 : _GEN_4570; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4572 = 6'h1c == _T_584 ? _T_48 : _GEN_4571; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4573 = 6'h1d == _T_584 ? _T_49 : _GEN_4572; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4574 = 6'h1e == _T_584 ? _T_50 : _GEN_4573; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4575 = 6'h1f == _T_584 ? _T_51 : _GEN_4574; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4576 = 6'h20 == _T_584 ? _T_52 : _GEN_4575; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4577 = 6'h21 == _T_584 ? _T_53 : _GEN_4576; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4578 = 6'h22 == _T_584 ? _T_54 : _GEN_4577; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4579 = 6'h23 == _T_584 ? _T_55 : _GEN_4578; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4580 = 6'h24 == _T_584 ? _T_56 : _GEN_4579; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4581 = 6'h25 == _T_584 ? _T_57 : _GEN_4580; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4582 = 6'h26 == _T_584 ? _T_58 : _GEN_4581; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4583 = 6'h27 == _T_584 ? _T_59 : _GEN_4582; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4584 = 6'h28 == _T_584 ? _T_60 : _GEN_4583; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4585 = 6'h29 == _T_584 ? _T_61 : _GEN_4584; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4586 = 6'h2a == _T_584 ? _T_62 : _GEN_4585; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4587 = 6'h2b == _T_584 ? _T_63 : _GEN_4586; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4588 = 6'h2c == _T_584 ? _T_64 : _GEN_4587; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4589 = 6'h2d == _T_584 ? _T_65 : _GEN_4588; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4590 = 6'h2e == _T_584 ? _T_66 : _GEN_4589; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4591 = 6'h2f == _T_584 ? _T_67 : _GEN_4590; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4592 = 6'h30 == _T_584 ? _T_68 : _GEN_4591; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4593 = 6'h31 == _T_584 ? _T_69 : _GEN_4592; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4594 = 6'h32 == _T_584 ? _T_70 : _GEN_4593; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4595 = 6'h33 == _T_584 ? _T_71 : _GEN_4594; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4596 = 6'h34 == _T_584 ? _T_72 : _GEN_4595; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4597 = 6'h35 == _T_584 ? _T_73 : _GEN_4596; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4598 = 6'h36 == _T_584 ? _T_74 : _GEN_4597; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4599 = 6'h37 == _T_584 ? _T_75 : _GEN_4598; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4600 = 6'h38 == _T_584 ? _T_76 : _GEN_4599; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4601 = 6'h39 == _T_584 ? _T_77 : _GEN_4600; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4602 = 6'h3a == _T_584 ? _T_78 : _GEN_4601; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4603 = 6'h3b == _T_584 ? _T_79 : _GEN_4602; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4604 = 6'h3c == _T_584 ? _T_80 : _GEN_4603; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4605 = 6'h3d == _T_584 ? _T_81 : _GEN_4604; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4606 = 6'h3e == _T_584 ? _T_82 : _GEN_4605; // @[execute.scala 79:10:@2102.4]
  assign _GEN_4607 = 6'h3f == _T_584 ? _T_83 : _GEN_4606; // @[execute.scala 79:10:@2102.4]
  assign _T_586 = _T_576 ? _GEN_4543 : _GEN_4607; // @[execute.scala 79:10:@2102.4]
  assign _T_588 = io_amount < 6'h1c; // @[execute.scala 79:15:@2103.4]
  assign _T_590 = io_amount - 6'h1c; // @[execute.scala 79:37:@2104.4]
  assign _T_591 = $unsigned(_T_590); // @[execute.scala 79:37:@2105.4]
  assign _T_592 = _T_591[5:0]; // @[execute.scala 79:37:@2106.4]
  assign _T_595 = 6'h24 + io_amount; // @[execute.scala 79:60:@2107.4]
  assign _T_596 = 6'h24 + io_amount; // @[execute.scala 79:60:@2108.4]
  assign _GEN_4609 = 6'h1 == _T_592 ? _T_21 : _T_20; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4610 = 6'h2 == _T_592 ? _T_22 : _GEN_4609; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4611 = 6'h3 == _T_592 ? _T_23 : _GEN_4610; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4612 = 6'h4 == _T_592 ? _T_24 : _GEN_4611; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4613 = 6'h5 == _T_592 ? _T_25 : _GEN_4612; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4614 = 6'h6 == _T_592 ? _T_26 : _GEN_4613; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4615 = 6'h7 == _T_592 ? _T_27 : _GEN_4614; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4616 = 6'h8 == _T_592 ? _T_28 : _GEN_4615; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4617 = 6'h9 == _T_592 ? _T_29 : _GEN_4616; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4618 = 6'ha == _T_592 ? _T_30 : _GEN_4617; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4619 = 6'hb == _T_592 ? _T_31 : _GEN_4618; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4620 = 6'hc == _T_592 ? _T_32 : _GEN_4619; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4621 = 6'hd == _T_592 ? _T_33 : _GEN_4620; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4622 = 6'he == _T_592 ? _T_34 : _GEN_4621; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4623 = 6'hf == _T_592 ? _T_35 : _GEN_4622; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4624 = 6'h10 == _T_592 ? _T_36 : _GEN_4623; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4625 = 6'h11 == _T_592 ? _T_37 : _GEN_4624; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4626 = 6'h12 == _T_592 ? _T_38 : _GEN_4625; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4627 = 6'h13 == _T_592 ? _T_39 : _GEN_4626; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4628 = 6'h14 == _T_592 ? _T_40 : _GEN_4627; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4629 = 6'h15 == _T_592 ? _T_41 : _GEN_4628; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4630 = 6'h16 == _T_592 ? _T_42 : _GEN_4629; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4631 = 6'h17 == _T_592 ? _T_43 : _GEN_4630; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4632 = 6'h18 == _T_592 ? _T_44 : _GEN_4631; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4633 = 6'h19 == _T_592 ? _T_45 : _GEN_4632; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4634 = 6'h1a == _T_592 ? _T_46 : _GEN_4633; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4635 = 6'h1b == _T_592 ? _T_47 : _GEN_4634; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4636 = 6'h1c == _T_592 ? _T_48 : _GEN_4635; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4637 = 6'h1d == _T_592 ? _T_49 : _GEN_4636; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4638 = 6'h1e == _T_592 ? _T_50 : _GEN_4637; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4639 = 6'h1f == _T_592 ? _T_51 : _GEN_4638; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4640 = 6'h20 == _T_592 ? _T_52 : _GEN_4639; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4641 = 6'h21 == _T_592 ? _T_53 : _GEN_4640; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4642 = 6'h22 == _T_592 ? _T_54 : _GEN_4641; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4643 = 6'h23 == _T_592 ? _T_55 : _GEN_4642; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4644 = 6'h24 == _T_592 ? _T_56 : _GEN_4643; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4645 = 6'h25 == _T_592 ? _T_57 : _GEN_4644; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4646 = 6'h26 == _T_592 ? _T_58 : _GEN_4645; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4647 = 6'h27 == _T_592 ? _T_59 : _GEN_4646; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4648 = 6'h28 == _T_592 ? _T_60 : _GEN_4647; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4649 = 6'h29 == _T_592 ? _T_61 : _GEN_4648; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4650 = 6'h2a == _T_592 ? _T_62 : _GEN_4649; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4651 = 6'h2b == _T_592 ? _T_63 : _GEN_4650; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4652 = 6'h2c == _T_592 ? _T_64 : _GEN_4651; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4653 = 6'h2d == _T_592 ? _T_65 : _GEN_4652; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4654 = 6'h2e == _T_592 ? _T_66 : _GEN_4653; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4655 = 6'h2f == _T_592 ? _T_67 : _GEN_4654; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4656 = 6'h30 == _T_592 ? _T_68 : _GEN_4655; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4657 = 6'h31 == _T_592 ? _T_69 : _GEN_4656; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4658 = 6'h32 == _T_592 ? _T_70 : _GEN_4657; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4659 = 6'h33 == _T_592 ? _T_71 : _GEN_4658; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4660 = 6'h34 == _T_592 ? _T_72 : _GEN_4659; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4661 = 6'h35 == _T_592 ? _T_73 : _GEN_4660; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4662 = 6'h36 == _T_592 ? _T_74 : _GEN_4661; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4663 = 6'h37 == _T_592 ? _T_75 : _GEN_4662; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4664 = 6'h38 == _T_592 ? _T_76 : _GEN_4663; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4665 = 6'h39 == _T_592 ? _T_77 : _GEN_4664; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4666 = 6'h3a == _T_592 ? _T_78 : _GEN_4665; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4667 = 6'h3b == _T_592 ? _T_79 : _GEN_4666; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4668 = 6'h3c == _T_592 ? _T_80 : _GEN_4667; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4669 = 6'h3d == _T_592 ? _T_81 : _GEN_4668; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4670 = 6'h3e == _T_592 ? _T_82 : _GEN_4669; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4671 = 6'h3f == _T_592 ? _T_83 : _GEN_4670; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4673 = 6'h1 == _T_596 ? _T_21 : _T_20; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4674 = 6'h2 == _T_596 ? _T_22 : _GEN_4673; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4675 = 6'h3 == _T_596 ? _T_23 : _GEN_4674; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4676 = 6'h4 == _T_596 ? _T_24 : _GEN_4675; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4677 = 6'h5 == _T_596 ? _T_25 : _GEN_4676; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4678 = 6'h6 == _T_596 ? _T_26 : _GEN_4677; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4679 = 6'h7 == _T_596 ? _T_27 : _GEN_4678; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4680 = 6'h8 == _T_596 ? _T_28 : _GEN_4679; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4681 = 6'h9 == _T_596 ? _T_29 : _GEN_4680; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4682 = 6'ha == _T_596 ? _T_30 : _GEN_4681; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4683 = 6'hb == _T_596 ? _T_31 : _GEN_4682; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4684 = 6'hc == _T_596 ? _T_32 : _GEN_4683; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4685 = 6'hd == _T_596 ? _T_33 : _GEN_4684; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4686 = 6'he == _T_596 ? _T_34 : _GEN_4685; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4687 = 6'hf == _T_596 ? _T_35 : _GEN_4686; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4688 = 6'h10 == _T_596 ? _T_36 : _GEN_4687; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4689 = 6'h11 == _T_596 ? _T_37 : _GEN_4688; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4690 = 6'h12 == _T_596 ? _T_38 : _GEN_4689; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4691 = 6'h13 == _T_596 ? _T_39 : _GEN_4690; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4692 = 6'h14 == _T_596 ? _T_40 : _GEN_4691; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4693 = 6'h15 == _T_596 ? _T_41 : _GEN_4692; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4694 = 6'h16 == _T_596 ? _T_42 : _GEN_4693; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4695 = 6'h17 == _T_596 ? _T_43 : _GEN_4694; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4696 = 6'h18 == _T_596 ? _T_44 : _GEN_4695; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4697 = 6'h19 == _T_596 ? _T_45 : _GEN_4696; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4698 = 6'h1a == _T_596 ? _T_46 : _GEN_4697; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4699 = 6'h1b == _T_596 ? _T_47 : _GEN_4698; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4700 = 6'h1c == _T_596 ? _T_48 : _GEN_4699; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4701 = 6'h1d == _T_596 ? _T_49 : _GEN_4700; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4702 = 6'h1e == _T_596 ? _T_50 : _GEN_4701; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4703 = 6'h1f == _T_596 ? _T_51 : _GEN_4702; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4704 = 6'h20 == _T_596 ? _T_52 : _GEN_4703; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4705 = 6'h21 == _T_596 ? _T_53 : _GEN_4704; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4706 = 6'h22 == _T_596 ? _T_54 : _GEN_4705; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4707 = 6'h23 == _T_596 ? _T_55 : _GEN_4706; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4708 = 6'h24 == _T_596 ? _T_56 : _GEN_4707; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4709 = 6'h25 == _T_596 ? _T_57 : _GEN_4708; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4710 = 6'h26 == _T_596 ? _T_58 : _GEN_4709; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4711 = 6'h27 == _T_596 ? _T_59 : _GEN_4710; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4712 = 6'h28 == _T_596 ? _T_60 : _GEN_4711; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4713 = 6'h29 == _T_596 ? _T_61 : _GEN_4712; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4714 = 6'h2a == _T_596 ? _T_62 : _GEN_4713; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4715 = 6'h2b == _T_596 ? _T_63 : _GEN_4714; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4716 = 6'h2c == _T_596 ? _T_64 : _GEN_4715; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4717 = 6'h2d == _T_596 ? _T_65 : _GEN_4716; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4718 = 6'h2e == _T_596 ? _T_66 : _GEN_4717; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4719 = 6'h2f == _T_596 ? _T_67 : _GEN_4718; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4720 = 6'h30 == _T_596 ? _T_68 : _GEN_4719; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4721 = 6'h31 == _T_596 ? _T_69 : _GEN_4720; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4722 = 6'h32 == _T_596 ? _T_70 : _GEN_4721; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4723 = 6'h33 == _T_596 ? _T_71 : _GEN_4722; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4724 = 6'h34 == _T_596 ? _T_72 : _GEN_4723; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4725 = 6'h35 == _T_596 ? _T_73 : _GEN_4724; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4726 = 6'h36 == _T_596 ? _T_74 : _GEN_4725; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4727 = 6'h37 == _T_596 ? _T_75 : _GEN_4726; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4728 = 6'h38 == _T_596 ? _T_76 : _GEN_4727; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4729 = 6'h39 == _T_596 ? _T_77 : _GEN_4728; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4730 = 6'h3a == _T_596 ? _T_78 : _GEN_4729; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4731 = 6'h3b == _T_596 ? _T_79 : _GEN_4730; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4732 = 6'h3c == _T_596 ? _T_80 : _GEN_4731; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4733 = 6'h3d == _T_596 ? _T_81 : _GEN_4732; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4734 = 6'h3e == _T_596 ? _T_82 : _GEN_4733; // @[execute.scala 79:10:@2109.4]
  assign _GEN_4735 = 6'h3f == _T_596 ? _T_83 : _GEN_4734; // @[execute.scala 79:10:@2109.4]
  assign _T_598 = _T_588 ? _GEN_4671 : _GEN_4735; // @[execute.scala 79:10:@2109.4]
  assign _T_600 = io_amount < 6'h1b; // @[execute.scala 79:15:@2110.4]
  assign _T_602 = io_amount - 6'h1b; // @[execute.scala 79:37:@2111.4]
  assign _T_603 = $unsigned(_T_602); // @[execute.scala 79:37:@2112.4]
  assign _T_604 = _T_603[5:0]; // @[execute.scala 79:37:@2113.4]
  assign _T_607 = 6'h25 + io_amount; // @[execute.scala 79:60:@2114.4]
  assign _T_608 = 6'h25 + io_amount; // @[execute.scala 79:60:@2115.4]
  assign _GEN_4737 = 6'h1 == _T_604 ? _T_21 : _T_20; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4738 = 6'h2 == _T_604 ? _T_22 : _GEN_4737; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4739 = 6'h3 == _T_604 ? _T_23 : _GEN_4738; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4740 = 6'h4 == _T_604 ? _T_24 : _GEN_4739; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4741 = 6'h5 == _T_604 ? _T_25 : _GEN_4740; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4742 = 6'h6 == _T_604 ? _T_26 : _GEN_4741; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4743 = 6'h7 == _T_604 ? _T_27 : _GEN_4742; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4744 = 6'h8 == _T_604 ? _T_28 : _GEN_4743; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4745 = 6'h9 == _T_604 ? _T_29 : _GEN_4744; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4746 = 6'ha == _T_604 ? _T_30 : _GEN_4745; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4747 = 6'hb == _T_604 ? _T_31 : _GEN_4746; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4748 = 6'hc == _T_604 ? _T_32 : _GEN_4747; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4749 = 6'hd == _T_604 ? _T_33 : _GEN_4748; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4750 = 6'he == _T_604 ? _T_34 : _GEN_4749; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4751 = 6'hf == _T_604 ? _T_35 : _GEN_4750; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4752 = 6'h10 == _T_604 ? _T_36 : _GEN_4751; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4753 = 6'h11 == _T_604 ? _T_37 : _GEN_4752; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4754 = 6'h12 == _T_604 ? _T_38 : _GEN_4753; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4755 = 6'h13 == _T_604 ? _T_39 : _GEN_4754; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4756 = 6'h14 == _T_604 ? _T_40 : _GEN_4755; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4757 = 6'h15 == _T_604 ? _T_41 : _GEN_4756; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4758 = 6'h16 == _T_604 ? _T_42 : _GEN_4757; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4759 = 6'h17 == _T_604 ? _T_43 : _GEN_4758; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4760 = 6'h18 == _T_604 ? _T_44 : _GEN_4759; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4761 = 6'h19 == _T_604 ? _T_45 : _GEN_4760; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4762 = 6'h1a == _T_604 ? _T_46 : _GEN_4761; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4763 = 6'h1b == _T_604 ? _T_47 : _GEN_4762; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4764 = 6'h1c == _T_604 ? _T_48 : _GEN_4763; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4765 = 6'h1d == _T_604 ? _T_49 : _GEN_4764; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4766 = 6'h1e == _T_604 ? _T_50 : _GEN_4765; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4767 = 6'h1f == _T_604 ? _T_51 : _GEN_4766; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4768 = 6'h20 == _T_604 ? _T_52 : _GEN_4767; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4769 = 6'h21 == _T_604 ? _T_53 : _GEN_4768; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4770 = 6'h22 == _T_604 ? _T_54 : _GEN_4769; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4771 = 6'h23 == _T_604 ? _T_55 : _GEN_4770; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4772 = 6'h24 == _T_604 ? _T_56 : _GEN_4771; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4773 = 6'h25 == _T_604 ? _T_57 : _GEN_4772; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4774 = 6'h26 == _T_604 ? _T_58 : _GEN_4773; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4775 = 6'h27 == _T_604 ? _T_59 : _GEN_4774; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4776 = 6'h28 == _T_604 ? _T_60 : _GEN_4775; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4777 = 6'h29 == _T_604 ? _T_61 : _GEN_4776; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4778 = 6'h2a == _T_604 ? _T_62 : _GEN_4777; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4779 = 6'h2b == _T_604 ? _T_63 : _GEN_4778; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4780 = 6'h2c == _T_604 ? _T_64 : _GEN_4779; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4781 = 6'h2d == _T_604 ? _T_65 : _GEN_4780; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4782 = 6'h2e == _T_604 ? _T_66 : _GEN_4781; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4783 = 6'h2f == _T_604 ? _T_67 : _GEN_4782; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4784 = 6'h30 == _T_604 ? _T_68 : _GEN_4783; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4785 = 6'h31 == _T_604 ? _T_69 : _GEN_4784; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4786 = 6'h32 == _T_604 ? _T_70 : _GEN_4785; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4787 = 6'h33 == _T_604 ? _T_71 : _GEN_4786; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4788 = 6'h34 == _T_604 ? _T_72 : _GEN_4787; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4789 = 6'h35 == _T_604 ? _T_73 : _GEN_4788; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4790 = 6'h36 == _T_604 ? _T_74 : _GEN_4789; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4791 = 6'h37 == _T_604 ? _T_75 : _GEN_4790; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4792 = 6'h38 == _T_604 ? _T_76 : _GEN_4791; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4793 = 6'h39 == _T_604 ? _T_77 : _GEN_4792; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4794 = 6'h3a == _T_604 ? _T_78 : _GEN_4793; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4795 = 6'h3b == _T_604 ? _T_79 : _GEN_4794; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4796 = 6'h3c == _T_604 ? _T_80 : _GEN_4795; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4797 = 6'h3d == _T_604 ? _T_81 : _GEN_4796; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4798 = 6'h3e == _T_604 ? _T_82 : _GEN_4797; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4799 = 6'h3f == _T_604 ? _T_83 : _GEN_4798; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4801 = 6'h1 == _T_608 ? _T_21 : _T_20; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4802 = 6'h2 == _T_608 ? _T_22 : _GEN_4801; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4803 = 6'h3 == _T_608 ? _T_23 : _GEN_4802; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4804 = 6'h4 == _T_608 ? _T_24 : _GEN_4803; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4805 = 6'h5 == _T_608 ? _T_25 : _GEN_4804; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4806 = 6'h6 == _T_608 ? _T_26 : _GEN_4805; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4807 = 6'h7 == _T_608 ? _T_27 : _GEN_4806; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4808 = 6'h8 == _T_608 ? _T_28 : _GEN_4807; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4809 = 6'h9 == _T_608 ? _T_29 : _GEN_4808; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4810 = 6'ha == _T_608 ? _T_30 : _GEN_4809; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4811 = 6'hb == _T_608 ? _T_31 : _GEN_4810; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4812 = 6'hc == _T_608 ? _T_32 : _GEN_4811; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4813 = 6'hd == _T_608 ? _T_33 : _GEN_4812; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4814 = 6'he == _T_608 ? _T_34 : _GEN_4813; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4815 = 6'hf == _T_608 ? _T_35 : _GEN_4814; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4816 = 6'h10 == _T_608 ? _T_36 : _GEN_4815; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4817 = 6'h11 == _T_608 ? _T_37 : _GEN_4816; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4818 = 6'h12 == _T_608 ? _T_38 : _GEN_4817; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4819 = 6'h13 == _T_608 ? _T_39 : _GEN_4818; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4820 = 6'h14 == _T_608 ? _T_40 : _GEN_4819; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4821 = 6'h15 == _T_608 ? _T_41 : _GEN_4820; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4822 = 6'h16 == _T_608 ? _T_42 : _GEN_4821; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4823 = 6'h17 == _T_608 ? _T_43 : _GEN_4822; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4824 = 6'h18 == _T_608 ? _T_44 : _GEN_4823; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4825 = 6'h19 == _T_608 ? _T_45 : _GEN_4824; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4826 = 6'h1a == _T_608 ? _T_46 : _GEN_4825; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4827 = 6'h1b == _T_608 ? _T_47 : _GEN_4826; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4828 = 6'h1c == _T_608 ? _T_48 : _GEN_4827; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4829 = 6'h1d == _T_608 ? _T_49 : _GEN_4828; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4830 = 6'h1e == _T_608 ? _T_50 : _GEN_4829; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4831 = 6'h1f == _T_608 ? _T_51 : _GEN_4830; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4832 = 6'h20 == _T_608 ? _T_52 : _GEN_4831; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4833 = 6'h21 == _T_608 ? _T_53 : _GEN_4832; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4834 = 6'h22 == _T_608 ? _T_54 : _GEN_4833; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4835 = 6'h23 == _T_608 ? _T_55 : _GEN_4834; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4836 = 6'h24 == _T_608 ? _T_56 : _GEN_4835; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4837 = 6'h25 == _T_608 ? _T_57 : _GEN_4836; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4838 = 6'h26 == _T_608 ? _T_58 : _GEN_4837; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4839 = 6'h27 == _T_608 ? _T_59 : _GEN_4838; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4840 = 6'h28 == _T_608 ? _T_60 : _GEN_4839; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4841 = 6'h29 == _T_608 ? _T_61 : _GEN_4840; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4842 = 6'h2a == _T_608 ? _T_62 : _GEN_4841; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4843 = 6'h2b == _T_608 ? _T_63 : _GEN_4842; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4844 = 6'h2c == _T_608 ? _T_64 : _GEN_4843; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4845 = 6'h2d == _T_608 ? _T_65 : _GEN_4844; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4846 = 6'h2e == _T_608 ? _T_66 : _GEN_4845; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4847 = 6'h2f == _T_608 ? _T_67 : _GEN_4846; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4848 = 6'h30 == _T_608 ? _T_68 : _GEN_4847; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4849 = 6'h31 == _T_608 ? _T_69 : _GEN_4848; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4850 = 6'h32 == _T_608 ? _T_70 : _GEN_4849; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4851 = 6'h33 == _T_608 ? _T_71 : _GEN_4850; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4852 = 6'h34 == _T_608 ? _T_72 : _GEN_4851; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4853 = 6'h35 == _T_608 ? _T_73 : _GEN_4852; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4854 = 6'h36 == _T_608 ? _T_74 : _GEN_4853; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4855 = 6'h37 == _T_608 ? _T_75 : _GEN_4854; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4856 = 6'h38 == _T_608 ? _T_76 : _GEN_4855; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4857 = 6'h39 == _T_608 ? _T_77 : _GEN_4856; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4858 = 6'h3a == _T_608 ? _T_78 : _GEN_4857; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4859 = 6'h3b == _T_608 ? _T_79 : _GEN_4858; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4860 = 6'h3c == _T_608 ? _T_80 : _GEN_4859; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4861 = 6'h3d == _T_608 ? _T_81 : _GEN_4860; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4862 = 6'h3e == _T_608 ? _T_82 : _GEN_4861; // @[execute.scala 79:10:@2116.4]
  assign _GEN_4863 = 6'h3f == _T_608 ? _T_83 : _GEN_4862; // @[execute.scala 79:10:@2116.4]
  assign _T_610 = _T_600 ? _GEN_4799 : _GEN_4863; // @[execute.scala 79:10:@2116.4]
  assign _T_612 = io_amount < 6'h1a; // @[execute.scala 79:15:@2117.4]
  assign _T_614 = io_amount - 6'h1a; // @[execute.scala 79:37:@2118.4]
  assign _T_615 = $unsigned(_T_614); // @[execute.scala 79:37:@2119.4]
  assign _T_616 = _T_615[5:0]; // @[execute.scala 79:37:@2120.4]
  assign _T_619 = 6'h26 + io_amount; // @[execute.scala 79:60:@2121.4]
  assign _T_620 = 6'h26 + io_amount; // @[execute.scala 79:60:@2122.4]
  assign _GEN_4865 = 6'h1 == _T_616 ? _T_21 : _T_20; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4866 = 6'h2 == _T_616 ? _T_22 : _GEN_4865; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4867 = 6'h3 == _T_616 ? _T_23 : _GEN_4866; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4868 = 6'h4 == _T_616 ? _T_24 : _GEN_4867; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4869 = 6'h5 == _T_616 ? _T_25 : _GEN_4868; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4870 = 6'h6 == _T_616 ? _T_26 : _GEN_4869; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4871 = 6'h7 == _T_616 ? _T_27 : _GEN_4870; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4872 = 6'h8 == _T_616 ? _T_28 : _GEN_4871; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4873 = 6'h9 == _T_616 ? _T_29 : _GEN_4872; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4874 = 6'ha == _T_616 ? _T_30 : _GEN_4873; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4875 = 6'hb == _T_616 ? _T_31 : _GEN_4874; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4876 = 6'hc == _T_616 ? _T_32 : _GEN_4875; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4877 = 6'hd == _T_616 ? _T_33 : _GEN_4876; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4878 = 6'he == _T_616 ? _T_34 : _GEN_4877; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4879 = 6'hf == _T_616 ? _T_35 : _GEN_4878; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4880 = 6'h10 == _T_616 ? _T_36 : _GEN_4879; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4881 = 6'h11 == _T_616 ? _T_37 : _GEN_4880; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4882 = 6'h12 == _T_616 ? _T_38 : _GEN_4881; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4883 = 6'h13 == _T_616 ? _T_39 : _GEN_4882; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4884 = 6'h14 == _T_616 ? _T_40 : _GEN_4883; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4885 = 6'h15 == _T_616 ? _T_41 : _GEN_4884; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4886 = 6'h16 == _T_616 ? _T_42 : _GEN_4885; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4887 = 6'h17 == _T_616 ? _T_43 : _GEN_4886; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4888 = 6'h18 == _T_616 ? _T_44 : _GEN_4887; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4889 = 6'h19 == _T_616 ? _T_45 : _GEN_4888; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4890 = 6'h1a == _T_616 ? _T_46 : _GEN_4889; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4891 = 6'h1b == _T_616 ? _T_47 : _GEN_4890; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4892 = 6'h1c == _T_616 ? _T_48 : _GEN_4891; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4893 = 6'h1d == _T_616 ? _T_49 : _GEN_4892; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4894 = 6'h1e == _T_616 ? _T_50 : _GEN_4893; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4895 = 6'h1f == _T_616 ? _T_51 : _GEN_4894; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4896 = 6'h20 == _T_616 ? _T_52 : _GEN_4895; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4897 = 6'h21 == _T_616 ? _T_53 : _GEN_4896; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4898 = 6'h22 == _T_616 ? _T_54 : _GEN_4897; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4899 = 6'h23 == _T_616 ? _T_55 : _GEN_4898; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4900 = 6'h24 == _T_616 ? _T_56 : _GEN_4899; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4901 = 6'h25 == _T_616 ? _T_57 : _GEN_4900; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4902 = 6'h26 == _T_616 ? _T_58 : _GEN_4901; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4903 = 6'h27 == _T_616 ? _T_59 : _GEN_4902; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4904 = 6'h28 == _T_616 ? _T_60 : _GEN_4903; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4905 = 6'h29 == _T_616 ? _T_61 : _GEN_4904; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4906 = 6'h2a == _T_616 ? _T_62 : _GEN_4905; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4907 = 6'h2b == _T_616 ? _T_63 : _GEN_4906; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4908 = 6'h2c == _T_616 ? _T_64 : _GEN_4907; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4909 = 6'h2d == _T_616 ? _T_65 : _GEN_4908; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4910 = 6'h2e == _T_616 ? _T_66 : _GEN_4909; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4911 = 6'h2f == _T_616 ? _T_67 : _GEN_4910; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4912 = 6'h30 == _T_616 ? _T_68 : _GEN_4911; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4913 = 6'h31 == _T_616 ? _T_69 : _GEN_4912; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4914 = 6'h32 == _T_616 ? _T_70 : _GEN_4913; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4915 = 6'h33 == _T_616 ? _T_71 : _GEN_4914; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4916 = 6'h34 == _T_616 ? _T_72 : _GEN_4915; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4917 = 6'h35 == _T_616 ? _T_73 : _GEN_4916; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4918 = 6'h36 == _T_616 ? _T_74 : _GEN_4917; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4919 = 6'h37 == _T_616 ? _T_75 : _GEN_4918; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4920 = 6'h38 == _T_616 ? _T_76 : _GEN_4919; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4921 = 6'h39 == _T_616 ? _T_77 : _GEN_4920; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4922 = 6'h3a == _T_616 ? _T_78 : _GEN_4921; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4923 = 6'h3b == _T_616 ? _T_79 : _GEN_4922; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4924 = 6'h3c == _T_616 ? _T_80 : _GEN_4923; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4925 = 6'h3d == _T_616 ? _T_81 : _GEN_4924; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4926 = 6'h3e == _T_616 ? _T_82 : _GEN_4925; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4927 = 6'h3f == _T_616 ? _T_83 : _GEN_4926; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4929 = 6'h1 == _T_620 ? _T_21 : _T_20; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4930 = 6'h2 == _T_620 ? _T_22 : _GEN_4929; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4931 = 6'h3 == _T_620 ? _T_23 : _GEN_4930; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4932 = 6'h4 == _T_620 ? _T_24 : _GEN_4931; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4933 = 6'h5 == _T_620 ? _T_25 : _GEN_4932; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4934 = 6'h6 == _T_620 ? _T_26 : _GEN_4933; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4935 = 6'h7 == _T_620 ? _T_27 : _GEN_4934; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4936 = 6'h8 == _T_620 ? _T_28 : _GEN_4935; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4937 = 6'h9 == _T_620 ? _T_29 : _GEN_4936; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4938 = 6'ha == _T_620 ? _T_30 : _GEN_4937; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4939 = 6'hb == _T_620 ? _T_31 : _GEN_4938; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4940 = 6'hc == _T_620 ? _T_32 : _GEN_4939; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4941 = 6'hd == _T_620 ? _T_33 : _GEN_4940; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4942 = 6'he == _T_620 ? _T_34 : _GEN_4941; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4943 = 6'hf == _T_620 ? _T_35 : _GEN_4942; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4944 = 6'h10 == _T_620 ? _T_36 : _GEN_4943; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4945 = 6'h11 == _T_620 ? _T_37 : _GEN_4944; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4946 = 6'h12 == _T_620 ? _T_38 : _GEN_4945; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4947 = 6'h13 == _T_620 ? _T_39 : _GEN_4946; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4948 = 6'h14 == _T_620 ? _T_40 : _GEN_4947; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4949 = 6'h15 == _T_620 ? _T_41 : _GEN_4948; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4950 = 6'h16 == _T_620 ? _T_42 : _GEN_4949; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4951 = 6'h17 == _T_620 ? _T_43 : _GEN_4950; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4952 = 6'h18 == _T_620 ? _T_44 : _GEN_4951; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4953 = 6'h19 == _T_620 ? _T_45 : _GEN_4952; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4954 = 6'h1a == _T_620 ? _T_46 : _GEN_4953; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4955 = 6'h1b == _T_620 ? _T_47 : _GEN_4954; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4956 = 6'h1c == _T_620 ? _T_48 : _GEN_4955; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4957 = 6'h1d == _T_620 ? _T_49 : _GEN_4956; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4958 = 6'h1e == _T_620 ? _T_50 : _GEN_4957; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4959 = 6'h1f == _T_620 ? _T_51 : _GEN_4958; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4960 = 6'h20 == _T_620 ? _T_52 : _GEN_4959; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4961 = 6'h21 == _T_620 ? _T_53 : _GEN_4960; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4962 = 6'h22 == _T_620 ? _T_54 : _GEN_4961; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4963 = 6'h23 == _T_620 ? _T_55 : _GEN_4962; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4964 = 6'h24 == _T_620 ? _T_56 : _GEN_4963; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4965 = 6'h25 == _T_620 ? _T_57 : _GEN_4964; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4966 = 6'h26 == _T_620 ? _T_58 : _GEN_4965; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4967 = 6'h27 == _T_620 ? _T_59 : _GEN_4966; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4968 = 6'h28 == _T_620 ? _T_60 : _GEN_4967; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4969 = 6'h29 == _T_620 ? _T_61 : _GEN_4968; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4970 = 6'h2a == _T_620 ? _T_62 : _GEN_4969; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4971 = 6'h2b == _T_620 ? _T_63 : _GEN_4970; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4972 = 6'h2c == _T_620 ? _T_64 : _GEN_4971; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4973 = 6'h2d == _T_620 ? _T_65 : _GEN_4972; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4974 = 6'h2e == _T_620 ? _T_66 : _GEN_4973; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4975 = 6'h2f == _T_620 ? _T_67 : _GEN_4974; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4976 = 6'h30 == _T_620 ? _T_68 : _GEN_4975; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4977 = 6'h31 == _T_620 ? _T_69 : _GEN_4976; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4978 = 6'h32 == _T_620 ? _T_70 : _GEN_4977; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4979 = 6'h33 == _T_620 ? _T_71 : _GEN_4978; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4980 = 6'h34 == _T_620 ? _T_72 : _GEN_4979; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4981 = 6'h35 == _T_620 ? _T_73 : _GEN_4980; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4982 = 6'h36 == _T_620 ? _T_74 : _GEN_4981; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4983 = 6'h37 == _T_620 ? _T_75 : _GEN_4982; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4984 = 6'h38 == _T_620 ? _T_76 : _GEN_4983; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4985 = 6'h39 == _T_620 ? _T_77 : _GEN_4984; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4986 = 6'h3a == _T_620 ? _T_78 : _GEN_4985; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4987 = 6'h3b == _T_620 ? _T_79 : _GEN_4986; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4988 = 6'h3c == _T_620 ? _T_80 : _GEN_4987; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4989 = 6'h3d == _T_620 ? _T_81 : _GEN_4988; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4990 = 6'h3e == _T_620 ? _T_82 : _GEN_4989; // @[execute.scala 79:10:@2123.4]
  assign _GEN_4991 = 6'h3f == _T_620 ? _T_83 : _GEN_4990; // @[execute.scala 79:10:@2123.4]
  assign _T_622 = _T_612 ? _GEN_4927 : _GEN_4991; // @[execute.scala 79:10:@2123.4]
  assign _T_624 = io_amount < 6'h19; // @[execute.scala 79:15:@2124.4]
  assign _T_626 = io_amount - 6'h19; // @[execute.scala 79:37:@2125.4]
  assign _T_627 = $unsigned(_T_626); // @[execute.scala 79:37:@2126.4]
  assign _T_628 = _T_627[5:0]; // @[execute.scala 79:37:@2127.4]
  assign _T_631 = 6'h27 + io_amount; // @[execute.scala 79:60:@2128.4]
  assign _T_632 = 6'h27 + io_amount; // @[execute.scala 79:60:@2129.4]
  assign _GEN_4993 = 6'h1 == _T_628 ? _T_21 : _T_20; // @[execute.scala 79:10:@2130.4]
  assign _GEN_4994 = 6'h2 == _T_628 ? _T_22 : _GEN_4993; // @[execute.scala 79:10:@2130.4]
  assign _GEN_4995 = 6'h3 == _T_628 ? _T_23 : _GEN_4994; // @[execute.scala 79:10:@2130.4]
  assign _GEN_4996 = 6'h4 == _T_628 ? _T_24 : _GEN_4995; // @[execute.scala 79:10:@2130.4]
  assign _GEN_4997 = 6'h5 == _T_628 ? _T_25 : _GEN_4996; // @[execute.scala 79:10:@2130.4]
  assign _GEN_4998 = 6'h6 == _T_628 ? _T_26 : _GEN_4997; // @[execute.scala 79:10:@2130.4]
  assign _GEN_4999 = 6'h7 == _T_628 ? _T_27 : _GEN_4998; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5000 = 6'h8 == _T_628 ? _T_28 : _GEN_4999; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5001 = 6'h9 == _T_628 ? _T_29 : _GEN_5000; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5002 = 6'ha == _T_628 ? _T_30 : _GEN_5001; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5003 = 6'hb == _T_628 ? _T_31 : _GEN_5002; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5004 = 6'hc == _T_628 ? _T_32 : _GEN_5003; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5005 = 6'hd == _T_628 ? _T_33 : _GEN_5004; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5006 = 6'he == _T_628 ? _T_34 : _GEN_5005; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5007 = 6'hf == _T_628 ? _T_35 : _GEN_5006; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5008 = 6'h10 == _T_628 ? _T_36 : _GEN_5007; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5009 = 6'h11 == _T_628 ? _T_37 : _GEN_5008; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5010 = 6'h12 == _T_628 ? _T_38 : _GEN_5009; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5011 = 6'h13 == _T_628 ? _T_39 : _GEN_5010; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5012 = 6'h14 == _T_628 ? _T_40 : _GEN_5011; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5013 = 6'h15 == _T_628 ? _T_41 : _GEN_5012; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5014 = 6'h16 == _T_628 ? _T_42 : _GEN_5013; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5015 = 6'h17 == _T_628 ? _T_43 : _GEN_5014; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5016 = 6'h18 == _T_628 ? _T_44 : _GEN_5015; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5017 = 6'h19 == _T_628 ? _T_45 : _GEN_5016; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5018 = 6'h1a == _T_628 ? _T_46 : _GEN_5017; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5019 = 6'h1b == _T_628 ? _T_47 : _GEN_5018; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5020 = 6'h1c == _T_628 ? _T_48 : _GEN_5019; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5021 = 6'h1d == _T_628 ? _T_49 : _GEN_5020; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5022 = 6'h1e == _T_628 ? _T_50 : _GEN_5021; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5023 = 6'h1f == _T_628 ? _T_51 : _GEN_5022; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5024 = 6'h20 == _T_628 ? _T_52 : _GEN_5023; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5025 = 6'h21 == _T_628 ? _T_53 : _GEN_5024; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5026 = 6'h22 == _T_628 ? _T_54 : _GEN_5025; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5027 = 6'h23 == _T_628 ? _T_55 : _GEN_5026; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5028 = 6'h24 == _T_628 ? _T_56 : _GEN_5027; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5029 = 6'h25 == _T_628 ? _T_57 : _GEN_5028; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5030 = 6'h26 == _T_628 ? _T_58 : _GEN_5029; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5031 = 6'h27 == _T_628 ? _T_59 : _GEN_5030; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5032 = 6'h28 == _T_628 ? _T_60 : _GEN_5031; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5033 = 6'h29 == _T_628 ? _T_61 : _GEN_5032; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5034 = 6'h2a == _T_628 ? _T_62 : _GEN_5033; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5035 = 6'h2b == _T_628 ? _T_63 : _GEN_5034; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5036 = 6'h2c == _T_628 ? _T_64 : _GEN_5035; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5037 = 6'h2d == _T_628 ? _T_65 : _GEN_5036; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5038 = 6'h2e == _T_628 ? _T_66 : _GEN_5037; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5039 = 6'h2f == _T_628 ? _T_67 : _GEN_5038; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5040 = 6'h30 == _T_628 ? _T_68 : _GEN_5039; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5041 = 6'h31 == _T_628 ? _T_69 : _GEN_5040; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5042 = 6'h32 == _T_628 ? _T_70 : _GEN_5041; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5043 = 6'h33 == _T_628 ? _T_71 : _GEN_5042; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5044 = 6'h34 == _T_628 ? _T_72 : _GEN_5043; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5045 = 6'h35 == _T_628 ? _T_73 : _GEN_5044; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5046 = 6'h36 == _T_628 ? _T_74 : _GEN_5045; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5047 = 6'h37 == _T_628 ? _T_75 : _GEN_5046; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5048 = 6'h38 == _T_628 ? _T_76 : _GEN_5047; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5049 = 6'h39 == _T_628 ? _T_77 : _GEN_5048; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5050 = 6'h3a == _T_628 ? _T_78 : _GEN_5049; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5051 = 6'h3b == _T_628 ? _T_79 : _GEN_5050; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5052 = 6'h3c == _T_628 ? _T_80 : _GEN_5051; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5053 = 6'h3d == _T_628 ? _T_81 : _GEN_5052; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5054 = 6'h3e == _T_628 ? _T_82 : _GEN_5053; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5055 = 6'h3f == _T_628 ? _T_83 : _GEN_5054; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5057 = 6'h1 == _T_632 ? _T_21 : _T_20; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5058 = 6'h2 == _T_632 ? _T_22 : _GEN_5057; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5059 = 6'h3 == _T_632 ? _T_23 : _GEN_5058; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5060 = 6'h4 == _T_632 ? _T_24 : _GEN_5059; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5061 = 6'h5 == _T_632 ? _T_25 : _GEN_5060; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5062 = 6'h6 == _T_632 ? _T_26 : _GEN_5061; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5063 = 6'h7 == _T_632 ? _T_27 : _GEN_5062; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5064 = 6'h8 == _T_632 ? _T_28 : _GEN_5063; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5065 = 6'h9 == _T_632 ? _T_29 : _GEN_5064; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5066 = 6'ha == _T_632 ? _T_30 : _GEN_5065; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5067 = 6'hb == _T_632 ? _T_31 : _GEN_5066; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5068 = 6'hc == _T_632 ? _T_32 : _GEN_5067; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5069 = 6'hd == _T_632 ? _T_33 : _GEN_5068; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5070 = 6'he == _T_632 ? _T_34 : _GEN_5069; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5071 = 6'hf == _T_632 ? _T_35 : _GEN_5070; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5072 = 6'h10 == _T_632 ? _T_36 : _GEN_5071; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5073 = 6'h11 == _T_632 ? _T_37 : _GEN_5072; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5074 = 6'h12 == _T_632 ? _T_38 : _GEN_5073; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5075 = 6'h13 == _T_632 ? _T_39 : _GEN_5074; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5076 = 6'h14 == _T_632 ? _T_40 : _GEN_5075; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5077 = 6'h15 == _T_632 ? _T_41 : _GEN_5076; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5078 = 6'h16 == _T_632 ? _T_42 : _GEN_5077; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5079 = 6'h17 == _T_632 ? _T_43 : _GEN_5078; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5080 = 6'h18 == _T_632 ? _T_44 : _GEN_5079; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5081 = 6'h19 == _T_632 ? _T_45 : _GEN_5080; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5082 = 6'h1a == _T_632 ? _T_46 : _GEN_5081; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5083 = 6'h1b == _T_632 ? _T_47 : _GEN_5082; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5084 = 6'h1c == _T_632 ? _T_48 : _GEN_5083; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5085 = 6'h1d == _T_632 ? _T_49 : _GEN_5084; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5086 = 6'h1e == _T_632 ? _T_50 : _GEN_5085; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5087 = 6'h1f == _T_632 ? _T_51 : _GEN_5086; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5088 = 6'h20 == _T_632 ? _T_52 : _GEN_5087; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5089 = 6'h21 == _T_632 ? _T_53 : _GEN_5088; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5090 = 6'h22 == _T_632 ? _T_54 : _GEN_5089; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5091 = 6'h23 == _T_632 ? _T_55 : _GEN_5090; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5092 = 6'h24 == _T_632 ? _T_56 : _GEN_5091; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5093 = 6'h25 == _T_632 ? _T_57 : _GEN_5092; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5094 = 6'h26 == _T_632 ? _T_58 : _GEN_5093; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5095 = 6'h27 == _T_632 ? _T_59 : _GEN_5094; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5096 = 6'h28 == _T_632 ? _T_60 : _GEN_5095; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5097 = 6'h29 == _T_632 ? _T_61 : _GEN_5096; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5098 = 6'h2a == _T_632 ? _T_62 : _GEN_5097; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5099 = 6'h2b == _T_632 ? _T_63 : _GEN_5098; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5100 = 6'h2c == _T_632 ? _T_64 : _GEN_5099; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5101 = 6'h2d == _T_632 ? _T_65 : _GEN_5100; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5102 = 6'h2e == _T_632 ? _T_66 : _GEN_5101; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5103 = 6'h2f == _T_632 ? _T_67 : _GEN_5102; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5104 = 6'h30 == _T_632 ? _T_68 : _GEN_5103; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5105 = 6'h31 == _T_632 ? _T_69 : _GEN_5104; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5106 = 6'h32 == _T_632 ? _T_70 : _GEN_5105; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5107 = 6'h33 == _T_632 ? _T_71 : _GEN_5106; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5108 = 6'h34 == _T_632 ? _T_72 : _GEN_5107; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5109 = 6'h35 == _T_632 ? _T_73 : _GEN_5108; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5110 = 6'h36 == _T_632 ? _T_74 : _GEN_5109; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5111 = 6'h37 == _T_632 ? _T_75 : _GEN_5110; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5112 = 6'h38 == _T_632 ? _T_76 : _GEN_5111; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5113 = 6'h39 == _T_632 ? _T_77 : _GEN_5112; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5114 = 6'h3a == _T_632 ? _T_78 : _GEN_5113; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5115 = 6'h3b == _T_632 ? _T_79 : _GEN_5114; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5116 = 6'h3c == _T_632 ? _T_80 : _GEN_5115; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5117 = 6'h3d == _T_632 ? _T_81 : _GEN_5116; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5118 = 6'h3e == _T_632 ? _T_82 : _GEN_5117; // @[execute.scala 79:10:@2130.4]
  assign _GEN_5119 = 6'h3f == _T_632 ? _T_83 : _GEN_5118; // @[execute.scala 79:10:@2130.4]
  assign _T_634 = _T_624 ? _GEN_5055 : _GEN_5119; // @[execute.scala 79:10:@2130.4]
  assign _T_636 = io_amount < 6'h18; // @[execute.scala 79:15:@2131.4]
  assign _T_638 = io_amount - 6'h18; // @[execute.scala 79:37:@2132.4]
  assign _T_639 = $unsigned(_T_638); // @[execute.scala 79:37:@2133.4]
  assign _T_640 = _T_639[5:0]; // @[execute.scala 79:37:@2134.4]
  assign _T_643 = 6'h28 + io_amount; // @[execute.scala 79:60:@2135.4]
  assign _T_644 = 6'h28 + io_amount; // @[execute.scala 79:60:@2136.4]
  assign _GEN_5121 = 6'h1 == _T_640 ? _T_21 : _T_20; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5122 = 6'h2 == _T_640 ? _T_22 : _GEN_5121; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5123 = 6'h3 == _T_640 ? _T_23 : _GEN_5122; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5124 = 6'h4 == _T_640 ? _T_24 : _GEN_5123; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5125 = 6'h5 == _T_640 ? _T_25 : _GEN_5124; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5126 = 6'h6 == _T_640 ? _T_26 : _GEN_5125; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5127 = 6'h7 == _T_640 ? _T_27 : _GEN_5126; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5128 = 6'h8 == _T_640 ? _T_28 : _GEN_5127; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5129 = 6'h9 == _T_640 ? _T_29 : _GEN_5128; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5130 = 6'ha == _T_640 ? _T_30 : _GEN_5129; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5131 = 6'hb == _T_640 ? _T_31 : _GEN_5130; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5132 = 6'hc == _T_640 ? _T_32 : _GEN_5131; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5133 = 6'hd == _T_640 ? _T_33 : _GEN_5132; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5134 = 6'he == _T_640 ? _T_34 : _GEN_5133; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5135 = 6'hf == _T_640 ? _T_35 : _GEN_5134; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5136 = 6'h10 == _T_640 ? _T_36 : _GEN_5135; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5137 = 6'h11 == _T_640 ? _T_37 : _GEN_5136; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5138 = 6'h12 == _T_640 ? _T_38 : _GEN_5137; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5139 = 6'h13 == _T_640 ? _T_39 : _GEN_5138; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5140 = 6'h14 == _T_640 ? _T_40 : _GEN_5139; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5141 = 6'h15 == _T_640 ? _T_41 : _GEN_5140; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5142 = 6'h16 == _T_640 ? _T_42 : _GEN_5141; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5143 = 6'h17 == _T_640 ? _T_43 : _GEN_5142; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5144 = 6'h18 == _T_640 ? _T_44 : _GEN_5143; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5145 = 6'h19 == _T_640 ? _T_45 : _GEN_5144; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5146 = 6'h1a == _T_640 ? _T_46 : _GEN_5145; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5147 = 6'h1b == _T_640 ? _T_47 : _GEN_5146; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5148 = 6'h1c == _T_640 ? _T_48 : _GEN_5147; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5149 = 6'h1d == _T_640 ? _T_49 : _GEN_5148; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5150 = 6'h1e == _T_640 ? _T_50 : _GEN_5149; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5151 = 6'h1f == _T_640 ? _T_51 : _GEN_5150; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5152 = 6'h20 == _T_640 ? _T_52 : _GEN_5151; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5153 = 6'h21 == _T_640 ? _T_53 : _GEN_5152; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5154 = 6'h22 == _T_640 ? _T_54 : _GEN_5153; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5155 = 6'h23 == _T_640 ? _T_55 : _GEN_5154; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5156 = 6'h24 == _T_640 ? _T_56 : _GEN_5155; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5157 = 6'h25 == _T_640 ? _T_57 : _GEN_5156; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5158 = 6'h26 == _T_640 ? _T_58 : _GEN_5157; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5159 = 6'h27 == _T_640 ? _T_59 : _GEN_5158; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5160 = 6'h28 == _T_640 ? _T_60 : _GEN_5159; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5161 = 6'h29 == _T_640 ? _T_61 : _GEN_5160; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5162 = 6'h2a == _T_640 ? _T_62 : _GEN_5161; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5163 = 6'h2b == _T_640 ? _T_63 : _GEN_5162; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5164 = 6'h2c == _T_640 ? _T_64 : _GEN_5163; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5165 = 6'h2d == _T_640 ? _T_65 : _GEN_5164; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5166 = 6'h2e == _T_640 ? _T_66 : _GEN_5165; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5167 = 6'h2f == _T_640 ? _T_67 : _GEN_5166; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5168 = 6'h30 == _T_640 ? _T_68 : _GEN_5167; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5169 = 6'h31 == _T_640 ? _T_69 : _GEN_5168; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5170 = 6'h32 == _T_640 ? _T_70 : _GEN_5169; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5171 = 6'h33 == _T_640 ? _T_71 : _GEN_5170; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5172 = 6'h34 == _T_640 ? _T_72 : _GEN_5171; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5173 = 6'h35 == _T_640 ? _T_73 : _GEN_5172; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5174 = 6'h36 == _T_640 ? _T_74 : _GEN_5173; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5175 = 6'h37 == _T_640 ? _T_75 : _GEN_5174; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5176 = 6'h38 == _T_640 ? _T_76 : _GEN_5175; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5177 = 6'h39 == _T_640 ? _T_77 : _GEN_5176; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5178 = 6'h3a == _T_640 ? _T_78 : _GEN_5177; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5179 = 6'h3b == _T_640 ? _T_79 : _GEN_5178; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5180 = 6'h3c == _T_640 ? _T_80 : _GEN_5179; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5181 = 6'h3d == _T_640 ? _T_81 : _GEN_5180; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5182 = 6'h3e == _T_640 ? _T_82 : _GEN_5181; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5183 = 6'h3f == _T_640 ? _T_83 : _GEN_5182; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5185 = 6'h1 == _T_644 ? _T_21 : _T_20; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5186 = 6'h2 == _T_644 ? _T_22 : _GEN_5185; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5187 = 6'h3 == _T_644 ? _T_23 : _GEN_5186; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5188 = 6'h4 == _T_644 ? _T_24 : _GEN_5187; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5189 = 6'h5 == _T_644 ? _T_25 : _GEN_5188; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5190 = 6'h6 == _T_644 ? _T_26 : _GEN_5189; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5191 = 6'h7 == _T_644 ? _T_27 : _GEN_5190; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5192 = 6'h8 == _T_644 ? _T_28 : _GEN_5191; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5193 = 6'h9 == _T_644 ? _T_29 : _GEN_5192; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5194 = 6'ha == _T_644 ? _T_30 : _GEN_5193; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5195 = 6'hb == _T_644 ? _T_31 : _GEN_5194; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5196 = 6'hc == _T_644 ? _T_32 : _GEN_5195; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5197 = 6'hd == _T_644 ? _T_33 : _GEN_5196; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5198 = 6'he == _T_644 ? _T_34 : _GEN_5197; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5199 = 6'hf == _T_644 ? _T_35 : _GEN_5198; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5200 = 6'h10 == _T_644 ? _T_36 : _GEN_5199; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5201 = 6'h11 == _T_644 ? _T_37 : _GEN_5200; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5202 = 6'h12 == _T_644 ? _T_38 : _GEN_5201; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5203 = 6'h13 == _T_644 ? _T_39 : _GEN_5202; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5204 = 6'h14 == _T_644 ? _T_40 : _GEN_5203; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5205 = 6'h15 == _T_644 ? _T_41 : _GEN_5204; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5206 = 6'h16 == _T_644 ? _T_42 : _GEN_5205; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5207 = 6'h17 == _T_644 ? _T_43 : _GEN_5206; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5208 = 6'h18 == _T_644 ? _T_44 : _GEN_5207; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5209 = 6'h19 == _T_644 ? _T_45 : _GEN_5208; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5210 = 6'h1a == _T_644 ? _T_46 : _GEN_5209; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5211 = 6'h1b == _T_644 ? _T_47 : _GEN_5210; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5212 = 6'h1c == _T_644 ? _T_48 : _GEN_5211; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5213 = 6'h1d == _T_644 ? _T_49 : _GEN_5212; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5214 = 6'h1e == _T_644 ? _T_50 : _GEN_5213; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5215 = 6'h1f == _T_644 ? _T_51 : _GEN_5214; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5216 = 6'h20 == _T_644 ? _T_52 : _GEN_5215; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5217 = 6'h21 == _T_644 ? _T_53 : _GEN_5216; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5218 = 6'h22 == _T_644 ? _T_54 : _GEN_5217; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5219 = 6'h23 == _T_644 ? _T_55 : _GEN_5218; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5220 = 6'h24 == _T_644 ? _T_56 : _GEN_5219; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5221 = 6'h25 == _T_644 ? _T_57 : _GEN_5220; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5222 = 6'h26 == _T_644 ? _T_58 : _GEN_5221; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5223 = 6'h27 == _T_644 ? _T_59 : _GEN_5222; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5224 = 6'h28 == _T_644 ? _T_60 : _GEN_5223; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5225 = 6'h29 == _T_644 ? _T_61 : _GEN_5224; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5226 = 6'h2a == _T_644 ? _T_62 : _GEN_5225; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5227 = 6'h2b == _T_644 ? _T_63 : _GEN_5226; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5228 = 6'h2c == _T_644 ? _T_64 : _GEN_5227; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5229 = 6'h2d == _T_644 ? _T_65 : _GEN_5228; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5230 = 6'h2e == _T_644 ? _T_66 : _GEN_5229; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5231 = 6'h2f == _T_644 ? _T_67 : _GEN_5230; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5232 = 6'h30 == _T_644 ? _T_68 : _GEN_5231; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5233 = 6'h31 == _T_644 ? _T_69 : _GEN_5232; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5234 = 6'h32 == _T_644 ? _T_70 : _GEN_5233; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5235 = 6'h33 == _T_644 ? _T_71 : _GEN_5234; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5236 = 6'h34 == _T_644 ? _T_72 : _GEN_5235; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5237 = 6'h35 == _T_644 ? _T_73 : _GEN_5236; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5238 = 6'h36 == _T_644 ? _T_74 : _GEN_5237; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5239 = 6'h37 == _T_644 ? _T_75 : _GEN_5238; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5240 = 6'h38 == _T_644 ? _T_76 : _GEN_5239; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5241 = 6'h39 == _T_644 ? _T_77 : _GEN_5240; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5242 = 6'h3a == _T_644 ? _T_78 : _GEN_5241; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5243 = 6'h3b == _T_644 ? _T_79 : _GEN_5242; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5244 = 6'h3c == _T_644 ? _T_80 : _GEN_5243; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5245 = 6'h3d == _T_644 ? _T_81 : _GEN_5244; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5246 = 6'h3e == _T_644 ? _T_82 : _GEN_5245; // @[execute.scala 79:10:@2137.4]
  assign _GEN_5247 = 6'h3f == _T_644 ? _T_83 : _GEN_5246; // @[execute.scala 79:10:@2137.4]
  assign _T_646 = _T_636 ? _GEN_5183 : _GEN_5247; // @[execute.scala 79:10:@2137.4]
  assign _T_648 = io_amount < 6'h17; // @[execute.scala 79:15:@2138.4]
  assign _T_650 = io_amount - 6'h17; // @[execute.scala 79:37:@2139.4]
  assign _T_651 = $unsigned(_T_650); // @[execute.scala 79:37:@2140.4]
  assign _T_652 = _T_651[5:0]; // @[execute.scala 79:37:@2141.4]
  assign _T_655 = 6'h29 + io_amount; // @[execute.scala 79:60:@2142.4]
  assign _T_656 = 6'h29 + io_amount; // @[execute.scala 79:60:@2143.4]
  assign _GEN_5249 = 6'h1 == _T_652 ? _T_21 : _T_20; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5250 = 6'h2 == _T_652 ? _T_22 : _GEN_5249; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5251 = 6'h3 == _T_652 ? _T_23 : _GEN_5250; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5252 = 6'h4 == _T_652 ? _T_24 : _GEN_5251; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5253 = 6'h5 == _T_652 ? _T_25 : _GEN_5252; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5254 = 6'h6 == _T_652 ? _T_26 : _GEN_5253; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5255 = 6'h7 == _T_652 ? _T_27 : _GEN_5254; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5256 = 6'h8 == _T_652 ? _T_28 : _GEN_5255; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5257 = 6'h9 == _T_652 ? _T_29 : _GEN_5256; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5258 = 6'ha == _T_652 ? _T_30 : _GEN_5257; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5259 = 6'hb == _T_652 ? _T_31 : _GEN_5258; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5260 = 6'hc == _T_652 ? _T_32 : _GEN_5259; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5261 = 6'hd == _T_652 ? _T_33 : _GEN_5260; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5262 = 6'he == _T_652 ? _T_34 : _GEN_5261; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5263 = 6'hf == _T_652 ? _T_35 : _GEN_5262; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5264 = 6'h10 == _T_652 ? _T_36 : _GEN_5263; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5265 = 6'h11 == _T_652 ? _T_37 : _GEN_5264; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5266 = 6'h12 == _T_652 ? _T_38 : _GEN_5265; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5267 = 6'h13 == _T_652 ? _T_39 : _GEN_5266; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5268 = 6'h14 == _T_652 ? _T_40 : _GEN_5267; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5269 = 6'h15 == _T_652 ? _T_41 : _GEN_5268; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5270 = 6'h16 == _T_652 ? _T_42 : _GEN_5269; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5271 = 6'h17 == _T_652 ? _T_43 : _GEN_5270; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5272 = 6'h18 == _T_652 ? _T_44 : _GEN_5271; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5273 = 6'h19 == _T_652 ? _T_45 : _GEN_5272; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5274 = 6'h1a == _T_652 ? _T_46 : _GEN_5273; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5275 = 6'h1b == _T_652 ? _T_47 : _GEN_5274; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5276 = 6'h1c == _T_652 ? _T_48 : _GEN_5275; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5277 = 6'h1d == _T_652 ? _T_49 : _GEN_5276; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5278 = 6'h1e == _T_652 ? _T_50 : _GEN_5277; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5279 = 6'h1f == _T_652 ? _T_51 : _GEN_5278; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5280 = 6'h20 == _T_652 ? _T_52 : _GEN_5279; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5281 = 6'h21 == _T_652 ? _T_53 : _GEN_5280; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5282 = 6'h22 == _T_652 ? _T_54 : _GEN_5281; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5283 = 6'h23 == _T_652 ? _T_55 : _GEN_5282; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5284 = 6'h24 == _T_652 ? _T_56 : _GEN_5283; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5285 = 6'h25 == _T_652 ? _T_57 : _GEN_5284; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5286 = 6'h26 == _T_652 ? _T_58 : _GEN_5285; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5287 = 6'h27 == _T_652 ? _T_59 : _GEN_5286; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5288 = 6'h28 == _T_652 ? _T_60 : _GEN_5287; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5289 = 6'h29 == _T_652 ? _T_61 : _GEN_5288; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5290 = 6'h2a == _T_652 ? _T_62 : _GEN_5289; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5291 = 6'h2b == _T_652 ? _T_63 : _GEN_5290; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5292 = 6'h2c == _T_652 ? _T_64 : _GEN_5291; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5293 = 6'h2d == _T_652 ? _T_65 : _GEN_5292; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5294 = 6'h2e == _T_652 ? _T_66 : _GEN_5293; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5295 = 6'h2f == _T_652 ? _T_67 : _GEN_5294; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5296 = 6'h30 == _T_652 ? _T_68 : _GEN_5295; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5297 = 6'h31 == _T_652 ? _T_69 : _GEN_5296; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5298 = 6'h32 == _T_652 ? _T_70 : _GEN_5297; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5299 = 6'h33 == _T_652 ? _T_71 : _GEN_5298; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5300 = 6'h34 == _T_652 ? _T_72 : _GEN_5299; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5301 = 6'h35 == _T_652 ? _T_73 : _GEN_5300; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5302 = 6'h36 == _T_652 ? _T_74 : _GEN_5301; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5303 = 6'h37 == _T_652 ? _T_75 : _GEN_5302; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5304 = 6'h38 == _T_652 ? _T_76 : _GEN_5303; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5305 = 6'h39 == _T_652 ? _T_77 : _GEN_5304; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5306 = 6'h3a == _T_652 ? _T_78 : _GEN_5305; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5307 = 6'h3b == _T_652 ? _T_79 : _GEN_5306; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5308 = 6'h3c == _T_652 ? _T_80 : _GEN_5307; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5309 = 6'h3d == _T_652 ? _T_81 : _GEN_5308; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5310 = 6'h3e == _T_652 ? _T_82 : _GEN_5309; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5311 = 6'h3f == _T_652 ? _T_83 : _GEN_5310; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5313 = 6'h1 == _T_656 ? _T_21 : _T_20; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5314 = 6'h2 == _T_656 ? _T_22 : _GEN_5313; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5315 = 6'h3 == _T_656 ? _T_23 : _GEN_5314; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5316 = 6'h4 == _T_656 ? _T_24 : _GEN_5315; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5317 = 6'h5 == _T_656 ? _T_25 : _GEN_5316; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5318 = 6'h6 == _T_656 ? _T_26 : _GEN_5317; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5319 = 6'h7 == _T_656 ? _T_27 : _GEN_5318; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5320 = 6'h8 == _T_656 ? _T_28 : _GEN_5319; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5321 = 6'h9 == _T_656 ? _T_29 : _GEN_5320; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5322 = 6'ha == _T_656 ? _T_30 : _GEN_5321; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5323 = 6'hb == _T_656 ? _T_31 : _GEN_5322; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5324 = 6'hc == _T_656 ? _T_32 : _GEN_5323; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5325 = 6'hd == _T_656 ? _T_33 : _GEN_5324; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5326 = 6'he == _T_656 ? _T_34 : _GEN_5325; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5327 = 6'hf == _T_656 ? _T_35 : _GEN_5326; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5328 = 6'h10 == _T_656 ? _T_36 : _GEN_5327; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5329 = 6'h11 == _T_656 ? _T_37 : _GEN_5328; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5330 = 6'h12 == _T_656 ? _T_38 : _GEN_5329; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5331 = 6'h13 == _T_656 ? _T_39 : _GEN_5330; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5332 = 6'h14 == _T_656 ? _T_40 : _GEN_5331; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5333 = 6'h15 == _T_656 ? _T_41 : _GEN_5332; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5334 = 6'h16 == _T_656 ? _T_42 : _GEN_5333; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5335 = 6'h17 == _T_656 ? _T_43 : _GEN_5334; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5336 = 6'h18 == _T_656 ? _T_44 : _GEN_5335; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5337 = 6'h19 == _T_656 ? _T_45 : _GEN_5336; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5338 = 6'h1a == _T_656 ? _T_46 : _GEN_5337; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5339 = 6'h1b == _T_656 ? _T_47 : _GEN_5338; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5340 = 6'h1c == _T_656 ? _T_48 : _GEN_5339; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5341 = 6'h1d == _T_656 ? _T_49 : _GEN_5340; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5342 = 6'h1e == _T_656 ? _T_50 : _GEN_5341; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5343 = 6'h1f == _T_656 ? _T_51 : _GEN_5342; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5344 = 6'h20 == _T_656 ? _T_52 : _GEN_5343; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5345 = 6'h21 == _T_656 ? _T_53 : _GEN_5344; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5346 = 6'h22 == _T_656 ? _T_54 : _GEN_5345; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5347 = 6'h23 == _T_656 ? _T_55 : _GEN_5346; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5348 = 6'h24 == _T_656 ? _T_56 : _GEN_5347; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5349 = 6'h25 == _T_656 ? _T_57 : _GEN_5348; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5350 = 6'h26 == _T_656 ? _T_58 : _GEN_5349; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5351 = 6'h27 == _T_656 ? _T_59 : _GEN_5350; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5352 = 6'h28 == _T_656 ? _T_60 : _GEN_5351; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5353 = 6'h29 == _T_656 ? _T_61 : _GEN_5352; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5354 = 6'h2a == _T_656 ? _T_62 : _GEN_5353; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5355 = 6'h2b == _T_656 ? _T_63 : _GEN_5354; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5356 = 6'h2c == _T_656 ? _T_64 : _GEN_5355; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5357 = 6'h2d == _T_656 ? _T_65 : _GEN_5356; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5358 = 6'h2e == _T_656 ? _T_66 : _GEN_5357; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5359 = 6'h2f == _T_656 ? _T_67 : _GEN_5358; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5360 = 6'h30 == _T_656 ? _T_68 : _GEN_5359; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5361 = 6'h31 == _T_656 ? _T_69 : _GEN_5360; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5362 = 6'h32 == _T_656 ? _T_70 : _GEN_5361; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5363 = 6'h33 == _T_656 ? _T_71 : _GEN_5362; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5364 = 6'h34 == _T_656 ? _T_72 : _GEN_5363; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5365 = 6'h35 == _T_656 ? _T_73 : _GEN_5364; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5366 = 6'h36 == _T_656 ? _T_74 : _GEN_5365; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5367 = 6'h37 == _T_656 ? _T_75 : _GEN_5366; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5368 = 6'h38 == _T_656 ? _T_76 : _GEN_5367; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5369 = 6'h39 == _T_656 ? _T_77 : _GEN_5368; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5370 = 6'h3a == _T_656 ? _T_78 : _GEN_5369; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5371 = 6'h3b == _T_656 ? _T_79 : _GEN_5370; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5372 = 6'h3c == _T_656 ? _T_80 : _GEN_5371; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5373 = 6'h3d == _T_656 ? _T_81 : _GEN_5372; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5374 = 6'h3e == _T_656 ? _T_82 : _GEN_5373; // @[execute.scala 79:10:@2144.4]
  assign _GEN_5375 = 6'h3f == _T_656 ? _T_83 : _GEN_5374; // @[execute.scala 79:10:@2144.4]
  assign _T_658 = _T_648 ? _GEN_5311 : _GEN_5375; // @[execute.scala 79:10:@2144.4]
  assign _T_660 = io_amount < 6'h16; // @[execute.scala 79:15:@2145.4]
  assign _T_662 = io_amount - 6'h16; // @[execute.scala 79:37:@2146.4]
  assign _T_663 = $unsigned(_T_662); // @[execute.scala 79:37:@2147.4]
  assign _T_664 = _T_663[5:0]; // @[execute.scala 79:37:@2148.4]
  assign _T_667 = 6'h2a + io_amount; // @[execute.scala 79:60:@2149.4]
  assign _T_668 = 6'h2a + io_amount; // @[execute.scala 79:60:@2150.4]
  assign _GEN_5377 = 6'h1 == _T_664 ? _T_21 : _T_20; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5378 = 6'h2 == _T_664 ? _T_22 : _GEN_5377; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5379 = 6'h3 == _T_664 ? _T_23 : _GEN_5378; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5380 = 6'h4 == _T_664 ? _T_24 : _GEN_5379; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5381 = 6'h5 == _T_664 ? _T_25 : _GEN_5380; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5382 = 6'h6 == _T_664 ? _T_26 : _GEN_5381; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5383 = 6'h7 == _T_664 ? _T_27 : _GEN_5382; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5384 = 6'h8 == _T_664 ? _T_28 : _GEN_5383; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5385 = 6'h9 == _T_664 ? _T_29 : _GEN_5384; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5386 = 6'ha == _T_664 ? _T_30 : _GEN_5385; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5387 = 6'hb == _T_664 ? _T_31 : _GEN_5386; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5388 = 6'hc == _T_664 ? _T_32 : _GEN_5387; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5389 = 6'hd == _T_664 ? _T_33 : _GEN_5388; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5390 = 6'he == _T_664 ? _T_34 : _GEN_5389; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5391 = 6'hf == _T_664 ? _T_35 : _GEN_5390; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5392 = 6'h10 == _T_664 ? _T_36 : _GEN_5391; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5393 = 6'h11 == _T_664 ? _T_37 : _GEN_5392; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5394 = 6'h12 == _T_664 ? _T_38 : _GEN_5393; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5395 = 6'h13 == _T_664 ? _T_39 : _GEN_5394; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5396 = 6'h14 == _T_664 ? _T_40 : _GEN_5395; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5397 = 6'h15 == _T_664 ? _T_41 : _GEN_5396; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5398 = 6'h16 == _T_664 ? _T_42 : _GEN_5397; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5399 = 6'h17 == _T_664 ? _T_43 : _GEN_5398; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5400 = 6'h18 == _T_664 ? _T_44 : _GEN_5399; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5401 = 6'h19 == _T_664 ? _T_45 : _GEN_5400; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5402 = 6'h1a == _T_664 ? _T_46 : _GEN_5401; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5403 = 6'h1b == _T_664 ? _T_47 : _GEN_5402; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5404 = 6'h1c == _T_664 ? _T_48 : _GEN_5403; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5405 = 6'h1d == _T_664 ? _T_49 : _GEN_5404; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5406 = 6'h1e == _T_664 ? _T_50 : _GEN_5405; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5407 = 6'h1f == _T_664 ? _T_51 : _GEN_5406; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5408 = 6'h20 == _T_664 ? _T_52 : _GEN_5407; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5409 = 6'h21 == _T_664 ? _T_53 : _GEN_5408; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5410 = 6'h22 == _T_664 ? _T_54 : _GEN_5409; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5411 = 6'h23 == _T_664 ? _T_55 : _GEN_5410; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5412 = 6'h24 == _T_664 ? _T_56 : _GEN_5411; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5413 = 6'h25 == _T_664 ? _T_57 : _GEN_5412; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5414 = 6'h26 == _T_664 ? _T_58 : _GEN_5413; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5415 = 6'h27 == _T_664 ? _T_59 : _GEN_5414; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5416 = 6'h28 == _T_664 ? _T_60 : _GEN_5415; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5417 = 6'h29 == _T_664 ? _T_61 : _GEN_5416; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5418 = 6'h2a == _T_664 ? _T_62 : _GEN_5417; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5419 = 6'h2b == _T_664 ? _T_63 : _GEN_5418; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5420 = 6'h2c == _T_664 ? _T_64 : _GEN_5419; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5421 = 6'h2d == _T_664 ? _T_65 : _GEN_5420; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5422 = 6'h2e == _T_664 ? _T_66 : _GEN_5421; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5423 = 6'h2f == _T_664 ? _T_67 : _GEN_5422; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5424 = 6'h30 == _T_664 ? _T_68 : _GEN_5423; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5425 = 6'h31 == _T_664 ? _T_69 : _GEN_5424; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5426 = 6'h32 == _T_664 ? _T_70 : _GEN_5425; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5427 = 6'h33 == _T_664 ? _T_71 : _GEN_5426; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5428 = 6'h34 == _T_664 ? _T_72 : _GEN_5427; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5429 = 6'h35 == _T_664 ? _T_73 : _GEN_5428; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5430 = 6'h36 == _T_664 ? _T_74 : _GEN_5429; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5431 = 6'h37 == _T_664 ? _T_75 : _GEN_5430; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5432 = 6'h38 == _T_664 ? _T_76 : _GEN_5431; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5433 = 6'h39 == _T_664 ? _T_77 : _GEN_5432; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5434 = 6'h3a == _T_664 ? _T_78 : _GEN_5433; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5435 = 6'h3b == _T_664 ? _T_79 : _GEN_5434; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5436 = 6'h3c == _T_664 ? _T_80 : _GEN_5435; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5437 = 6'h3d == _T_664 ? _T_81 : _GEN_5436; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5438 = 6'h3e == _T_664 ? _T_82 : _GEN_5437; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5439 = 6'h3f == _T_664 ? _T_83 : _GEN_5438; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5441 = 6'h1 == _T_668 ? _T_21 : _T_20; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5442 = 6'h2 == _T_668 ? _T_22 : _GEN_5441; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5443 = 6'h3 == _T_668 ? _T_23 : _GEN_5442; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5444 = 6'h4 == _T_668 ? _T_24 : _GEN_5443; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5445 = 6'h5 == _T_668 ? _T_25 : _GEN_5444; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5446 = 6'h6 == _T_668 ? _T_26 : _GEN_5445; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5447 = 6'h7 == _T_668 ? _T_27 : _GEN_5446; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5448 = 6'h8 == _T_668 ? _T_28 : _GEN_5447; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5449 = 6'h9 == _T_668 ? _T_29 : _GEN_5448; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5450 = 6'ha == _T_668 ? _T_30 : _GEN_5449; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5451 = 6'hb == _T_668 ? _T_31 : _GEN_5450; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5452 = 6'hc == _T_668 ? _T_32 : _GEN_5451; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5453 = 6'hd == _T_668 ? _T_33 : _GEN_5452; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5454 = 6'he == _T_668 ? _T_34 : _GEN_5453; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5455 = 6'hf == _T_668 ? _T_35 : _GEN_5454; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5456 = 6'h10 == _T_668 ? _T_36 : _GEN_5455; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5457 = 6'h11 == _T_668 ? _T_37 : _GEN_5456; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5458 = 6'h12 == _T_668 ? _T_38 : _GEN_5457; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5459 = 6'h13 == _T_668 ? _T_39 : _GEN_5458; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5460 = 6'h14 == _T_668 ? _T_40 : _GEN_5459; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5461 = 6'h15 == _T_668 ? _T_41 : _GEN_5460; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5462 = 6'h16 == _T_668 ? _T_42 : _GEN_5461; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5463 = 6'h17 == _T_668 ? _T_43 : _GEN_5462; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5464 = 6'h18 == _T_668 ? _T_44 : _GEN_5463; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5465 = 6'h19 == _T_668 ? _T_45 : _GEN_5464; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5466 = 6'h1a == _T_668 ? _T_46 : _GEN_5465; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5467 = 6'h1b == _T_668 ? _T_47 : _GEN_5466; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5468 = 6'h1c == _T_668 ? _T_48 : _GEN_5467; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5469 = 6'h1d == _T_668 ? _T_49 : _GEN_5468; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5470 = 6'h1e == _T_668 ? _T_50 : _GEN_5469; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5471 = 6'h1f == _T_668 ? _T_51 : _GEN_5470; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5472 = 6'h20 == _T_668 ? _T_52 : _GEN_5471; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5473 = 6'h21 == _T_668 ? _T_53 : _GEN_5472; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5474 = 6'h22 == _T_668 ? _T_54 : _GEN_5473; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5475 = 6'h23 == _T_668 ? _T_55 : _GEN_5474; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5476 = 6'h24 == _T_668 ? _T_56 : _GEN_5475; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5477 = 6'h25 == _T_668 ? _T_57 : _GEN_5476; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5478 = 6'h26 == _T_668 ? _T_58 : _GEN_5477; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5479 = 6'h27 == _T_668 ? _T_59 : _GEN_5478; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5480 = 6'h28 == _T_668 ? _T_60 : _GEN_5479; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5481 = 6'h29 == _T_668 ? _T_61 : _GEN_5480; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5482 = 6'h2a == _T_668 ? _T_62 : _GEN_5481; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5483 = 6'h2b == _T_668 ? _T_63 : _GEN_5482; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5484 = 6'h2c == _T_668 ? _T_64 : _GEN_5483; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5485 = 6'h2d == _T_668 ? _T_65 : _GEN_5484; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5486 = 6'h2e == _T_668 ? _T_66 : _GEN_5485; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5487 = 6'h2f == _T_668 ? _T_67 : _GEN_5486; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5488 = 6'h30 == _T_668 ? _T_68 : _GEN_5487; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5489 = 6'h31 == _T_668 ? _T_69 : _GEN_5488; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5490 = 6'h32 == _T_668 ? _T_70 : _GEN_5489; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5491 = 6'h33 == _T_668 ? _T_71 : _GEN_5490; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5492 = 6'h34 == _T_668 ? _T_72 : _GEN_5491; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5493 = 6'h35 == _T_668 ? _T_73 : _GEN_5492; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5494 = 6'h36 == _T_668 ? _T_74 : _GEN_5493; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5495 = 6'h37 == _T_668 ? _T_75 : _GEN_5494; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5496 = 6'h38 == _T_668 ? _T_76 : _GEN_5495; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5497 = 6'h39 == _T_668 ? _T_77 : _GEN_5496; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5498 = 6'h3a == _T_668 ? _T_78 : _GEN_5497; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5499 = 6'h3b == _T_668 ? _T_79 : _GEN_5498; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5500 = 6'h3c == _T_668 ? _T_80 : _GEN_5499; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5501 = 6'h3d == _T_668 ? _T_81 : _GEN_5500; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5502 = 6'h3e == _T_668 ? _T_82 : _GEN_5501; // @[execute.scala 79:10:@2151.4]
  assign _GEN_5503 = 6'h3f == _T_668 ? _T_83 : _GEN_5502; // @[execute.scala 79:10:@2151.4]
  assign _T_670 = _T_660 ? _GEN_5439 : _GEN_5503; // @[execute.scala 79:10:@2151.4]
  assign _T_672 = io_amount < 6'h15; // @[execute.scala 79:15:@2152.4]
  assign _T_674 = io_amount - 6'h15; // @[execute.scala 79:37:@2153.4]
  assign _T_675 = $unsigned(_T_674); // @[execute.scala 79:37:@2154.4]
  assign _T_676 = _T_675[5:0]; // @[execute.scala 79:37:@2155.4]
  assign _T_679 = 6'h2b + io_amount; // @[execute.scala 79:60:@2156.4]
  assign _T_680 = 6'h2b + io_amount; // @[execute.scala 79:60:@2157.4]
  assign _GEN_5505 = 6'h1 == _T_676 ? _T_21 : _T_20; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5506 = 6'h2 == _T_676 ? _T_22 : _GEN_5505; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5507 = 6'h3 == _T_676 ? _T_23 : _GEN_5506; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5508 = 6'h4 == _T_676 ? _T_24 : _GEN_5507; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5509 = 6'h5 == _T_676 ? _T_25 : _GEN_5508; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5510 = 6'h6 == _T_676 ? _T_26 : _GEN_5509; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5511 = 6'h7 == _T_676 ? _T_27 : _GEN_5510; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5512 = 6'h8 == _T_676 ? _T_28 : _GEN_5511; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5513 = 6'h9 == _T_676 ? _T_29 : _GEN_5512; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5514 = 6'ha == _T_676 ? _T_30 : _GEN_5513; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5515 = 6'hb == _T_676 ? _T_31 : _GEN_5514; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5516 = 6'hc == _T_676 ? _T_32 : _GEN_5515; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5517 = 6'hd == _T_676 ? _T_33 : _GEN_5516; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5518 = 6'he == _T_676 ? _T_34 : _GEN_5517; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5519 = 6'hf == _T_676 ? _T_35 : _GEN_5518; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5520 = 6'h10 == _T_676 ? _T_36 : _GEN_5519; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5521 = 6'h11 == _T_676 ? _T_37 : _GEN_5520; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5522 = 6'h12 == _T_676 ? _T_38 : _GEN_5521; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5523 = 6'h13 == _T_676 ? _T_39 : _GEN_5522; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5524 = 6'h14 == _T_676 ? _T_40 : _GEN_5523; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5525 = 6'h15 == _T_676 ? _T_41 : _GEN_5524; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5526 = 6'h16 == _T_676 ? _T_42 : _GEN_5525; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5527 = 6'h17 == _T_676 ? _T_43 : _GEN_5526; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5528 = 6'h18 == _T_676 ? _T_44 : _GEN_5527; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5529 = 6'h19 == _T_676 ? _T_45 : _GEN_5528; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5530 = 6'h1a == _T_676 ? _T_46 : _GEN_5529; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5531 = 6'h1b == _T_676 ? _T_47 : _GEN_5530; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5532 = 6'h1c == _T_676 ? _T_48 : _GEN_5531; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5533 = 6'h1d == _T_676 ? _T_49 : _GEN_5532; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5534 = 6'h1e == _T_676 ? _T_50 : _GEN_5533; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5535 = 6'h1f == _T_676 ? _T_51 : _GEN_5534; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5536 = 6'h20 == _T_676 ? _T_52 : _GEN_5535; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5537 = 6'h21 == _T_676 ? _T_53 : _GEN_5536; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5538 = 6'h22 == _T_676 ? _T_54 : _GEN_5537; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5539 = 6'h23 == _T_676 ? _T_55 : _GEN_5538; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5540 = 6'h24 == _T_676 ? _T_56 : _GEN_5539; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5541 = 6'h25 == _T_676 ? _T_57 : _GEN_5540; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5542 = 6'h26 == _T_676 ? _T_58 : _GEN_5541; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5543 = 6'h27 == _T_676 ? _T_59 : _GEN_5542; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5544 = 6'h28 == _T_676 ? _T_60 : _GEN_5543; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5545 = 6'h29 == _T_676 ? _T_61 : _GEN_5544; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5546 = 6'h2a == _T_676 ? _T_62 : _GEN_5545; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5547 = 6'h2b == _T_676 ? _T_63 : _GEN_5546; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5548 = 6'h2c == _T_676 ? _T_64 : _GEN_5547; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5549 = 6'h2d == _T_676 ? _T_65 : _GEN_5548; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5550 = 6'h2e == _T_676 ? _T_66 : _GEN_5549; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5551 = 6'h2f == _T_676 ? _T_67 : _GEN_5550; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5552 = 6'h30 == _T_676 ? _T_68 : _GEN_5551; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5553 = 6'h31 == _T_676 ? _T_69 : _GEN_5552; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5554 = 6'h32 == _T_676 ? _T_70 : _GEN_5553; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5555 = 6'h33 == _T_676 ? _T_71 : _GEN_5554; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5556 = 6'h34 == _T_676 ? _T_72 : _GEN_5555; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5557 = 6'h35 == _T_676 ? _T_73 : _GEN_5556; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5558 = 6'h36 == _T_676 ? _T_74 : _GEN_5557; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5559 = 6'h37 == _T_676 ? _T_75 : _GEN_5558; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5560 = 6'h38 == _T_676 ? _T_76 : _GEN_5559; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5561 = 6'h39 == _T_676 ? _T_77 : _GEN_5560; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5562 = 6'h3a == _T_676 ? _T_78 : _GEN_5561; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5563 = 6'h3b == _T_676 ? _T_79 : _GEN_5562; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5564 = 6'h3c == _T_676 ? _T_80 : _GEN_5563; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5565 = 6'h3d == _T_676 ? _T_81 : _GEN_5564; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5566 = 6'h3e == _T_676 ? _T_82 : _GEN_5565; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5567 = 6'h3f == _T_676 ? _T_83 : _GEN_5566; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5569 = 6'h1 == _T_680 ? _T_21 : _T_20; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5570 = 6'h2 == _T_680 ? _T_22 : _GEN_5569; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5571 = 6'h3 == _T_680 ? _T_23 : _GEN_5570; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5572 = 6'h4 == _T_680 ? _T_24 : _GEN_5571; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5573 = 6'h5 == _T_680 ? _T_25 : _GEN_5572; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5574 = 6'h6 == _T_680 ? _T_26 : _GEN_5573; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5575 = 6'h7 == _T_680 ? _T_27 : _GEN_5574; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5576 = 6'h8 == _T_680 ? _T_28 : _GEN_5575; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5577 = 6'h9 == _T_680 ? _T_29 : _GEN_5576; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5578 = 6'ha == _T_680 ? _T_30 : _GEN_5577; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5579 = 6'hb == _T_680 ? _T_31 : _GEN_5578; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5580 = 6'hc == _T_680 ? _T_32 : _GEN_5579; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5581 = 6'hd == _T_680 ? _T_33 : _GEN_5580; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5582 = 6'he == _T_680 ? _T_34 : _GEN_5581; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5583 = 6'hf == _T_680 ? _T_35 : _GEN_5582; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5584 = 6'h10 == _T_680 ? _T_36 : _GEN_5583; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5585 = 6'h11 == _T_680 ? _T_37 : _GEN_5584; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5586 = 6'h12 == _T_680 ? _T_38 : _GEN_5585; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5587 = 6'h13 == _T_680 ? _T_39 : _GEN_5586; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5588 = 6'h14 == _T_680 ? _T_40 : _GEN_5587; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5589 = 6'h15 == _T_680 ? _T_41 : _GEN_5588; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5590 = 6'h16 == _T_680 ? _T_42 : _GEN_5589; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5591 = 6'h17 == _T_680 ? _T_43 : _GEN_5590; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5592 = 6'h18 == _T_680 ? _T_44 : _GEN_5591; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5593 = 6'h19 == _T_680 ? _T_45 : _GEN_5592; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5594 = 6'h1a == _T_680 ? _T_46 : _GEN_5593; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5595 = 6'h1b == _T_680 ? _T_47 : _GEN_5594; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5596 = 6'h1c == _T_680 ? _T_48 : _GEN_5595; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5597 = 6'h1d == _T_680 ? _T_49 : _GEN_5596; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5598 = 6'h1e == _T_680 ? _T_50 : _GEN_5597; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5599 = 6'h1f == _T_680 ? _T_51 : _GEN_5598; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5600 = 6'h20 == _T_680 ? _T_52 : _GEN_5599; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5601 = 6'h21 == _T_680 ? _T_53 : _GEN_5600; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5602 = 6'h22 == _T_680 ? _T_54 : _GEN_5601; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5603 = 6'h23 == _T_680 ? _T_55 : _GEN_5602; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5604 = 6'h24 == _T_680 ? _T_56 : _GEN_5603; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5605 = 6'h25 == _T_680 ? _T_57 : _GEN_5604; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5606 = 6'h26 == _T_680 ? _T_58 : _GEN_5605; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5607 = 6'h27 == _T_680 ? _T_59 : _GEN_5606; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5608 = 6'h28 == _T_680 ? _T_60 : _GEN_5607; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5609 = 6'h29 == _T_680 ? _T_61 : _GEN_5608; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5610 = 6'h2a == _T_680 ? _T_62 : _GEN_5609; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5611 = 6'h2b == _T_680 ? _T_63 : _GEN_5610; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5612 = 6'h2c == _T_680 ? _T_64 : _GEN_5611; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5613 = 6'h2d == _T_680 ? _T_65 : _GEN_5612; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5614 = 6'h2e == _T_680 ? _T_66 : _GEN_5613; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5615 = 6'h2f == _T_680 ? _T_67 : _GEN_5614; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5616 = 6'h30 == _T_680 ? _T_68 : _GEN_5615; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5617 = 6'h31 == _T_680 ? _T_69 : _GEN_5616; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5618 = 6'h32 == _T_680 ? _T_70 : _GEN_5617; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5619 = 6'h33 == _T_680 ? _T_71 : _GEN_5618; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5620 = 6'h34 == _T_680 ? _T_72 : _GEN_5619; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5621 = 6'h35 == _T_680 ? _T_73 : _GEN_5620; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5622 = 6'h36 == _T_680 ? _T_74 : _GEN_5621; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5623 = 6'h37 == _T_680 ? _T_75 : _GEN_5622; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5624 = 6'h38 == _T_680 ? _T_76 : _GEN_5623; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5625 = 6'h39 == _T_680 ? _T_77 : _GEN_5624; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5626 = 6'h3a == _T_680 ? _T_78 : _GEN_5625; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5627 = 6'h3b == _T_680 ? _T_79 : _GEN_5626; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5628 = 6'h3c == _T_680 ? _T_80 : _GEN_5627; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5629 = 6'h3d == _T_680 ? _T_81 : _GEN_5628; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5630 = 6'h3e == _T_680 ? _T_82 : _GEN_5629; // @[execute.scala 79:10:@2158.4]
  assign _GEN_5631 = 6'h3f == _T_680 ? _T_83 : _GEN_5630; // @[execute.scala 79:10:@2158.4]
  assign _T_682 = _T_672 ? _GEN_5567 : _GEN_5631; // @[execute.scala 79:10:@2158.4]
  assign _T_684 = io_amount < 6'h14; // @[execute.scala 79:15:@2159.4]
  assign _T_686 = io_amount - 6'h14; // @[execute.scala 79:37:@2160.4]
  assign _T_687 = $unsigned(_T_686); // @[execute.scala 79:37:@2161.4]
  assign _T_688 = _T_687[5:0]; // @[execute.scala 79:37:@2162.4]
  assign _T_691 = 6'h2c + io_amount; // @[execute.scala 79:60:@2163.4]
  assign _T_692 = 6'h2c + io_amount; // @[execute.scala 79:60:@2164.4]
  assign _GEN_5633 = 6'h1 == _T_688 ? _T_21 : _T_20; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5634 = 6'h2 == _T_688 ? _T_22 : _GEN_5633; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5635 = 6'h3 == _T_688 ? _T_23 : _GEN_5634; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5636 = 6'h4 == _T_688 ? _T_24 : _GEN_5635; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5637 = 6'h5 == _T_688 ? _T_25 : _GEN_5636; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5638 = 6'h6 == _T_688 ? _T_26 : _GEN_5637; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5639 = 6'h7 == _T_688 ? _T_27 : _GEN_5638; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5640 = 6'h8 == _T_688 ? _T_28 : _GEN_5639; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5641 = 6'h9 == _T_688 ? _T_29 : _GEN_5640; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5642 = 6'ha == _T_688 ? _T_30 : _GEN_5641; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5643 = 6'hb == _T_688 ? _T_31 : _GEN_5642; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5644 = 6'hc == _T_688 ? _T_32 : _GEN_5643; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5645 = 6'hd == _T_688 ? _T_33 : _GEN_5644; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5646 = 6'he == _T_688 ? _T_34 : _GEN_5645; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5647 = 6'hf == _T_688 ? _T_35 : _GEN_5646; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5648 = 6'h10 == _T_688 ? _T_36 : _GEN_5647; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5649 = 6'h11 == _T_688 ? _T_37 : _GEN_5648; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5650 = 6'h12 == _T_688 ? _T_38 : _GEN_5649; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5651 = 6'h13 == _T_688 ? _T_39 : _GEN_5650; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5652 = 6'h14 == _T_688 ? _T_40 : _GEN_5651; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5653 = 6'h15 == _T_688 ? _T_41 : _GEN_5652; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5654 = 6'h16 == _T_688 ? _T_42 : _GEN_5653; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5655 = 6'h17 == _T_688 ? _T_43 : _GEN_5654; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5656 = 6'h18 == _T_688 ? _T_44 : _GEN_5655; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5657 = 6'h19 == _T_688 ? _T_45 : _GEN_5656; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5658 = 6'h1a == _T_688 ? _T_46 : _GEN_5657; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5659 = 6'h1b == _T_688 ? _T_47 : _GEN_5658; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5660 = 6'h1c == _T_688 ? _T_48 : _GEN_5659; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5661 = 6'h1d == _T_688 ? _T_49 : _GEN_5660; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5662 = 6'h1e == _T_688 ? _T_50 : _GEN_5661; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5663 = 6'h1f == _T_688 ? _T_51 : _GEN_5662; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5664 = 6'h20 == _T_688 ? _T_52 : _GEN_5663; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5665 = 6'h21 == _T_688 ? _T_53 : _GEN_5664; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5666 = 6'h22 == _T_688 ? _T_54 : _GEN_5665; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5667 = 6'h23 == _T_688 ? _T_55 : _GEN_5666; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5668 = 6'h24 == _T_688 ? _T_56 : _GEN_5667; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5669 = 6'h25 == _T_688 ? _T_57 : _GEN_5668; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5670 = 6'h26 == _T_688 ? _T_58 : _GEN_5669; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5671 = 6'h27 == _T_688 ? _T_59 : _GEN_5670; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5672 = 6'h28 == _T_688 ? _T_60 : _GEN_5671; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5673 = 6'h29 == _T_688 ? _T_61 : _GEN_5672; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5674 = 6'h2a == _T_688 ? _T_62 : _GEN_5673; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5675 = 6'h2b == _T_688 ? _T_63 : _GEN_5674; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5676 = 6'h2c == _T_688 ? _T_64 : _GEN_5675; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5677 = 6'h2d == _T_688 ? _T_65 : _GEN_5676; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5678 = 6'h2e == _T_688 ? _T_66 : _GEN_5677; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5679 = 6'h2f == _T_688 ? _T_67 : _GEN_5678; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5680 = 6'h30 == _T_688 ? _T_68 : _GEN_5679; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5681 = 6'h31 == _T_688 ? _T_69 : _GEN_5680; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5682 = 6'h32 == _T_688 ? _T_70 : _GEN_5681; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5683 = 6'h33 == _T_688 ? _T_71 : _GEN_5682; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5684 = 6'h34 == _T_688 ? _T_72 : _GEN_5683; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5685 = 6'h35 == _T_688 ? _T_73 : _GEN_5684; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5686 = 6'h36 == _T_688 ? _T_74 : _GEN_5685; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5687 = 6'h37 == _T_688 ? _T_75 : _GEN_5686; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5688 = 6'h38 == _T_688 ? _T_76 : _GEN_5687; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5689 = 6'h39 == _T_688 ? _T_77 : _GEN_5688; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5690 = 6'h3a == _T_688 ? _T_78 : _GEN_5689; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5691 = 6'h3b == _T_688 ? _T_79 : _GEN_5690; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5692 = 6'h3c == _T_688 ? _T_80 : _GEN_5691; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5693 = 6'h3d == _T_688 ? _T_81 : _GEN_5692; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5694 = 6'h3e == _T_688 ? _T_82 : _GEN_5693; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5695 = 6'h3f == _T_688 ? _T_83 : _GEN_5694; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5697 = 6'h1 == _T_692 ? _T_21 : _T_20; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5698 = 6'h2 == _T_692 ? _T_22 : _GEN_5697; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5699 = 6'h3 == _T_692 ? _T_23 : _GEN_5698; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5700 = 6'h4 == _T_692 ? _T_24 : _GEN_5699; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5701 = 6'h5 == _T_692 ? _T_25 : _GEN_5700; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5702 = 6'h6 == _T_692 ? _T_26 : _GEN_5701; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5703 = 6'h7 == _T_692 ? _T_27 : _GEN_5702; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5704 = 6'h8 == _T_692 ? _T_28 : _GEN_5703; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5705 = 6'h9 == _T_692 ? _T_29 : _GEN_5704; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5706 = 6'ha == _T_692 ? _T_30 : _GEN_5705; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5707 = 6'hb == _T_692 ? _T_31 : _GEN_5706; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5708 = 6'hc == _T_692 ? _T_32 : _GEN_5707; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5709 = 6'hd == _T_692 ? _T_33 : _GEN_5708; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5710 = 6'he == _T_692 ? _T_34 : _GEN_5709; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5711 = 6'hf == _T_692 ? _T_35 : _GEN_5710; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5712 = 6'h10 == _T_692 ? _T_36 : _GEN_5711; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5713 = 6'h11 == _T_692 ? _T_37 : _GEN_5712; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5714 = 6'h12 == _T_692 ? _T_38 : _GEN_5713; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5715 = 6'h13 == _T_692 ? _T_39 : _GEN_5714; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5716 = 6'h14 == _T_692 ? _T_40 : _GEN_5715; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5717 = 6'h15 == _T_692 ? _T_41 : _GEN_5716; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5718 = 6'h16 == _T_692 ? _T_42 : _GEN_5717; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5719 = 6'h17 == _T_692 ? _T_43 : _GEN_5718; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5720 = 6'h18 == _T_692 ? _T_44 : _GEN_5719; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5721 = 6'h19 == _T_692 ? _T_45 : _GEN_5720; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5722 = 6'h1a == _T_692 ? _T_46 : _GEN_5721; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5723 = 6'h1b == _T_692 ? _T_47 : _GEN_5722; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5724 = 6'h1c == _T_692 ? _T_48 : _GEN_5723; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5725 = 6'h1d == _T_692 ? _T_49 : _GEN_5724; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5726 = 6'h1e == _T_692 ? _T_50 : _GEN_5725; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5727 = 6'h1f == _T_692 ? _T_51 : _GEN_5726; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5728 = 6'h20 == _T_692 ? _T_52 : _GEN_5727; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5729 = 6'h21 == _T_692 ? _T_53 : _GEN_5728; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5730 = 6'h22 == _T_692 ? _T_54 : _GEN_5729; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5731 = 6'h23 == _T_692 ? _T_55 : _GEN_5730; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5732 = 6'h24 == _T_692 ? _T_56 : _GEN_5731; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5733 = 6'h25 == _T_692 ? _T_57 : _GEN_5732; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5734 = 6'h26 == _T_692 ? _T_58 : _GEN_5733; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5735 = 6'h27 == _T_692 ? _T_59 : _GEN_5734; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5736 = 6'h28 == _T_692 ? _T_60 : _GEN_5735; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5737 = 6'h29 == _T_692 ? _T_61 : _GEN_5736; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5738 = 6'h2a == _T_692 ? _T_62 : _GEN_5737; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5739 = 6'h2b == _T_692 ? _T_63 : _GEN_5738; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5740 = 6'h2c == _T_692 ? _T_64 : _GEN_5739; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5741 = 6'h2d == _T_692 ? _T_65 : _GEN_5740; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5742 = 6'h2e == _T_692 ? _T_66 : _GEN_5741; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5743 = 6'h2f == _T_692 ? _T_67 : _GEN_5742; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5744 = 6'h30 == _T_692 ? _T_68 : _GEN_5743; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5745 = 6'h31 == _T_692 ? _T_69 : _GEN_5744; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5746 = 6'h32 == _T_692 ? _T_70 : _GEN_5745; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5747 = 6'h33 == _T_692 ? _T_71 : _GEN_5746; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5748 = 6'h34 == _T_692 ? _T_72 : _GEN_5747; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5749 = 6'h35 == _T_692 ? _T_73 : _GEN_5748; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5750 = 6'h36 == _T_692 ? _T_74 : _GEN_5749; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5751 = 6'h37 == _T_692 ? _T_75 : _GEN_5750; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5752 = 6'h38 == _T_692 ? _T_76 : _GEN_5751; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5753 = 6'h39 == _T_692 ? _T_77 : _GEN_5752; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5754 = 6'h3a == _T_692 ? _T_78 : _GEN_5753; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5755 = 6'h3b == _T_692 ? _T_79 : _GEN_5754; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5756 = 6'h3c == _T_692 ? _T_80 : _GEN_5755; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5757 = 6'h3d == _T_692 ? _T_81 : _GEN_5756; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5758 = 6'h3e == _T_692 ? _T_82 : _GEN_5757; // @[execute.scala 79:10:@2165.4]
  assign _GEN_5759 = 6'h3f == _T_692 ? _T_83 : _GEN_5758; // @[execute.scala 79:10:@2165.4]
  assign _T_694 = _T_684 ? _GEN_5695 : _GEN_5759; // @[execute.scala 79:10:@2165.4]
  assign _T_696 = io_amount < 6'h13; // @[execute.scala 79:15:@2166.4]
  assign _T_698 = io_amount - 6'h13; // @[execute.scala 79:37:@2167.4]
  assign _T_699 = $unsigned(_T_698); // @[execute.scala 79:37:@2168.4]
  assign _T_700 = _T_699[5:0]; // @[execute.scala 79:37:@2169.4]
  assign _T_703 = 6'h2d + io_amount; // @[execute.scala 79:60:@2170.4]
  assign _T_704 = 6'h2d + io_amount; // @[execute.scala 79:60:@2171.4]
  assign _GEN_5761 = 6'h1 == _T_700 ? _T_21 : _T_20; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5762 = 6'h2 == _T_700 ? _T_22 : _GEN_5761; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5763 = 6'h3 == _T_700 ? _T_23 : _GEN_5762; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5764 = 6'h4 == _T_700 ? _T_24 : _GEN_5763; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5765 = 6'h5 == _T_700 ? _T_25 : _GEN_5764; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5766 = 6'h6 == _T_700 ? _T_26 : _GEN_5765; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5767 = 6'h7 == _T_700 ? _T_27 : _GEN_5766; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5768 = 6'h8 == _T_700 ? _T_28 : _GEN_5767; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5769 = 6'h9 == _T_700 ? _T_29 : _GEN_5768; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5770 = 6'ha == _T_700 ? _T_30 : _GEN_5769; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5771 = 6'hb == _T_700 ? _T_31 : _GEN_5770; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5772 = 6'hc == _T_700 ? _T_32 : _GEN_5771; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5773 = 6'hd == _T_700 ? _T_33 : _GEN_5772; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5774 = 6'he == _T_700 ? _T_34 : _GEN_5773; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5775 = 6'hf == _T_700 ? _T_35 : _GEN_5774; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5776 = 6'h10 == _T_700 ? _T_36 : _GEN_5775; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5777 = 6'h11 == _T_700 ? _T_37 : _GEN_5776; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5778 = 6'h12 == _T_700 ? _T_38 : _GEN_5777; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5779 = 6'h13 == _T_700 ? _T_39 : _GEN_5778; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5780 = 6'h14 == _T_700 ? _T_40 : _GEN_5779; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5781 = 6'h15 == _T_700 ? _T_41 : _GEN_5780; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5782 = 6'h16 == _T_700 ? _T_42 : _GEN_5781; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5783 = 6'h17 == _T_700 ? _T_43 : _GEN_5782; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5784 = 6'h18 == _T_700 ? _T_44 : _GEN_5783; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5785 = 6'h19 == _T_700 ? _T_45 : _GEN_5784; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5786 = 6'h1a == _T_700 ? _T_46 : _GEN_5785; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5787 = 6'h1b == _T_700 ? _T_47 : _GEN_5786; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5788 = 6'h1c == _T_700 ? _T_48 : _GEN_5787; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5789 = 6'h1d == _T_700 ? _T_49 : _GEN_5788; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5790 = 6'h1e == _T_700 ? _T_50 : _GEN_5789; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5791 = 6'h1f == _T_700 ? _T_51 : _GEN_5790; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5792 = 6'h20 == _T_700 ? _T_52 : _GEN_5791; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5793 = 6'h21 == _T_700 ? _T_53 : _GEN_5792; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5794 = 6'h22 == _T_700 ? _T_54 : _GEN_5793; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5795 = 6'h23 == _T_700 ? _T_55 : _GEN_5794; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5796 = 6'h24 == _T_700 ? _T_56 : _GEN_5795; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5797 = 6'h25 == _T_700 ? _T_57 : _GEN_5796; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5798 = 6'h26 == _T_700 ? _T_58 : _GEN_5797; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5799 = 6'h27 == _T_700 ? _T_59 : _GEN_5798; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5800 = 6'h28 == _T_700 ? _T_60 : _GEN_5799; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5801 = 6'h29 == _T_700 ? _T_61 : _GEN_5800; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5802 = 6'h2a == _T_700 ? _T_62 : _GEN_5801; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5803 = 6'h2b == _T_700 ? _T_63 : _GEN_5802; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5804 = 6'h2c == _T_700 ? _T_64 : _GEN_5803; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5805 = 6'h2d == _T_700 ? _T_65 : _GEN_5804; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5806 = 6'h2e == _T_700 ? _T_66 : _GEN_5805; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5807 = 6'h2f == _T_700 ? _T_67 : _GEN_5806; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5808 = 6'h30 == _T_700 ? _T_68 : _GEN_5807; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5809 = 6'h31 == _T_700 ? _T_69 : _GEN_5808; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5810 = 6'h32 == _T_700 ? _T_70 : _GEN_5809; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5811 = 6'h33 == _T_700 ? _T_71 : _GEN_5810; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5812 = 6'h34 == _T_700 ? _T_72 : _GEN_5811; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5813 = 6'h35 == _T_700 ? _T_73 : _GEN_5812; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5814 = 6'h36 == _T_700 ? _T_74 : _GEN_5813; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5815 = 6'h37 == _T_700 ? _T_75 : _GEN_5814; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5816 = 6'h38 == _T_700 ? _T_76 : _GEN_5815; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5817 = 6'h39 == _T_700 ? _T_77 : _GEN_5816; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5818 = 6'h3a == _T_700 ? _T_78 : _GEN_5817; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5819 = 6'h3b == _T_700 ? _T_79 : _GEN_5818; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5820 = 6'h3c == _T_700 ? _T_80 : _GEN_5819; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5821 = 6'h3d == _T_700 ? _T_81 : _GEN_5820; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5822 = 6'h3e == _T_700 ? _T_82 : _GEN_5821; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5823 = 6'h3f == _T_700 ? _T_83 : _GEN_5822; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5825 = 6'h1 == _T_704 ? _T_21 : _T_20; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5826 = 6'h2 == _T_704 ? _T_22 : _GEN_5825; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5827 = 6'h3 == _T_704 ? _T_23 : _GEN_5826; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5828 = 6'h4 == _T_704 ? _T_24 : _GEN_5827; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5829 = 6'h5 == _T_704 ? _T_25 : _GEN_5828; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5830 = 6'h6 == _T_704 ? _T_26 : _GEN_5829; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5831 = 6'h7 == _T_704 ? _T_27 : _GEN_5830; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5832 = 6'h8 == _T_704 ? _T_28 : _GEN_5831; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5833 = 6'h9 == _T_704 ? _T_29 : _GEN_5832; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5834 = 6'ha == _T_704 ? _T_30 : _GEN_5833; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5835 = 6'hb == _T_704 ? _T_31 : _GEN_5834; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5836 = 6'hc == _T_704 ? _T_32 : _GEN_5835; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5837 = 6'hd == _T_704 ? _T_33 : _GEN_5836; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5838 = 6'he == _T_704 ? _T_34 : _GEN_5837; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5839 = 6'hf == _T_704 ? _T_35 : _GEN_5838; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5840 = 6'h10 == _T_704 ? _T_36 : _GEN_5839; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5841 = 6'h11 == _T_704 ? _T_37 : _GEN_5840; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5842 = 6'h12 == _T_704 ? _T_38 : _GEN_5841; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5843 = 6'h13 == _T_704 ? _T_39 : _GEN_5842; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5844 = 6'h14 == _T_704 ? _T_40 : _GEN_5843; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5845 = 6'h15 == _T_704 ? _T_41 : _GEN_5844; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5846 = 6'h16 == _T_704 ? _T_42 : _GEN_5845; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5847 = 6'h17 == _T_704 ? _T_43 : _GEN_5846; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5848 = 6'h18 == _T_704 ? _T_44 : _GEN_5847; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5849 = 6'h19 == _T_704 ? _T_45 : _GEN_5848; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5850 = 6'h1a == _T_704 ? _T_46 : _GEN_5849; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5851 = 6'h1b == _T_704 ? _T_47 : _GEN_5850; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5852 = 6'h1c == _T_704 ? _T_48 : _GEN_5851; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5853 = 6'h1d == _T_704 ? _T_49 : _GEN_5852; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5854 = 6'h1e == _T_704 ? _T_50 : _GEN_5853; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5855 = 6'h1f == _T_704 ? _T_51 : _GEN_5854; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5856 = 6'h20 == _T_704 ? _T_52 : _GEN_5855; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5857 = 6'h21 == _T_704 ? _T_53 : _GEN_5856; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5858 = 6'h22 == _T_704 ? _T_54 : _GEN_5857; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5859 = 6'h23 == _T_704 ? _T_55 : _GEN_5858; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5860 = 6'h24 == _T_704 ? _T_56 : _GEN_5859; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5861 = 6'h25 == _T_704 ? _T_57 : _GEN_5860; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5862 = 6'h26 == _T_704 ? _T_58 : _GEN_5861; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5863 = 6'h27 == _T_704 ? _T_59 : _GEN_5862; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5864 = 6'h28 == _T_704 ? _T_60 : _GEN_5863; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5865 = 6'h29 == _T_704 ? _T_61 : _GEN_5864; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5866 = 6'h2a == _T_704 ? _T_62 : _GEN_5865; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5867 = 6'h2b == _T_704 ? _T_63 : _GEN_5866; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5868 = 6'h2c == _T_704 ? _T_64 : _GEN_5867; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5869 = 6'h2d == _T_704 ? _T_65 : _GEN_5868; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5870 = 6'h2e == _T_704 ? _T_66 : _GEN_5869; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5871 = 6'h2f == _T_704 ? _T_67 : _GEN_5870; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5872 = 6'h30 == _T_704 ? _T_68 : _GEN_5871; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5873 = 6'h31 == _T_704 ? _T_69 : _GEN_5872; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5874 = 6'h32 == _T_704 ? _T_70 : _GEN_5873; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5875 = 6'h33 == _T_704 ? _T_71 : _GEN_5874; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5876 = 6'h34 == _T_704 ? _T_72 : _GEN_5875; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5877 = 6'h35 == _T_704 ? _T_73 : _GEN_5876; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5878 = 6'h36 == _T_704 ? _T_74 : _GEN_5877; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5879 = 6'h37 == _T_704 ? _T_75 : _GEN_5878; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5880 = 6'h38 == _T_704 ? _T_76 : _GEN_5879; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5881 = 6'h39 == _T_704 ? _T_77 : _GEN_5880; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5882 = 6'h3a == _T_704 ? _T_78 : _GEN_5881; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5883 = 6'h3b == _T_704 ? _T_79 : _GEN_5882; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5884 = 6'h3c == _T_704 ? _T_80 : _GEN_5883; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5885 = 6'h3d == _T_704 ? _T_81 : _GEN_5884; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5886 = 6'h3e == _T_704 ? _T_82 : _GEN_5885; // @[execute.scala 79:10:@2172.4]
  assign _GEN_5887 = 6'h3f == _T_704 ? _T_83 : _GEN_5886; // @[execute.scala 79:10:@2172.4]
  assign _T_706 = _T_696 ? _GEN_5823 : _GEN_5887; // @[execute.scala 79:10:@2172.4]
  assign _T_708 = io_amount < 6'h12; // @[execute.scala 79:15:@2173.4]
  assign _T_710 = io_amount - 6'h12; // @[execute.scala 79:37:@2174.4]
  assign _T_711 = $unsigned(_T_710); // @[execute.scala 79:37:@2175.4]
  assign _T_712 = _T_711[5:0]; // @[execute.scala 79:37:@2176.4]
  assign _T_715 = 6'h2e + io_amount; // @[execute.scala 79:60:@2177.4]
  assign _T_716 = 6'h2e + io_amount; // @[execute.scala 79:60:@2178.4]
  assign _GEN_5889 = 6'h1 == _T_712 ? _T_21 : _T_20; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5890 = 6'h2 == _T_712 ? _T_22 : _GEN_5889; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5891 = 6'h3 == _T_712 ? _T_23 : _GEN_5890; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5892 = 6'h4 == _T_712 ? _T_24 : _GEN_5891; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5893 = 6'h5 == _T_712 ? _T_25 : _GEN_5892; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5894 = 6'h6 == _T_712 ? _T_26 : _GEN_5893; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5895 = 6'h7 == _T_712 ? _T_27 : _GEN_5894; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5896 = 6'h8 == _T_712 ? _T_28 : _GEN_5895; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5897 = 6'h9 == _T_712 ? _T_29 : _GEN_5896; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5898 = 6'ha == _T_712 ? _T_30 : _GEN_5897; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5899 = 6'hb == _T_712 ? _T_31 : _GEN_5898; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5900 = 6'hc == _T_712 ? _T_32 : _GEN_5899; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5901 = 6'hd == _T_712 ? _T_33 : _GEN_5900; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5902 = 6'he == _T_712 ? _T_34 : _GEN_5901; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5903 = 6'hf == _T_712 ? _T_35 : _GEN_5902; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5904 = 6'h10 == _T_712 ? _T_36 : _GEN_5903; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5905 = 6'h11 == _T_712 ? _T_37 : _GEN_5904; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5906 = 6'h12 == _T_712 ? _T_38 : _GEN_5905; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5907 = 6'h13 == _T_712 ? _T_39 : _GEN_5906; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5908 = 6'h14 == _T_712 ? _T_40 : _GEN_5907; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5909 = 6'h15 == _T_712 ? _T_41 : _GEN_5908; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5910 = 6'h16 == _T_712 ? _T_42 : _GEN_5909; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5911 = 6'h17 == _T_712 ? _T_43 : _GEN_5910; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5912 = 6'h18 == _T_712 ? _T_44 : _GEN_5911; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5913 = 6'h19 == _T_712 ? _T_45 : _GEN_5912; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5914 = 6'h1a == _T_712 ? _T_46 : _GEN_5913; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5915 = 6'h1b == _T_712 ? _T_47 : _GEN_5914; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5916 = 6'h1c == _T_712 ? _T_48 : _GEN_5915; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5917 = 6'h1d == _T_712 ? _T_49 : _GEN_5916; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5918 = 6'h1e == _T_712 ? _T_50 : _GEN_5917; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5919 = 6'h1f == _T_712 ? _T_51 : _GEN_5918; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5920 = 6'h20 == _T_712 ? _T_52 : _GEN_5919; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5921 = 6'h21 == _T_712 ? _T_53 : _GEN_5920; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5922 = 6'h22 == _T_712 ? _T_54 : _GEN_5921; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5923 = 6'h23 == _T_712 ? _T_55 : _GEN_5922; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5924 = 6'h24 == _T_712 ? _T_56 : _GEN_5923; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5925 = 6'h25 == _T_712 ? _T_57 : _GEN_5924; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5926 = 6'h26 == _T_712 ? _T_58 : _GEN_5925; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5927 = 6'h27 == _T_712 ? _T_59 : _GEN_5926; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5928 = 6'h28 == _T_712 ? _T_60 : _GEN_5927; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5929 = 6'h29 == _T_712 ? _T_61 : _GEN_5928; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5930 = 6'h2a == _T_712 ? _T_62 : _GEN_5929; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5931 = 6'h2b == _T_712 ? _T_63 : _GEN_5930; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5932 = 6'h2c == _T_712 ? _T_64 : _GEN_5931; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5933 = 6'h2d == _T_712 ? _T_65 : _GEN_5932; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5934 = 6'h2e == _T_712 ? _T_66 : _GEN_5933; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5935 = 6'h2f == _T_712 ? _T_67 : _GEN_5934; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5936 = 6'h30 == _T_712 ? _T_68 : _GEN_5935; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5937 = 6'h31 == _T_712 ? _T_69 : _GEN_5936; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5938 = 6'h32 == _T_712 ? _T_70 : _GEN_5937; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5939 = 6'h33 == _T_712 ? _T_71 : _GEN_5938; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5940 = 6'h34 == _T_712 ? _T_72 : _GEN_5939; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5941 = 6'h35 == _T_712 ? _T_73 : _GEN_5940; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5942 = 6'h36 == _T_712 ? _T_74 : _GEN_5941; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5943 = 6'h37 == _T_712 ? _T_75 : _GEN_5942; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5944 = 6'h38 == _T_712 ? _T_76 : _GEN_5943; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5945 = 6'h39 == _T_712 ? _T_77 : _GEN_5944; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5946 = 6'h3a == _T_712 ? _T_78 : _GEN_5945; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5947 = 6'h3b == _T_712 ? _T_79 : _GEN_5946; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5948 = 6'h3c == _T_712 ? _T_80 : _GEN_5947; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5949 = 6'h3d == _T_712 ? _T_81 : _GEN_5948; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5950 = 6'h3e == _T_712 ? _T_82 : _GEN_5949; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5951 = 6'h3f == _T_712 ? _T_83 : _GEN_5950; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5953 = 6'h1 == _T_716 ? _T_21 : _T_20; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5954 = 6'h2 == _T_716 ? _T_22 : _GEN_5953; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5955 = 6'h3 == _T_716 ? _T_23 : _GEN_5954; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5956 = 6'h4 == _T_716 ? _T_24 : _GEN_5955; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5957 = 6'h5 == _T_716 ? _T_25 : _GEN_5956; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5958 = 6'h6 == _T_716 ? _T_26 : _GEN_5957; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5959 = 6'h7 == _T_716 ? _T_27 : _GEN_5958; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5960 = 6'h8 == _T_716 ? _T_28 : _GEN_5959; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5961 = 6'h9 == _T_716 ? _T_29 : _GEN_5960; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5962 = 6'ha == _T_716 ? _T_30 : _GEN_5961; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5963 = 6'hb == _T_716 ? _T_31 : _GEN_5962; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5964 = 6'hc == _T_716 ? _T_32 : _GEN_5963; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5965 = 6'hd == _T_716 ? _T_33 : _GEN_5964; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5966 = 6'he == _T_716 ? _T_34 : _GEN_5965; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5967 = 6'hf == _T_716 ? _T_35 : _GEN_5966; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5968 = 6'h10 == _T_716 ? _T_36 : _GEN_5967; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5969 = 6'h11 == _T_716 ? _T_37 : _GEN_5968; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5970 = 6'h12 == _T_716 ? _T_38 : _GEN_5969; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5971 = 6'h13 == _T_716 ? _T_39 : _GEN_5970; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5972 = 6'h14 == _T_716 ? _T_40 : _GEN_5971; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5973 = 6'h15 == _T_716 ? _T_41 : _GEN_5972; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5974 = 6'h16 == _T_716 ? _T_42 : _GEN_5973; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5975 = 6'h17 == _T_716 ? _T_43 : _GEN_5974; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5976 = 6'h18 == _T_716 ? _T_44 : _GEN_5975; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5977 = 6'h19 == _T_716 ? _T_45 : _GEN_5976; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5978 = 6'h1a == _T_716 ? _T_46 : _GEN_5977; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5979 = 6'h1b == _T_716 ? _T_47 : _GEN_5978; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5980 = 6'h1c == _T_716 ? _T_48 : _GEN_5979; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5981 = 6'h1d == _T_716 ? _T_49 : _GEN_5980; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5982 = 6'h1e == _T_716 ? _T_50 : _GEN_5981; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5983 = 6'h1f == _T_716 ? _T_51 : _GEN_5982; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5984 = 6'h20 == _T_716 ? _T_52 : _GEN_5983; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5985 = 6'h21 == _T_716 ? _T_53 : _GEN_5984; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5986 = 6'h22 == _T_716 ? _T_54 : _GEN_5985; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5987 = 6'h23 == _T_716 ? _T_55 : _GEN_5986; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5988 = 6'h24 == _T_716 ? _T_56 : _GEN_5987; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5989 = 6'h25 == _T_716 ? _T_57 : _GEN_5988; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5990 = 6'h26 == _T_716 ? _T_58 : _GEN_5989; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5991 = 6'h27 == _T_716 ? _T_59 : _GEN_5990; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5992 = 6'h28 == _T_716 ? _T_60 : _GEN_5991; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5993 = 6'h29 == _T_716 ? _T_61 : _GEN_5992; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5994 = 6'h2a == _T_716 ? _T_62 : _GEN_5993; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5995 = 6'h2b == _T_716 ? _T_63 : _GEN_5994; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5996 = 6'h2c == _T_716 ? _T_64 : _GEN_5995; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5997 = 6'h2d == _T_716 ? _T_65 : _GEN_5996; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5998 = 6'h2e == _T_716 ? _T_66 : _GEN_5997; // @[execute.scala 79:10:@2179.4]
  assign _GEN_5999 = 6'h2f == _T_716 ? _T_67 : _GEN_5998; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6000 = 6'h30 == _T_716 ? _T_68 : _GEN_5999; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6001 = 6'h31 == _T_716 ? _T_69 : _GEN_6000; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6002 = 6'h32 == _T_716 ? _T_70 : _GEN_6001; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6003 = 6'h33 == _T_716 ? _T_71 : _GEN_6002; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6004 = 6'h34 == _T_716 ? _T_72 : _GEN_6003; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6005 = 6'h35 == _T_716 ? _T_73 : _GEN_6004; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6006 = 6'h36 == _T_716 ? _T_74 : _GEN_6005; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6007 = 6'h37 == _T_716 ? _T_75 : _GEN_6006; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6008 = 6'h38 == _T_716 ? _T_76 : _GEN_6007; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6009 = 6'h39 == _T_716 ? _T_77 : _GEN_6008; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6010 = 6'h3a == _T_716 ? _T_78 : _GEN_6009; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6011 = 6'h3b == _T_716 ? _T_79 : _GEN_6010; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6012 = 6'h3c == _T_716 ? _T_80 : _GEN_6011; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6013 = 6'h3d == _T_716 ? _T_81 : _GEN_6012; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6014 = 6'h3e == _T_716 ? _T_82 : _GEN_6013; // @[execute.scala 79:10:@2179.4]
  assign _GEN_6015 = 6'h3f == _T_716 ? _T_83 : _GEN_6014; // @[execute.scala 79:10:@2179.4]
  assign _T_718 = _T_708 ? _GEN_5951 : _GEN_6015; // @[execute.scala 79:10:@2179.4]
  assign _T_720 = io_amount < 6'h11; // @[execute.scala 79:15:@2180.4]
  assign _T_722 = io_amount - 6'h11; // @[execute.scala 79:37:@2181.4]
  assign _T_723 = $unsigned(_T_722); // @[execute.scala 79:37:@2182.4]
  assign _T_724 = _T_723[5:0]; // @[execute.scala 79:37:@2183.4]
  assign _T_727 = 6'h2f + io_amount; // @[execute.scala 79:60:@2184.4]
  assign _T_728 = 6'h2f + io_amount; // @[execute.scala 79:60:@2185.4]
  assign _GEN_6017 = 6'h1 == _T_724 ? _T_21 : _T_20; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6018 = 6'h2 == _T_724 ? _T_22 : _GEN_6017; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6019 = 6'h3 == _T_724 ? _T_23 : _GEN_6018; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6020 = 6'h4 == _T_724 ? _T_24 : _GEN_6019; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6021 = 6'h5 == _T_724 ? _T_25 : _GEN_6020; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6022 = 6'h6 == _T_724 ? _T_26 : _GEN_6021; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6023 = 6'h7 == _T_724 ? _T_27 : _GEN_6022; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6024 = 6'h8 == _T_724 ? _T_28 : _GEN_6023; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6025 = 6'h9 == _T_724 ? _T_29 : _GEN_6024; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6026 = 6'ha == _T_724 ? _T_30 : _GEN_6025; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6027 = 6'hb == _T_724 ? _T_31 : _GEN_6026; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6028 = 6'hc == _T_724 ? _T_32 : _GEN_6027; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6029 = 6'hd == _T_724 ? _T_33 : _GEN_6028; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6030 = 6'he == _T_724 ? _T_34 : _GEN_6029; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6031 = 6'hf == _T_724 ? _T_35 : _GEN_6030; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6032 = 6'h10 == _T_724 ? _T_36 : _GEN_6031; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6033 = 6'h11 == _T_724 ? _T_37 : _GEN_6032; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6034 = 6'h12 == _T_724 ? _T_38 : _GEN_6033; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6035 = 6'h13 == _T_724 ? _T_39 : _GEN_6034; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6036 = 6'h14 == _T_724 ? _T_40 : _GEN_6035; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6037 = 6'h15 == _T_724 ? _T_41 : _GEN_6036; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6038 = 6'h16 == _T_724 ? _T_42 : _GEN_6037; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6039 = 6'h17 == _T_724 ? _T_43 : _GEN_6038; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6040 = 6'h18 == _T_724 ? _T_44 : _GEN_6039; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6041 = 6'h19 == _T_724 ? _T_45 : _GEN_6040; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6042 = 6'h1a == _T_724 ? _T_46 : _GEN_6041; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6043 = 6'h1b == _T_724 ? _T_47 : _GEN_6042; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6044 = 6'h1c == _T_724 ? _T_48 : _GEN_6043; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6045 = 6'h1d == _T_724 ? _T_49 : _GEN_6044; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6046 = 6'h1e == _T_724 ? _T_50 : _GEN_6045; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6047 = 6'h1f == _T_724 ? _T_51 : _GEN_6046; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6048 = 6'h20 == _T_724 ? _T_52 : _GEN_6047; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6049 = 6'h21 == _T_724 ? _T_53 : _GEN_6048; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6050 = 6'h22 == _T_724 ? _T_54 : _GEN_6049; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6051 = 6'h23 == _T_724 ? _T_55 : _GEN_6050; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6052 = 6'h24 == _T_724 ? _T_56 : _GEN_6051; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6053 = 6'h25 == _T_724 ? _T_57 : _GEN_6052; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6054 = 6'h26 == _T_724 ? _T_58 : _GEN_6053; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6055 = 6'h27 == _T_724 ? _T_59 : _GEN_6054; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6056 = 6'h28 == _T_724 ? _T_60 : _GEN_6055; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6057 = 6'h29 == _T_724 ? _T_61 : _GEN_6056; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6058 = 6'h2a == _T_724 ? _T_62 : _GEN_6057; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6059 = 6'h2b == _T_724 ? _T_63 : _GEN_6058; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6060 = 6'h2c == _T_724 ? _T_64 : _GEN_6059; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6061 = 6'h2d == _T_724 ? _T_65 : _GEN_6060; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6062 = 6'h2e == _T_724 ? _T_66 : _GEN_6061; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6063 = 6'h2f == _T_724 ? _T_67 : _GEN_6062; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6064 = 6'h30 == _T_724 ? _T_68 : _GEN_6063; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6065 = 6'h31 == _T_724 ? _T_69 : _GEN_6064; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6066 = 6'h32 == _T_724 ? _T_70 : _GEN_6065; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6067 = 6'h33 == _T_724 ? _T_71 : _GEN_6066; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6068 = 6'h34 == _T_724 ? _T_72 : _GEN_6067; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6069 = 6'h35 == _T_724 ? _T_73 : _GEN_6068; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6070 = 6'h36 == _T_724 ? _T_74 : _GEN_6069; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6071 = 6'h37 == _T_724 ? _T_75 : _GEN_6070; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6072 = 6'h38 == _T_724 ? _T_76 : _GEN_6071; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6073 = 6'h39 == _T_724 ? _T_77 : _GEN_6072; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6074 = 6'h3a == _T_724 ? _T_78 : _GEN_6073; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6075 = 6'h3b == _T_724 ? _T_79 : _GEN_6074; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6076 = 6'h3c == _T_724 ? _T_80 : _GEN_6075; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6077 = 6'h3d == _T_724 ? _T_81 : _GEN_6076; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6078 = 6'h3e == _T_724 ? _T_82 : _GEN_6077; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6079 = 6'h3f == _T_724 ? _T_83 : _GEN_6078; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6081 = 6'h1 == _T_728 ? _T_21 : _T_20; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6082 = 6'h2 == _T_728 ? _T_22 : _GEN_6081; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6083 = 6'h3 == _T_728 ? _T_23 : _GEN_6082; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6084 = 6'h4 == _T_728 ? _T_24 : _GEN_6083; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6085 = 6'h5 == _T_728 ? _T_25 : _GEN_6084; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6086 = 6'h6 == _T_728 ? _T_26 : _GEN_6085; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6087 = 6'h7 == _T_728 ? _T_27 : _GEN_6086; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6088 = 6'h8 == _T_728 ? _T_28 : _GEN_6087; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6089 = 6'h9 == _T_728 ? _T_29 : _GEN_6088; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6090 = 6'ha == _T_728 ? _T_30 : _GEN_6089; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6091 = 6'hb == _T_728 ? _T_31 : _GEN_6090; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6092 = 6'hc == _T_728 ? _T_32 : _GEN_6091; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6093 = 6'hd == _T_728 ? _T_33 : _GEN_6092; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6094 = 6'he == _T_728 ? _T_34 : _GEN_6093; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6095 = 6'hf == _T_728 ? _T_35 : _GEN_6094; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6096 = 6'h10 == _T_728 ? _T_36 : _GEN_6095; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6097 = 6'h11 == _T_728 ? _T_37 : _GEN_6096; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6098 = 6'h12 == _T_728 ? _T_38 : _GEN_6097; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6099 = 6'h13 == _T_728 ? _T_39 : _GEN_6098; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6100 = 6'h14 == _T_728 ? _T_40 : _GEN_6099; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6101 = 6'h15 == _T_728 ? _T_41 : _GEN_6100; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6102 = 6'h16 == _T_728 ? _T_42 : _GEN_6101; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6103 = 6'h17 == _T_728 ? _T_43 : _GEN_6102; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6104 = 6'h18 == _T_728 ? _T_44 : _GEN_6103; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6105 = 6'h19 == _T_728 ? _T_45 : _GEN_6104; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6106 = 6'h1a == _T_728 ? _T_46 : _GEN_6105; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6107 = 6'h1b == _T_728 ? _T_47 : _GEN_6106; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6108 = 6'h1c == _T_728 ? _T_48 : _GEN_6107; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6109 = 6'h1d == _T_728 ? _T_49 : _GEN_6108; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6110 = 6'h1e == _T_728 ? _T_50 : _GEN_6109; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6111 = 6'h1f == _T_728 ? _T_51 : _GEN_6110; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6112 = 6'h20 == _T_728 ? _T_52 : _GEN_6111; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6113 = 6'h21 == _T_728 ? _T_53 : _GEN_6112; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6114 = 6'h22 == _T_728 ? _T_54 : _GEN_6113; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6115 = 6'h23 == _T_728 ? _T_55 : _GEN_6114; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6116 = 6'h24 == _T_728 ? _T_56 : _GEN_6115; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6117 = 6'h25 == _T_728 ? _T_57 : _GEN_6116; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6118 = 6'h26 == _T_728 ? _T_58 : _GEN_6117; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6119 = 6'h27 == _T_728 ? _T_59 : _GEN_6118; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6120 = 6'h28 == _T_728 ? _T_60 : _GEN_6119; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6121 = 6'h29 == _T_728 ? _T_61 : _GEN_6120; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6122 = 6'h2a == _T_728 ? _T_62 : _GEN_6121; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6123 = 6'h2b == _T_728 ? _T_63 : _GEN_6122; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6124 = 6'h2c == _T_728 ? _T_64 : _GEN_6123; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6125 = 6'h2d == _T_728 ? _T_65 : _GEN_6124; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6126 = 6'h2e == _T_728 ? _T_66 : _GEN_6125; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6127 = 6'h2f == _T_728 ? _T_67 : _GEN_6126; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6128 = 6'h30 == _T_728 ? _T_68 : _GEN_6127; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6129 = 6'h31 == _T_728 ? _T_69 : _GEN_6128; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6130 = 6'h32 == _T_728 ? _T_70 : _GEN_6129; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6131 = 6'h33 == _T_728 ? _T_71 : _GEN_6130; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6132 = 6'h34 == _T_728 ? _T_72 : _GEN_6131; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6133 = 6'h35 == _T_728 ? _T_73 : _GEN_6132; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6134 = 6'h36 == _T_728 ? _T_74 : _GEN_6133; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6135 = 6'h37 == _T_728 ? _T_75 : _GEN_6134; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6136 = 6'h38 == _T_728 ? _T_76 : _GEN_6135; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6137 = 6'h39 == _T_728 ? _T_77 : _GEN_6136; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6138 = 6'h3a == _T_728 ? _T_78 : _GEN_6137; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6139 = 6'h3b == _T_728 ? _T_79 : _GEN_6138; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6140 = 6'h3c == _T_728 ? _T_80 : _GEN_6139; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6141 = 6'h3d == _T_728 ? _T_81 : _GEN_6140; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6142 = 6'h3e == _T_728 ? _T_82 : _GEN_6141; // @[execute.scala 79:10:@2186.4]
  assign _GEN_6143 = 6'h3f == _T_728 ? _T_83 : _GEN_6142; // @[execute.scala 79:10:@2186.4]
  assign _T_730 = _T_720 ? _GEN_6079 : _GEN_6143; // @[execute.scala 79:10:@2186.4]
  assign _T_732 = io_amount < 6'h10; // @[execute.scala 79:15:@2187.4]
  assign _T_734 = io_amount - 6'h10; // @[execute.scala 79:37:@2188.4]
  assign _T_735 = $unsigned(_T_734); // @[execute.scala 79:37:@2189.4]
  assign _T_736 = _T_735[5:0]; // @[execute.scala 79:37:@2190.4]
  assign _T_739 = 6'h30 + io_amount; // @[execute.scala 79:60:@2191.4]
  assign _T_740 = 6'h30 + io_amount; // @[execute.scala 79:60:@2192.4]
  assign _GEN_6145 = 6'h1 == _T_736 ? _T_21 : _T_20; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6146 = 6'h2 == _T_736 ? _T_22 : _GEN_6145; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6147 = 6'h3 == _T_736 ? _T_23 : _GEN_6146; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6148 = 6'h4 == _T_736 ? _T_24 : _GEN_6147; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6149 = 6'h5 == _T_736 ? _T_25 : _GEN_6148; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6150 = 6'h6 == _T_736 ? _T_26 : _GEN_6149; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6151 = 6'h7 == _T_736 ? _T_27 : _GEN_6150; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6152 = 6'h8 == _T_736 ? _T_28 : _GEN_6151; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6153 = 6'h9 == _T_736 ? _T_29 : _GEN_6152; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6154 = 6'ha == _T_736 ? _T_30 : _GEN_6153; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6155 = 6'hb == _T_736 ? _T_31 : _GEN_6154; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6156 = 6'hc == _T_736 ? _T_32 : _GEN_6155; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6157 = 6'hd == _T_736 ? _T_33 : _GEN_6156; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6158 = 6'he == _T_736 ? _T_34 : _GEN_6157; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6159 = 6'hf == _T_736 ? _T_35 : _GEN_6158; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6160 = 6'h10 == _T_736 ? _T_36 : _GEN_6159; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6161 = 6'h11 == _T_736 ? _T_37 : _GEN_6160; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6162 = 6'h12 == _T_736 ? _T_38 : _GEN_6161; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6163 = 6'h13 == _T_736 ? _T_39 : _GEN_6162; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6164 = 6'h14 == _T_736 ? _T_40 : _GEN_6163; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6165 = 6'h15 == _T_736 ? _T_41 : _GEN_6164; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6166 = 6'h16 == _T_736 ? _T_42 : _GEN_6165; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6167 = 6'h17 == _T_736 ? _T_43 : _GEN_6166; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6168 = 6'h18 == _T_736 ? _T_44 : _GEN_6167; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6169 = 6'h19 == _T_736 ? _T_45 : _GEN_6168; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6170 = 6'h1a == _T_736 ? _T_46 : _GEN_6169; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6171 = 6'h1b == _T_736 ? _T_47 : _GEN_6170; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6172 = 6'h1c == _T_736 ? _T_48 : _GEN_6171; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6173 = 6'h1d == _T_736 ? _T_49 : _GEN_6172; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6174 = 6'h1e == _T_736 ? _T_50 : _GEN_6173; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6175 = 6'h1f == _T_736 ? _T_51 : _GEN_6174; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6176 = 6'h20 == _T_736 ? _T_52 : _GEN_6175; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6177 = 6'h21 == _T_736 ? _T_53 : _GEN_6176; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6178 = 6'h22 == _T_736 ? _T_54 : _GEN_6177; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6179 = 6'h23 == _T_736 ? _T_55 : _GEN_6178; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6180 = 6'h24 == _T_736 ? _T_56 : _GEN_6179; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6181 = 6'h25 == _T_736 ? _T_57 : _GEN_6180; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6182 = 6'h26 == _T_736 ? _T_58 : _GEN_6181; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6183 = 6'h27 == _T_736 ? _T_59 : _GEN_6182; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6184 = 6'h28 == _T_736 ? _T_60 : _GEN_6183; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6185 = 6'h29 == _T_736 ? _T_61 : _GEN_6184; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6186 = 6'h2a == _T_736 ? _T_62 : _GEN_6185; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6187 = 6'h2b == _T_736 ? _T_63 : _GEN_6186; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6188 = 6'h2c == _T_736 ? _T_64 : _GEN_6187; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6189 = 6'h2d == _T_736 ? _T_65 : _GEN_6188; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6190 = 6'h2e == _T_736 ? _T_66 : _GEN_6189; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6191 = 6'h2f == _T_736 ? _T_67 : _GEN_6190; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6192 = 6'h30 == _T_736 ? _T_68 : _GEN_6191; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6193 = 6'h31 == _T_736 ? _T_69 : _GEN_6192; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6194 = 6'h32 == _T_736 ? _T_70 : _GEN_6193; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6195 = 6'h33 == _T_736 ? _T_71 : _GEN_6194; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6196 = 6'h34 == _T_736 ? _T_72 : _GEN_6195; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6197 = 6'h35 == _T_736 ? _T_73 : _GEN_6196; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6198 = 6'h36 == _T_736 ? _T_74 : _GEN_6197; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6199 = 6'h37 == _T_736 ? _T_75 : _GEN_6198; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6200 = 6'h38 == _T_736 ? _T_76 : _GEN_6199; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6201 = 6'h39 == _T_736 ? _T_77 : _GEN_6200; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6202 = 6'h3a == _T_736 ? _T_78 : _GEN_6201; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6203 = 6'h3b == _T_736 ? _T_79 : _GEN_6202; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6204 = 6'h3c == _T_736 ? _T_80 : _GEN_6203; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6205 = 6'h3d == _T_736 ? _T_81 : _GEN_6204; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6206 = 6'h3e == _T_736 ? _T_82 : _GEN_6205; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6207 = 6'h3f == _T_736 ? _T_83 : _GEN_6206; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6209 = 6'h1 == _T_740 ? _T_21 : _T_20; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6210 = 6'h2 == _T_740 ? _T_22 : _GEN_6209; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6211 = 6'h3 == _T_740 ? _T_23 : _GEN_6210; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6212 = 6'h4 == _T_740 ? _T_24 : _GEN_6211; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6213 = 6'h5 == _T_740 ? _T_25 : _GEN_6212; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6214 = 6'h6 == _T_740 ? _T_26 : _GEN_6213; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6215 = 6'h7 == _T_740 ? _T_27 : _GEN_6214; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6216 = 6'h8 == _T_740 ? _T_28 : _GEN_6215; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6217 = 6'h9 == _T_740 ? _T_29 : _GEN_6216; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6218 = 6'ha == _T_740 ? _T_30 : _GEN_6217; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6219 = 6'hb == _T_740 ? _T_31 : _GEN_6218; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6220 = 6'hc == _T_740 ? _T_32 : _GEN_6219; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6221 = 6'hd == _T_740 ? _T_33 : _GEN_6220; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6222 = 6'he == _T_740 ? _T_34 : _GEN_6221; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6223 = 6'hf == _T_740 ? _T_35 : _GEN_6222; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6224 = 6'h10 == _T_740 ? _T_36 : _GEN_6223; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6225 = 6'h11 == _T_740 ? _T_37 : _GEN_6224; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6226 = 6'h12 == _T_740 ? _T_38 : _GEN_6225; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6227 = 6'h13 == _T_740 ? _T_39 : _GEN_6226; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6228 = 6'h14 == _T_740 ? _T_40 : _GEN_6227; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6229 = 6'h15 == _T_740 ? _T_41 : _GEN_6228; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6230 = 6'h16 == _T_740 ? _T_42 : _GEN_6229; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6231 = 6'h17 == _T_740 ? _T_43 : _GEN_6230; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6232 = 6'h18 == _T_740 ? _T_44 : _GEN_6231; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6233 = 6'h19 == _T_740 ? _T_45 : _GEN_6232; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6234 = 6'h1a == _T_740 ? _T_46 : _GEN_6233; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6235 = 6'h1b == _T_740 ? _T_47 : _GEN_6234; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6236 = 6'h1c == _T_740 ? _T_48 : _GEN_6235; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6237 = 6'h1d == _T_740 ? _T_49 : _GEN_6236; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6238 = 6'h1e == _T_740 ? _T_50 : _GEN_6237; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6239 = 6'h1f == _T_740 ? _T_51 : _GEN_6238; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6240 = 6'h20 == _T_740 ? _T_52 : _GEN_6239; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6241 = 6'h21 == _T_740 ? _T_53 : _GEN_6240; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6242 = 6'h22 == _T_740 ? _T_54 : _GEN_6241; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6243 = 6'h23 == _T_740 ? _T_55 : _GEN_6242; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6244 = 6'h24 == _T_740 ? _T_56 : _GEN_6243; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6245 = 6'h25 == _T_740 ? _T_57 : _GEN_6244; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6246 = 6'h26 == _T_740 ? _T_58 : _GEN_6245; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6247 = 6'h27 == _T_740 ? _T_59 : _GEN_6246; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6248 = 6'h28 == _T_740 ? _T_60 : _GEN_6247; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6249 = 6'h29 == _T_740 ? _T_61 : _GEN_6248; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6250 = 6'h2a == _T_740 ? _T_62 : _GEN_6249; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6251 = 6'h2b == _T_740 ? _T_63 : _GEN_6250; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6252 = 6'h2c == _T_740 ? _T_64 : _GEN_6251; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6253 = 6'h2d == _T_740 ? _T_65 : _GEN_6252; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6254 = 6'h2e == _T_740 ? _T_66 : _GEN_6253; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6255 = 6'h2f == _T_740 ? _T_67 : _GEN_6254; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6256 = 6'h30 == _T_740 ? _T_68 : _GEN_6255; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6257 = 6'h31 == _T_740 ? _T_69 : _GEN_6256; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6258 = 6'h32 == _T_740 ? _T_70 : _GEN_6257; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6259 = 6'h33 == _T_740 ? _T_71 : _GEN_6258; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6260 = 6'h34 == _T_740 ? _T_72 : _GEN_6259; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6261 = 6'h35 == _T_740 ? _T_73 : _GEN_6260; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6262 = 6'h36 == _T_740 ? _T_74 : _GEN_6261; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6263 = 6'h37 == _T_740 ? _T_75 : _GEN_6262; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6264 = 6'h38 == _T_740 ? _T_76 : _GEN_6263; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6265 = 6'h39 == _T_740 ? _T_77 : _GEN_6264; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6266 = 6'h3a == _T_740 ? _T_78 : _GEN_6265; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6267 = 6'h3b == _T_740 ? _T_79 : _GEN_6266; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6268 = 6'h3c == _T_740 ? _T_80 : _GEN_6267; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6269 = 6'h3d == _T_740 ? _T_81 : _GEN_6268; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6270 = 6'h3e == _T_740 ? _T_82 : _GEN_6269; // @[execute.scala 79:10:@2193.4]
  assign _GEN_6271 = 6'h3f == _T_740 ? _T_83 : _GEN_6270; // @[execute.scala 79:10:@2193.4]
  assign _T_742 = _T_732 ? _GEN_6207 : _GEN_6271; // @[execute.scala 79:10:@2193.4]
  assign _T_744 = io_amount < 6'hf; // @[execute.scala 79:15:@2194.4]
  assign _T_746 = io_amount - 6'hf; // @[execute.scala 79:37:@2195.4]
  assign _T_747 = $unsigned(_T_746); // @[execute.scala 79:37:@2196.4]
  assign _T_748 = _T_747[5:0]; // @[execute.scala 79:37:@2197.4]
  assign _T_751 = 6'h31 + io_amount; // @[execute.scala 79:60:@2198.4]
  assign _T_752 = 6'h31 + io_amount; // @[execute.scala 79:60:@2199.4]
  assign _GEN_6273 = 6'h1 == _T_748 ? _T_21 : _T_20; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6274 = 6'h2 == _T_748 ? _T_22 : _GEN_6273; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6275 = 6'h3 == _T_748 ? _T_23 : _GEN_6274; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6276 = 6'h4 == _T_748 ? _T_24 : _GEN_6275; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6277 = 6'h5 == _T_748 ? _T_25 : _GEN_6276; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6278 = 6'h6 == _T_748 ? _T_26 : _GEN_6277; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6279 = 6'h7 == _T_748 ? _T_27 : _GEN_6278; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6280 = 6'h8 == _T_748 ? _T_28 : _GEN_6279; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6281 = 6'h9 == _T_748 ? _T_29 : _GEN_6280; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6282 = 6'ha == _T_748 ? _T_30 : _GEN_6281; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6283 = 6'hb == _T_748 ? _T_31 : _GEN_6282; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6284 = 6'hc == _T_748 ? _T_32 : _GEN_6283; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6285 = 6'hd == _T_748 ? _T_33 : _GEN_6284; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6286 = 6'he == _T_748 ? _T_34 : _GEN_6285; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6287 = 6'hf == _T_748 ? _T_35 : _GEN_6286; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6288 = 6'h10 == _T_748 ? _T_36 : _GEN_6287; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6289 = 6'h11 == _T_748 ? _T_37 : _GEN_6288; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6290 = 6'h12 == _T_748 ? _T_38 : _GEN_6289; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6291 = 6'h13 == _T_748 ? _T_39 : _GEN_6290; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6292 = 6'h14 == _T_748 ? _T_40 : _GEN_6291; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6293 = 6'h15 == _T_748 ? _T_41 : _GEN_6292; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6294 = 6'h16 == _T_748 ? _T_42 : _GEN_6293; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6295 = 6'h17 == _T_748 ? _T_43 : _GEN_6294; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6296 = 6'h18 == _T_748 ? _T_44 : _GEN_6295; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6297 = 6'h19 == _T_748 ? _T_45 : _GEN_6296; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6298 = 6'h1a == _T_748 ? _T_46 : _GEN_6297; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6299 = 6'h1b == _T_748 ? _T_47 : _GEN_6298; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6300 = 6'h1c == _T_748 ? _T_48 : _GEN_6299; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6301 = 6'h1d == _T_748 ? _T_49 : _GEN_6300; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6302 = 6'h1e == _T_748 ? _T_50 : _GEN_6301; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6303 = 6'h1f == _T_748 ? _T_51 : _GEN_6302; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6304 = 6'h20 == _T_748 ? _T_52 : _GEN_6303; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6305 = 6'h21 == _T_748 ? _T_53 : _GEN_6304; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6306 = 6'h22 == _T_748 ? _T_54 : _GEN_6305; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6307 = 6'h23 == _T_748 ? _T_55 : _GEN_6306; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6308 = 6'h24 == _T_748 ? _T_56 : _GEN_6307; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6309 = 6'h25 == _T_748 ? _T_57 : _GEN_6308; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6310 = 6'h26 == _T_748 ? _T_58 : _GEN_6309; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6311 = 6'h27 == _T_748 ? _T_59 : _GEN_6310; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6312 = 6'h28 == _T_748 ? _T_60 : _GEN_6311; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6313 = 6'h29 == _T_748 ? _T_61 : _GEN_6312; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6314 = 6'h2a == _T_748 ? _T_62 : _GEN_6313; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6315 = 6'h2b == _T_748 ? _T_63 : _GEN_6314; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6316 = 6'h2c == _T_748 ? _T_64 : _GEN_6315; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6317 = 6'h2d == _T_748 ? _T_65 : _GEN_6316; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6318 = 6'h2e == _T_748 ? _T_66 : _GEN_6317; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6319 = 6'h2f == _T_748 ? _T_67 : _GEN_6318; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6320 = 6'h30 == _T_748 ? _T_68 : _GEN_6319; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6321 = 6'h31 == _T_748 ? _T_69 : _GEN_6320; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6322 = 6'h32 == _T_748 ? _T_70 : _GEN_6321; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6323 = 6'h33 == _T_748 ? _T_71 : _GEN_6322; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6324 = 6'h34 == _T_748 ? _T_72 : _GEN_6323; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6325 = 6'h35 == _T_748 ? _T_73 : _GEN_6324; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6326 = 6'h36 == _T_748 ? _T_74 : _GEN_6325; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6327 = 6'h37 == _T_748 ? _T_75 : _GEN_6326; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6328 = 6'h38 == _T_748 ? _T_76 : _GEN_6327; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6329 = 6'h39 == _T_748 ? _T_77 : _GEN_6328; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6330 = 6'h3a == _T_748 ? _T_78 : _GEN_6329; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6331 = 6'h3b == _T_748 ? _T_79 : _GEN_6330; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6332 = 6'h3c == _T_748 ? _T_80 : _GEN_6331; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6333 = 6'h3d == _T_748 ? _T_81 : _GEN_6332; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6334 = 6'h3e == _T_748 ? _T_82 : _GEN_6333; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6335 = 6'h3f == _T_748 ? _T_83 : _GEN_6334; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6337 = 6'h1 == _T_752 ? _T_21 : _T_20; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6338 = 6'h2 == _T_752 ? _T_22 : _GEN_6337; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6339 = 6'h3 == _T_752 ? _T_23 : _GEN_6338; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6340 = 6'h4 == _T_752 ? _T_24 : _GEN_6339; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6341 = 6'h5 == _T_752 ? _T_25 : _GEN_6340; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6342 = 6'h6 == _T_752 ? _T_26 : _GEN_6341; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6343 = 6'h7 == _T_752 ? _T_27 : _GEN_6342; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6344 = 6'h8 == _T_752 ? _T_28 : _GEN_6343; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6345 = 6'h9 == _T_752 ? _T_29 : _GEN_6344; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6346 = 6'ha == _T_752 ? _T_30 : _GEN_6345; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6347 = 6'hb == _T_752 ? _T_31 : _GEN_6346; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6348 = 6'hc == _T_752 ? _T_32 : _GEN_6347; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6349 = 6'hd == _T_752 ? _T_33 : _GEN_6348; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6350 = 6'he == _T_752 ? _T_34 : _GEN_6349; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6351 = 6'hf == _T_752 ? _T_35 : _GEN_6350; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6352 = 6'h10 == _T_752 ? _T_36 : _GEN_6351; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6353 = 6'h11 == _T_752 ? _T_37 : _GEN_6352; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6354 = 6'h12 == _T_752 ? _T_38 : _GEN_6353; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6355 = 6'h13 == _T_752 ? _T_39 : _GEN_6354; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6356 = 6'h14 == _T_752 ? _T_40 : _GEN_6355; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6357 = 6'h15 == _T_752 ? _T_41 : _GEN_6356; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6358 = 6'h16 == _T_752 ? _T_42 : _GEN_6357; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6359 = 6'h17 == _T_752 ? _T_43 : _GEN_6358; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6360 = 6'h18 == _T_752 ? _T_44 : _GEN_6359; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6361 = 6'h19 == _T_752 ? _T_45 : _GEN_6360; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6362 = 6'h1a == _T_752 ? _T_46 : _GEN_6361; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6363 = 6'h1b == _T_752 ? _T_47 : _GEN_6362; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6364 = 6'h1c == _T_752 ? _T_48 : _GEN_6363; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6365 = 6'h1d == _T_752 ? _T_49 : _GEN_6364; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6366 = 6'h1e == _T_752 ? _T_50 : _GEN_6365; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6367 = 6'h1f == _T_752 ? _T_51 : _GEN_6366; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6368 = 6'h20 == _T_752 ? _T_52 : _GEN_6367; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6369 = 6'h21 == _T_752 ? _T_53 : _GEN_6368; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6370 = 6'h22 == _T_752 ? _T_54 : _GEN_6369; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6371 = 6'h23 == _T_752 ? _T_55 : _GEN_6370; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6372 = 6'h24 == _T_752 ? _T_56 : _GEN_6371; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6373 = 6'h25 == _T_752 ? _T_57 : _GEN_6372; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6374 = 6'h26 == _T_752 ? _T_58 : _GEN_6373; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6375 = 6'h27 == _T_752 ? _T_59 : _GEN_6374; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6376 = 6'h28 == _T_752 ? _T_60 : _GEN_6375; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6377 = 6'h29 == _T_752 ? _T_61 : _GEN_6376; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6378 = 6'h2a == _T_752 ? _T_62 : _GEN_6377; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6379 = 6'h2b == _T_752 ? _T_63 : _GEN_6378; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6380 = 6'h2c == _T_752 ? _T_64 : _GEN_6379; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6381 = 6'h2d == _T_752 ? _T_65 : _GEN_6380; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6382 = 6'h2e == _T_752 ? _T_66 : _GEN_6381; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6383 = 6'h2f == _T_752 ? _T_67 : _GEN_6382; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6384 = 6'h30 == _T_752 ? _T_68 : _GEN_6383; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6385 = 6'h31 == _T_752 ? _T_69 : _GEN_6384; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6386 = 6'h32 == _T_752 ? _T_70 : _GEN_6385; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6387 = 6'h33 == _T_752 ? _T_71 : _GEN_6386; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6388 = 6'h34 == _T_752 ? _T_72 : _GEN_6387; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6389 = 6'h35 == _T_752 ? _T_73 : _GEN_6388; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6390 = 6'h36 == _T_752 ? _T_74 : _GEN_6389; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6391 = 6'h37 == _T_752 ? _T_75 : _GEN_6390; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6392 = 6'h38 == _T_752 ? _T_76 : _GEN_6391; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6393 = 6'h39 == _T_752 ? _T_77 : _GEN_6392; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6394 = 6'h3a == _T_752 ? _T_78 : _GEN_6393; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6395 = 6'h3b == _T_752 ? _T_79 : _GEN_6394; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6396 = 6'h3c == _T_752 ? _T_80 : _GEN_6395; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6397 = 6'h3d == _T_752 ? _T_81 : _GEN_6396; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6398 = 6'h3e == _T_752 ? _T_82 : _GEN_6397; // @[execute.scala 79:10:@2200.4]
  assign _GEN_6399 = 6'h3f == _T_752 ? _T_83 : _GEN_6398; // @[execute.scala 79:10:@2200.4]
  assign _T_754 = _T_744 ? _GEN_6335 : _GEN_6399; // @[execute.scala 79:10:@2200.4]
  assign _T_756 = io_amount < 6'he; // @[execute.scala 79:15:@2201.4]
  assign _T_758 = io_amount - 6'he; // @[execute.scala 79:37:@2202.4]
  assign _T_759 = $unsigned(_T_758); // @[execute.scala 79:37:@2203.4]
  assign _T_760 = _T_759[5:0]; // @[execute.scala 79:37:@2204.4]
  assign _T_763 = 6'h32 + io_amount; // @[execute.scala 79:60:@2205.4]
  assign _T_764 = 6'h32 + io_amount; // @[execute.scala 79:60:@2206.4]
  assign _GEN_6401 = 6'h1 == _T_760 ? _T_21 : _T_20; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6402 = 6'h2 == _T_760 ? _T_22 : _GEN_6401; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6403 = 6'h3 == _T_760 ? _T_23 : _GEN_6402; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6404 = 6'h4 == _T_760 ? _T_24 : _GEN_6403; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6405 = 6'h5 == _T_760 ? _T_25 : _GEN_6404; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6406 = 6'h6 == _T_760 ? _T_26 : _GEN_6405; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6407 = 6'h7 == _T_760 ? _T_27 : _GEN_6406; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6408 = 6'h8 == _T_760 ? _T_28 : _GEN_6407; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6409 = 6'h9 == _T_760 ? _T_29 : _GEN_6408; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6410 = 6'ha == _T_760 ? _T_30 : _GEN_6409; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6411 = 6'hb == _T_760 ? _T_31 : _GEN_6410; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6412 = 6'hc == _T_760 ? _T_32 : _GEN_6411; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6413 = 6'hd == _T_760 ? _T_33 : _GEN_6412; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6414 = 6'he == _T_760 ? _T_34 : _GEN_6413; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6415 = 6'hf == _T_760 ? _T_35 : _GEN_6414; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6416 = 6'h10 == _T_760 ? _T_36 : _GEN_6415; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6417 = 6'h11 == _T_760 ? _T_37 : _GEN_6416; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6418 = 6'h12 == _T_760 ? _T_38 : _GEN_6417; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6419 = 6'h13 == _T_760 ? _T_39 : _GEN_6418; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6420 = 6'h14 == _T_760 ? _T_40 : _GEN_6419; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6421 = 6'h15 == _T_760 ? _T_41 : _GEN_6420; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6422 = 6'h16 == _T_760 ? _T_42 : _GEN_6421; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6423 = 6'h17 == _T_760 ? _T_43 : _GEN_6422; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6424 = 6'h18 == _T_760 ? _T_44 : _GEN_6423; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6425 = 6'h19 == _T_760 ? _T_45 : _GEN_6424; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6426 = 6'h1a == _T_760 ? _T_46 : _GEN_6425; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6427 = 6'h1b == _T_760 ? _T_47 : _GEN_6426; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6428 = 6'h1c == _T_760 ? _T_48 : _GEN_6427; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6429 = 6'h1d == _T_760 ? _T_49 : _GEN_6428; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6430 = 6'h1e == _T_760 ? _T_50 : _GEN_6429; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6431 = 6'h1f == _T_760 ? _T_51 : _GEN_6430; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6432 = 6'h20 == _T_760 ? _T_52 : _GEN_6431; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6433 = 6'h21 == _T_760 ? _T_53 : _GEN_6432; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6434 = 6'h22 == _T_760 ? _T_54 : _GEN_6433; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6435 = 6'h23 == _T_760 ? _T_55 : _GEN_6434; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6436 = 6'h24 == _T_760 ? _T_56 : _GEN_6435; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6437 = 6'h25 == _T_760 ? _T_57 : _GEN_6436; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6438 = 6'h26 == _T_760 ? _T_58 : _GEN_6437; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6439 = 6'h27 == _T_760 ? _T_59 : _GEN_6438; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6440 = 6'h28 == _T_760 ? _T_60 : _GEN_6439; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6441 = 6'h29 == _T_760 ? _T_61 : _GEN_6440; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6442 = 6'h2a == _T_760 ? _T_62 : _GEN_6441; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6443 = 6'h2b == _T_760 ? _T_63 : _GEN_6442; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6444 = 6'h2c == _T_760 ? _T_64 : _GEN_6443; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6445 = 6'h2d == _T_760 ? _T_65 : _GEN_6444; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6446 = 6'h2e == _T_760 ? _T_66 : _GEN_6445; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6447 = 6'h2f == _T_760 ? _T_67 : _GEN_6446; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6448 = 6'h30 == _T_760 ? _T_68 : _GEN_6447; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6449 = 6'h31 == _T_760 ? _T_69 : _GEN_6448; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6450 = 6'h32 == _T_760 ? _T_70 : _GEN_6449; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6451 = 6'h33 == _T_760 ? _T_71 : _GEN_6450; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6452 = 6'h34 == _T_760 ? _T_72 : _GEN_6451; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6453 = 6'h35 == _T_760 ? _T_73 : _GEN_6452; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6454 = 6'h36 == _T_760 ? _T_74 : _GEN_6453; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6455 = 6'h37 == _T_760 ? _T_75 : _GEN_6454; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6456 = 6'h38 == _T_760 ? _T_76 : _GEN_6455; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6457 = 6'h39 == _T_760 ? _T_77 : _GEN_6456; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6458 = 6'h3a == _T_760 ? _T_78 : _GEN_6457; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6459 = 6'h3b == _T_760 ? _T_79 : _GEN_6458; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6460 = 6'h3c == _T_760 ? _T_80 : _GEN_6459; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6461 = 6'h3d == _T_760 ? _T_81 : _GEN_6460; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6462 = 6'h3e == _T_760 ? _T_82 : _GEN_6461; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6463 = 6'h3f == _T_760 ? _T_83 : _GEN_6462; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6465 = 6'h1 == _T_764 ? _T_21 : _T_20; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6466 = 6'h2 == _T_764 ? _T_22 : _GEN_6465; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6467 = 6'h3 == _T_764 ? _T_23 : _GEN_6466; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6468 = 6'h4 == _T_764 ? _T_24 : _GEN_6467; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6469 = 6'h5 == _T_764 ? _T_25 : _GEN_6468; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6470 = 6'h6 == _T_764 ? _T_26 : _GEN_6469; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6471 = 6'h7 == _T_764 ? _T_27 : _GEN_6470; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6472 = 6'h8 == _T_764 ? _T_28 : _GEN_6471; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6473 = 6'h9 == _T_764 ? _T_29 : _GEN_6472; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6474 = 6'ha == _T_764 ? _T_30 : _GEN_6473; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6475 = 6'hb == _T_764 ? _T_31 : _GEN_6474; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6476 = 6'hc == _T_764 ? _T_32 : _GEN_6475; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6477 = 6'hd == _T_764 ? _T_33 : _GEN_6476; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6478 = 6'he == _T_764 ? _T_34 : _GEN_6477; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6479 = 6'hf == _T_764 ? _T_35 : _GEN_6478; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6480 = 6'h10 == _T_764 ? _T_36 : _GEN_6479; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6481 = 6'h11 == _T_764 ? _T_37 : _GEN_6480; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6482 = 6'h12 == _T_764 ? _T_38 : _GEN_6481; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6483 = 6'h13 == _T_764 ? _T_39 : _GEN_6482; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6484 = 6'h14 == _T_764 ? _T_40 : _GEN_6483; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6485 = 6'h15 == _T_764 ? _T_41 : _GEN_6484; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6486 = 6'h16 == _T_764 ? _T_42 : _GEN_6485; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6487 = 6'h17 == _T_764 ? _T_43 : _GEN_6486; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6488 = 6'h18 == _T_764 ? _T_44 : _GEN_6487; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6489 = 6'h19 == _T_764 ? _T_45 : _GEN_6488; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6490 = 6'h1a == _T_764 ? _T_46 : _GEN_6489; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6491 = 6'h1b == _T_764 ? _T_47 : _GEN_6490; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6492 = 6'h1c == _T_764 ? _T_48 : _GEN_6491; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6493 = 6'h1d == _T_764 ? _T_49 : _GEN_6492; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6494 = 6'h1e == _T_764 ? _T_50 : _GEN_6493; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6495 = 6'h1f == _T_764 ? _T_51 : _GEN_6494; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6496 = 6'h20 == _T_764 ? _T_52 : _GEN_6495; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6497 = 6'h21 == _T_764 ? _T_53 : _GEN_6496; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6498 = 6'h22 == _T_764 ? _T_54 : _GEN_6497; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6499 = 6'h23 == _T_764 ? _T_55 : _GEN_6498; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6500 = 6'h24 == _T_764 ? _T_56 : _GEN_6499; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6501 = 6'h25 == _T_764 ? _T_57 : _GEN_6500; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6502 = 6'h26 == _T_764 ? _T_58 : _GEN_6501; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6503 = 6'h27 == _T_764 ? _T_59 : _GEN_6502; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6504 = 6'h28 == _T_764 ? _T_60 : _GEN_6503; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6505 = 6'h29 == _T_764 ? _T_61 : _GEN_6504; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6506 = 6'h2a == _T_764 ? _T_62 : _GEN_6505; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6507 = 6'h2b == _T_764 ? _T_63 : _GEN_6506; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6508 = 6'h2c == _T_764 ? _T_64 : _GEN_6507; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6509 = 6'h2d == _T_764 ? _T_65 : _GEN_6508; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6510 = 6'h2e == _T_764 ? _T_66 : _GEN_6509; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6511 = 6'h2f == _T_764 ? _T_67 : _GEN_6510; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6512 = 6'h30 == _T_764 ? _T_68 : _GEN_6511; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6513 = 6'h31 == _T_764 ? _T_69 : _GEN_6512; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6514 = 6'h32 == _T_764 ? _T_70 : _GEN_6513; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6515 = 6'h33 == _T_764 ? _T_71 : _GEN_6514; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6516 = 6'h34 == _T_764 ? _T_72 : _GEN_6515; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6517 = 6'h35 == _T_764 ? _T_73 : _GEN_6516; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6518 = 6'h36 == _T_764 ? _T_74 : _GEN_6517; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6519 = 6'h37 == _T_764 ? _T_75 : _GEN_6518; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6520 = 6'h38 == _T_764 ? _T_76 : _GEN_6519; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6521 = 6'h39 == _T_764 ? _T_77 : _GEN_6520; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6522 = 6'h3a == _T_764 ? _T_78 : _GEN_6521; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6523 = 6'h3b == _T_764 ? _T_79 : _GEN_6522; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6524 = 6'h3c == _T_764 ? _T_80 : _GEN_6523; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6525 = 6'h3d == _T_764 ? _T_81 : _GEN_6524; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6526 = 6'h3e == _T_764 ? _T_82 : _GEN_6525; // @[execute.scala 79:10:@2207.4]
  assign _GEN_6527 = 6'h3f == _T_764 ? _T_83 : _GEN_6526; // @[execute.scala 79:10:@2207.4]
  assign _T_766 = _T_756 ? _GEN_6463 : _GEN_6527; // @[execute.scala 79:10:@2207.4]
  assign _T_768 = io_amount < 6'hd; // @[execute.scala 79:15:@2208.4]
  assign _T_770 = io_amount - 6'hd; // @[execute.scala 79:37:@2209.4]
  assign _T_771 = $unsigned(_T_770); // @[execute.scala 79:37:@2210.4]
  assign _T_772 = _T_771[5:0]; // @[execute.scala 79:37:@2211.4]
  assign _T_775 = 6'h33 + io_amount; // @[execute.scala 79:60:@2212.4]
  assign _T_776 = 6'h33 + io_amount; // @[execute.scala 79:60:@2213.4]
  assign _GEN_6529 = 6'h1 == _T_772 ? _T_21 : _T_20; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6530 = 6'h2 == _T_772 ? _T_22 : _GEN_6529; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6531 = 6'h3 == _T_772 ? _T_23 : _GEN_6530; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6532 = 6'h4 == _T_772 ? _T_24 : _GEN_6531; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6533 = 6'h5 == _T_772 ? _T_25 : _GEN_6532; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6534 = 6'h6 == _T_772 ? _T_26 : _GEN_6533; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6535 = 6'h7 == _T_772 ? _T_27 : _GEN_6534; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6536 = 6'h8 == _T_772 ? _T_28 : _GEN_6535; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6537 = 6'h9 == _T_772 ? _T_29 : _GEN_6536; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6538 = 6'ha == _T_772 ? _T_30 : _GEN_6537; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6539 = 6'hb == _T_772 ? _T_31 : _GEN_6538; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6540 = 6'hc == _T_772 ? _T_32 : _GEN_6539; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6541 = 6'hd == _T_772 ? _T_33 : _GEN_6540; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6542 = 6'he == _T_772 ? _T_34 : _GEN_6541; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6543 = 6'hf == _T_772 ? _T_35 : _GEN_6542; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6544 = 6'h10 == _T_772 ? _T_36 : _GEN_6543; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6545 = 6'h11 == _T_772 ? _T_37 : _GEN_6544; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6546 = 6'h12 == _T_772 ? _T_38 : _GEN_6545; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6547 = 6'h13 == _T_772 ? _T_39 : _GEN_6546; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6548 = 6'h14 == _T_772 ? _T_40 : _GEN_6547; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6549 = 6'h15 == _T_772 ? _T_41 : _GEN_6548; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6550 = 6'h16 == _T_772 ? _T_42 : _GEN_6549; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6551 = 6'h17 == _T_772 ? _T_43 : _GEN_6550; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6552 = 6'h18 == _T_772 ? _T_44 : _GEN_6551; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6553 = 6'h19 == _T_772 ? _T_45 : _GEN_6552; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6554 = 6'h1a == _T_772 ? _T_46 : _GEN_6553; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6555 = 6'h1b == _T_772 ? _T_47 : _GEN_6554; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6556 = 6'h1c == _T_772 ? _T_48 : _GEN_6555; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6557 = 6'h1d == _T_772 ? _T_49 : _GEN_6556; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6558 = 6'h1e == _T_772 ? _T_50 : _GEN_6557; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6559 = 6'h1f == _T_772 ? _T_51 : _GEN_6558; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6560 = 6'h20 == _T_772 ? _T_52 : _GEN_6559; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6561 = 6'h21 == _T_772 ? _T_53 : _GEN_6560; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6562 = 6'h22 == _T_772 ? _T_54 : _GEN_6561; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6563 = 6'h23 == _T_772 ? _T_55 : _GEN_6562; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6564 = 6'h24 == _T_772 ? _T_56 : _GEN_6563; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6565 = 6'h25 == _T_772 ? _T_57 : _GEN_6564; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6566 = 6'h26 == _T_772 ? _T_58 : _GEN_6565; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6567 = 6'h27 == _T_772 ? _T_59 : _GEN_6566; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6568 = 6'h28 == _T_772 ? _T_60 : _GEN_6567; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6569 = 6'h29 == _T_772 ? _T_61 : _GEN_6568; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6570 = 6'h2a == _T_772 ? _T_62 : _GEN_6569; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6571 = 6'h2b == _T_772 ? _T_63 : _GEN_6570; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6572 = 6'h2c == _T_772 ? _T_64 : _GEN_6571; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6573 = 6'h2d == _T_772 ? _T_65 : _GEN_6572; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6574 = 6'h2e == _T_772 ? _T_66 : _GEN_6573; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6575 = 6'h2f == _T_772 ? _T_67 : _GEN_6574; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6576 = 6'h30 == _T_772 ? _T_68 : _GEN_6575; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6577 = 6'h31 == _T_772 ? _T_69 : _GEN_6576; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6578 = 6'h32 == _T_772 ? _T_70 : _GEN_6577; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6579 = 6'h33 == _T_772 ? _T_71 : _GEN_6578; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6580 = 6'h34 == _T_772 ? _T_72 : _GEN_6579; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6581 = 6'h35 == _T_772 ? _T_73 : _GEN_6580; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6582 = 6'h36 == _T_772 ? _T_74 : _GEN_6581; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6583 = 6'h37 == _T_772 ? _T_75 : _GEN_6582; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6584 = 6'h38 == _T_772 ? _T_76 : _GEN_6583; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6585 = 6'h39 == _T_772 ? _T_77 : _GEN_6584; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6586 = 6'h3a == _T_772 ? _T_78 : _GEN_6585; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6587 = 6'h3b == _T_772 ? _T_79 : _GEN_6586; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6588 = 6'h3c == _T_772 ? _T_80 : _GEN_6587; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6589 = 6'h3d == _T_772 ? _T_81 : _GEN_6588; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6590 = 6'h3e == _T_772 ? _T_82 : _GEN_6589; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6591 = 6'h3f == _T_772 ? _T_83 : _GEN_6590; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6593 = 6'h1 == _T_776 ? _T_21 : _T_20; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6594 = 6'h2 == _T_776 ? _T_22 : _GEN_6593; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6595 = 6'h3 == _T_776 ? _T_23 : _GEN_6594; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6596 = 6'h4 == _T_776 ? _T_24 : _GEN_6595; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6597 = 6'h5 == _T_776 ? _T_25 : _GEN_6596; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6598 = 6'h6 == _T_776 ? _T_26 : _GEN_6597; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6599 = 6'h7 == _T_776 ? _T_27 : _GEN_6598; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6600 = 6'h8 == _T_776 ? _T_28 : _GEN_6599; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6601 = 6'h9 == _T_776 ? _T_29 : _GEN_6600; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6602 = 6'ha == _T_776 ? _T_30 : _GEN_6601; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6603 = 6'hb == _T_776 ? _T_31 : _GEN_6602; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6604 = 6'hc == _T_776 ? _T_32 : _GEN_6603; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6605 = 6'hd == _T_776 ? _T_33 : _GEN_6604; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6606 = 6'he == _T_776 ? _T_34 : _GEN_6605; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6607 = 6'hf == _T_776 ? _T_35 : _GEN_6606; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6608 = 6'h10 == _T_776 ? _T_36 : _GEN_6607; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6609 = 6'h11 == _T_776 ? _T_37 : _GEN_6608; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6610 = 6'h12 == _T_776 ? _T_38 : _GEN_6609; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6611 = 6'h13 == _T_776 ? _T_39 : _GEN_6610; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6612 = 6'h14 == _T_776 ? _T_40 : _GEN_6611; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6613 = 6'h15 == _T_776 ? _T_41 : _GEN_6612; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6614 = 6'h16 == _T_776 ? _T_42 : _GEN_6613; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6615 = 6'h17 == _T_776 ? _T_43 : _GEN_6614; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6616 = 6'h18 == _T_776 ? _T_44 : _GEN_6615; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6617 = 6'h19 == _T_776 ? _T_45 : _GEN_6616; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6618 = 6'h1a == _T_776 ? _T_46 : _GEN_6617; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6619 = 6'h1b == _T_776 ? _T_47 : _GEN_6618; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6620 = 6'h1c == _T_776 ? _T_48 : _GEN_6619; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6621 = 6'h1d == _T_776 ? _T_49 : _GEN_6620; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6622 = 6'h1e == _T_776 ? _T_50 : _GEN_6621; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6623 = 6'h1f == _T_776 ? _T_51 : _GEN_6622; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6624 = 6'h20 == _T_776 ? _T_52 : _GEN_6623; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6625 = 6'h21 == _T_776 ? _T_53 : _GEN_6624; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6626 = 6'h22 == _T_776 ? _T_54 : _GEN_6625; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6627 = 6'h23 == _T_776 ? _T_55 : _GEN_6626; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6628 = 6'h24 == _T_776 ? _T_56 : _GEN_6627; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6629 = 6'h25 == _T_776 ? _T_57 : _GEN_6628; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6630 = 6'h26 == _T_776 ? _T_58 : _GEN_6629; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6631 = 6'h27 == _T_776 ? _T_59 : _GEN_6630; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6632 = 6'h28 == _T_776 ? _T_60 : _GEN_6631; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6633 = 6'h29 == _T_776 ? _T_61 : _GEN_6632; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6634 = 6'h2a == _T_776 ? _T_62 : _GEN_6633; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6635 = 6'h2b == _T_776 ? _T_63 : _GEN_6634; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6636 = 6'h2c == _T_776 ? _T_64 : _GEN_6635; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6637 = 6'h2d == _T_776 ? _T_65 : _GEN_6636; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6638 = 6'h2e == _T_776 ? _T_66 : _GEN_6637; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6639 = 6'h2f == _T_776 ? _T_67 : _GEN_6638; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6640 = 6'h30 == _T_776 ? _T_68 : _GEN_6639; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6641 = 6'h31 == _T_776 ? _T_69 : _GEN_6640; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6642 = 6'h32 == _T_776 ? _T_70 : _GEN_6641; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6643 = 6'h33 == _T_776 ? _T_71 : _GEN_6642; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6644 = 6'h34 == _T_776 ? _T_72 : _GEN_6643; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6645 = 6'h35 == _T_776 ? _T_73 : _GEN_6644; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6646 = 6'h36 == _T_776 ? _T_74 : _GEN_6645; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6647 = 6'h37 == _T_776 ? _T_75 : _GEN_6646; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6648 = 6'h38 == _T_776 ? _T_76 : _GEN_6647; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6649 = 6'h39 == _T_776 ? _T_77 : _GEN_6648; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6650 = 6'h3a == _T_776 ? _T_78 : _GEN_6649; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6651 = 6'h3b == _T_776 ? _T_79 : _GEN_6650; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6652 = 6'h3c == _T_776 ? _T_80 : _GEN_6651; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6653 = 6'h3d == _T_776 ? _T_81 : _GEN_6652; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6654 = 6'h3e == _T_776 ? _T_82 : _GEN_6653; // @[execute.scala 79:10:@2214.4]
  assign _GEN_6655 = 6'h3f == _T_776 ? _T_83 : _GEN_6654; // @[execute.scala 79:10:@2214.4]
  assign _T_778 = _T_768 ? _GEN_6591 : _GEN_6655; // @[execute.scala 79:10:@2214.4]
  assign _T_780 = io_amount < 6'hc; // @[execute.scala 79:15:@2215.4]
  assign _T_782 = io_amount - 6'hc; // @[execute.scala 79:37:@2216.4]
  assign _T_783 = $unsigned(_T_782); // @[execute.scala 79:37:@2217.4]
  assign _T_784 = _T_783[5:0]; // @[execute.scala 79:37:@2218.4]
  assign _T_787 = 6'h34 + io_amount; // @[execute.scala 79:60:@2219.4]
  assign _T_788 = 6'h34 + io_amount; // @[execute.scala 79:60:@2220.4]
  assign _GEN_6657 = 6'h1 == _T_784 ? _T_21 : _T_20; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6658 = 6'h2 == _T_784 ? _T_22 : _GEN_6657; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6659 = 6'h3 == _T_784 ? _T_23 : _GEN_6658; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6660 = 6'h4 == _T_784 ? _T_24 : _GEN_6659; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6661 = 6'h5 == _T_784 ? _T_25 : _GEN_6660; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6662 = 6'h6 == _T_784 ? _T_26 : _GEN_6661; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6663 = 6'h7 == _T_784 ? _T_27 : _GEN_6662; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6664 = 6'h8 == _T_784 ? _T_28 : _GEN_6663; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6665 = 6'h9 == _T_784 ? _T_29 : _GEN_6664; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6666 = 6'ha == _T_784 ? _T_30 : _GEN_6665; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6667 = 6'hb == _T_784 ? _T_31 : _GEN_6666; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6668 = 6'hc == _T_784 ? _T_32 : _GEN_6667; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6669 = 6'hd == _T_784 ? _T_33 : _GEN_6668; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6670 = 6'he == _T_784 ? _T_34 : _GEN_6669; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6671 = 6'hf == _T_784 ? _T_35 : _GEN_6670; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6672 = 6'h10 == _T_784 ? _T_36 : _GEN_6671; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6673 = 6'h11 == _T_784 ? _T_37 : _GEN_6672; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6674 = 6'h12 == _T_784 ? _T_38 : _GEN_6673; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6675 = 6'h13 == _T_784 ? _T_39 : _GEN_6674; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6676 = 6'h14 == _T_784 ? _T_40 : _GEN_6675; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6677 = 6'h15 == _T_784 ? _T_41 : _GEN_6676; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6678 = 6'h16 == _T_784 ? _T_42 : _GEN_6677; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6679 = 6'h17 == _T_784 ? _T_43 : _GEN_6678; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6680 = 6'h18 == _T_784 ? _T_44 : _GEN_6679; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6681 = 6'h19 == _T_784 ? _T_45 : _GEN_6680; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6682 = 6'h1a == _T_784 ? _T_46 : _GEN_6681; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6683 = 6'h1b == _T_784 ? _T_47 : _GEN_6682; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6684 = 6'h1c == _T_784 ? _T_48 : _GEN_6683; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6685 = 6'h1d == _T_784 ? _T_49 : _GEN_6684; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6686 = 6'h1e == _T_784 ? _T_50 : _GEN_6685; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6687 = 6'h1f == _T_784 ? _T_51 : _GEN_6686; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6688 = 6'h20 == _T_784 ? _T_52 : _GEN_6687; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6689 = 6'h21 == _T_784 ? _T_53 : _GEN_6688; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6690 = 6'h22 == _T_784 ? _T_54 : _GEN_6689; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6691 = 6'h23 == _T_784 ? _T_55 : _GEN_6690; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6692 = 6'h24 == _T_784 ? _T_56 : _GEN_6691; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6693 = 6'h25 == _T_784 ? _T_57 : _GEN_6692; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6694 = 6'h26 == _T_784 ? _T_58 : _GEN_6693; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6695 = 6'h27 == _T_784 ? _T_59 : _GEN_6694; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6696 = 6'h28 == _T_784 ? _T_60 : _GEN_6695; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6697 = 6'h29 == _T_784 ? _T_61 : _GEN_6696; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6698 = 6'h2a == _T_784 ? _T_62 : _GEN_6697; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6699 = 6'h2b == _T_784 ? _T_63 : _GEN_6698; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6700 = 6'h2c == _T_784 ? _T_64 : _GEN_6699; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6701 = 6'h2d == _T_784 ? _T_65 : _GEN_6700; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6702 = 6'h2e == _T_784 ? _T_66 : _GEN_6701; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6703 = 6'h2f == _T_784 ? _T_67 : _GEN_6702; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6704 = 6'h30 == _T_784 ? _T_68 : _GEN_6703; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6705 = 6'h31 == _T_784 ? _T_69 : _GEN_6704; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6706 = 6'h32 == _T_784 ? _T_70 : _GEN_6705; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6707 = 6'h33 == _T_784 ? _T_71 : _GEN_6706; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6708 = 6'h34 == _T_784 ? _T_72 : _GEN_6707; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6709 = 6'h35 == _T_784 ? _T_73 : _GEN_6708; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6710 = 6'h36 == _T_784 ? _T_74 : _GEN_6709; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6711 = 6'h37 == _T_784 ? _T_75 : _GEN_6710; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6712 = 6'h38 == _T_784 ? _T_76 : _GEN_6711; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6713 = 6'h39 == _T_784 ? _T_77 : _GEN_6712; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6714 = 6'h3a == _T_784 ? _T_78 : _GEN_6713; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6715 = 6'h3b == _T_784 ? _T_79 : _GEN_6714; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6716 = 6'h3c == _T_784 ? _T_80 : _GEN_6715; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6717 = 6'h3d == _T_784 ? _T_81 : _GEN_6716; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6718 = 6'h3e == _T_784 ? _T_82 : _GEN_6717; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6719 = 6'h3f == _T_784 ? _T_83 : _GEN_6718; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6721 = 6'h1 == _T_788 ? _T_21 : _T_20; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6722 = 6'h2 == _T_788 ? _T_22 : _GEN_6721; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6723 = 6'h3 == _T_788 ? _T_23 : _GEN_6722; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6724 = 6'h4 == _T_788 ? _T_24 : _GEN_6723; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6725 = 6'h5 == _T_788 ? _T_25 : _GEN_6724; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6726 = 6'h6 == _T_788 ? _T_26 : _GEN_6725; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6727 = 6'h7 == _T_788 ? _T_27 : _GEN_6726; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6728 = 6'h8 == _T_788 ? _T_28 : _GEN_6727; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6729 = 6'h9 == _T_788 ? _T_29 : _GEN_6728; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6730 = 6'ha == _T_788 ? _T_30 : _GEN_6729; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6731 = 6'hb == _T_788 ? _T_31 : _GEN_6730; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6732 = 6'hc == _T_788 ? _T_32 : _GEN_6731; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6733 = 6'hd == _T_788 ? _T_33 : _GEN_6732; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6734 = 6'he == _T_788 ? _T_34 : _GEN_6733; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6735 = 6'hf == _T_788 ? _T_35 : _GEN_6734; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6736 = 6'h10 == _T_788 ? _T_36 : _GEN_6735; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6737 = 6'h11 == _T_788 ? _T_37 : _GEN_6736; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6738 = 6'h12 == _T_788 ? _T_38 : _GEN_6737; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6739 = 6'h13 == _T_788 ? _T_39 : _GEN_6738; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6740 = 6'h14 == _T_788 ? _T_40 : _GEN_6739; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6741 = 6'h15 == _T_788 ? _T_41 : _GEN_6740; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6742 = 6'h16 == _T_788 ? _T_42 : _GEN_6741; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6743 = 6'h17 == _T_788 ? _T_43 : _GEN_6742; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6744 = 6'h18 == _T_788 ? _T_44 : _GEN_6743; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6745 = 6'h19 == _T_788 ? _T_45 : _GEN_6744; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6746 = 6'h1a == _T_788 ? _T_46 : _GEN_6745; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6747 = 6'h1b == _T_788 ? _T_47 : _GEN_6746; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6748 = 6'h1c == _T_788 ? _T_48 : _GEN_6747; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6749 = 6'h1d == _T_788 ? _T_49 : _GEN_6748; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6750 = 6'h1e == _T_788 ? _T_50 : _GEN_6749; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6751 = 6'h1f == _T_788 ? _T_51 : _GEN_6750; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6752 = 6'h20 == _T_788 ? _T_52 : _GEN_6751; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6753 = 6'h21 == _T_788 ? _T_53 : _GEN_6752; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6754 = 6'h22 == _T_788 ? _T_54 : _GEN_6753; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6755 = 6'h23 == _T_788 ? _T_55 : _GEN_6754; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6756 = 6'h24 == _T_788 ? _T_56 : _GEN_6755; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6757 = 6'h25 == _T_788 ? _T_57 : _GEN_6756; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6758 = 6'h26 == _T_788 ? _T_58 : _GEN_6757; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6759 = 6'h27 == _T_788 ? _T_59 : _GEN_6758; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6760 = 6'h28 == _T_788 ? _T_60 : _GEN_6759; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6761 = 6'h29 == _T_788 ? _T_61 : _GEN_6760; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6762 = 6'h2a == _T_788 ? _T_62 : _GEN_6761; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6763 = 6'h2b == _T_788 ? _T_63 : _GEN_6762; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6764 = 6'h2c == _T_788 ? _T_64 : _GEN_6763; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6765 = 6'h2d == _T_788 ? _T_65 : _GEN_6764; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6766 = 6'h2e == _T_788 ? _T_66 : _GEN_6765; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6767 = 6'h2f == _T_788 ? _T_67 : _GEN_6766; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6768 = 6'h30 == _T_788 ? _T_68 : _GEN_6767; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6769 = 6'h31 == _T_788 ? _T_69 : _GEN_6768; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6770 = 6'h32 == _T_788 ? _T_70 : _GEN_6769; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6771 = 6'h33 == _T_788 ? _T_71 : _GEN_6770; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6772 = 6'h34 == _T_788 ? _T_72 : _GEN_6771; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6773 = 6'h35 == _T_788 ? _T_73 : _GEN_6772; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6774 = 6'h36 == _T_788 ? _T_74 : _GEN_6773; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6775 = 6'h37 == _T_788 ? _T_75 : _GEN_6774; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6776 = 6'h38 == _T_788 ? _T_76 : _GEN_6775; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6777 = 6'h39 == _T_788 ? _T_77 : _GEN_6776; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6778 = 6'h3a == _T_788 ? _T_78 : _GEN_6777; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6779 = 6'h3b == _T_788 ? _T_79 : _GEN_6778; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6780 = 6'h3c == _T_788 ? _T_80 : _GEN_6779; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6781 = 6'h3d == _T_788 ? _T_81 : _GEN_6780; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6782 = 6'h3e == _T_788 ? _T_82 : _GEN_6781; // @[execute.scala 79:10:@2221.4]
  assign _GEN_6783 = 6'h3f == _T_788 ? _T_83 : _GEN_6782; // @[execute.scala 79:10:@2221.4]
  assign _T_790 = _T_780 ? _GEN_6719 : _GEN_6783; // @[execute.scala 79:10:@2221.4]
  assign _T_792 = io_amount < 6'hb; // @[execute.scala 79:15:@2222.4]
  assign _T_794 = io_amount - 6'hb; // @[execute.scala 79:37:@2223.4]
  assign _T_795 = $unsigned(_T_794); // @[execute.scala 79:37:@2224.4]
  assign _T_796 = _T_795[5:0]; // @[execute.scala 79:37:@2225.4]
  assign _T_799 = 6'h35 + io_amount; // @[execute.scala 79:60:@2226.4]
  assign _T_800 = 6'h35 + io_amount; // @[execute.scala 79:60:@2227.4]
  assign _GEN_6785 = 6'h1 == _T_796 ? _T_21 : _T_20; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6786 = 6'h2 == _T_796 ? _T_22 : _GEN_6785; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6787 = 6'h3 == _T_796 ? _T_23 : _GEN_6786; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6788 = 6'h4 == _T_796 ? _T_24 : _GEN_6787; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6789 = 6'h5 == _T_796 ? _T_25 : _GEN_6788; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6790 = 6'h6 == _T_796 ? _T_26 : _GEN_6789; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6791 = 6'h7 == _T_796 ? _T_27 : _GEN_6790; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6792 = 6'h8 == _T_796 ? _T_28 : _GEN_6791; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6793 = 6'h9 == _T_796 ? _T_29 : _GEN_6792; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6794 = 6'ha == _T_796 ? _T_30 : _GEN_6793; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6795 = 6'hb == _T_796 ? _T_31 : _GEN_6794; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6796 = 6'hc == _T_796 ? _T_32 : _GEN_6795; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6797 = 6'hd == _T_796 ? _T_33 : _GEN_6796; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6798 = 6'he == _T_796 ? _T_34 : _GEN_6797; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6799 = 6'hf == _T_796 ? _T_35 : _GEN_6798; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6800 = 6'h10 == _T_796 ? _T_36 : _GEN_6799; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6801 = 6'h11 == _T_796 ? _T_37 : _GEN_6800; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6802 = 6'h12 == _T_796 ? _T_38 : _GEN_6801; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6803 = 6'h13 == _T_796 ? _T_39 : _GEN_6802; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6804 = 6'h14 == _T_796 ? _T_40 : _GEN_6803; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6805 = 6'h15 == _T_796 ? _T_41 : _GEN_6804; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6806 = 6'h16 == _T_796 ? _T_42 : _GEN_6805; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6807 = 6'h17 == _T_796 ? _T_43 : _GEN_6806; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6808 = 6'h18 == _T_796 ? _T_44 : _GEN_6807; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6809 = 6'h19 == _T_796 ? _T_45 : _GEN_6808; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6810 = 6'h1a == _T_796 ? _T_46 : _GEN_6809; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6811 = 6'h1b == _T_796 ? _T_47 : _GEN_6810; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6812 = 6'h1c == _T_796 ? _T_48 : _GEN_6811; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6813 = 6'h1d == _T_796 ? _T_49 : _GEN_6812; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6814 = 6'h1e == _T_796 ? _T_50 : _GEN_6813; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6815 = 6'h1f == _T_796 ? _T_51 : _GEN_6814; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6816 = 6'h20 == _T_796 ? _T_52 : _GEN_6815; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6817 = 6'h21 == _T_796 ? _T_53 : _GEN_6816; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6818 = 6'h22 == _T_796 ? _T_54 : _GEN_6817; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6819 = 6'h23 == _T_796 ? _T_55 : _GEN_6818; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6820 = 6'h24 == _T_796 ? _T_56 : _GEN_6819; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6821 = 6'h25 == _T_796 ? _T_57 : _GEN_6820; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6822 = 6'h26 == _T_796 ? _T_58 : _GEN_6821; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6823 = 6'h27 == _T_796 ? _T_59 : _GEN_6822; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6824 = 6'h28 == _T_796 ? _T_60 : _GEN_6823; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6825 = 6'h29 == _T_796 ? _T_61 : _GEN_6824; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6826 = 6'h2a == _T_796 ? _T_62 : _GEN_6825; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6827 = 6'h2b == _T_796 ? _T_63 : _GEN_6826; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6828 = 6'h2c == _T_796 ? _T_64 : _GEN_6827; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6829 = 6'h2d == _T_796 ? _T_65 : _GEN_6828; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6830 = 6'h2e == _T_796 ? _T_66 : _GEN_6829; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6831 = 6'h2f == _T_796 ? _T_67 : _GEN_6830; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6832 = 6'h30 == _T_796 ? _T_68 : _GEN_6831; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6833 = 6'h31 == _T_796 ? _T_69 : _GEN_6832; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6834 = 6'h32 == _T_796 ? _T_70 : _GEN_6833; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6835 = 6'h33 == _T_796 ? _T_71 : _GEN_6834; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6836 = 6'h34 == _T_796 ? _T_72 : _GEN_6835; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6837 = 6'h35 == _T_796 ? _T_73 : _GEN_6836; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6838 = 6'h36 == _T_796 ? _T_74 : _GEN_6837; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6839 = 6'h37 == _T_796 ? _T_75 : _GEN_6838; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6840 = 6'h38 == _T_796 ? _T_76 : _GEN_6839; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6841 = 6'h39 == _T_796 ? _T_77 : _GEN_6840; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6842 = 6'h3a == _T_796 ? _T_78 : _GEN_6841; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6843 = 6'h3b == _T_796 ? _T_79 : _GEN_6842; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6844 = 6'h3c == _T_796 ? _T_80 : _GEN_6843; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6845 = 6'h3d == _T_796 ? _T_81 : _GEN_6844; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6846 = 6'h3e == _T_796 ? _T_82 : _GEN_6845; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6847 = 6'h3f == _T_796 ? _T_83 : _GEN_6846; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6849 = 6'h1 == _T_800 ? _T_21 : _T_20; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6850 = 6'h2 == _T_800 ? _T_22 : _GEN_6849; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6851 = 6'h3 == _T_800 ? _T_23 : _GEN_6850; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6852 = 6'h4 == _T_800 ? _T_24 : _GEN_6851; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6853 = 6'h5 == _T_800 ? _T_25 : _GEN_6852; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6854 = 6'h6 == _T_800 ? _T_26 : _GEN_6853; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6855 = 6'h7 == _T_800 ? _T_27 : _GEN_6854; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6856 = 6'h8 == _T_800 ? _T_28 : _GEN_6855; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6857 = 6'h9 == _T_800 ? _T_29 : _GEN_6856; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6858 = 6'ha == _T_800 ? _T_30 : _GEN_6857; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6859 = 6'hb == _T_800 ? _T_31 : _GEN_6858; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6860 = 6'hc == _T_800 ? _T_32 : _GEN_6859; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6861 = 6'hd == _T_800 ? _T_33 : _GEN_6860; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6862 = 6'he == _T_800 ? _T_34 : _GEN_6861; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6863 = 6'hf == _T_800 ? _T_35 : _GEN_6862; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6864 = 6'h10 == _T_800 ? _T_36 : _GEN_6863; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6865 = 6'h11 == _T_800 ? _T_37 : _GEN_6864; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6866 = 6'h12 == _T_800 ? _T_38 : _GEN_6865; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6867 = 6'h13 == _T_800 ? _T_39 : _GEN_6866; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6868 = 6'h14 == _T_800 ? _T_40 : _GEN_6867; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6869 = 6'h15 == _T_800 ? _T_41 : _GEN_6868; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6870 = 6'h16 == _T_800 ? _T_42 : _GEN_6869; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6871 = 6'h17 == _T_800 ? _T_43 : _GEN_6870; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6872 = 6'h18 == _T_800 ? _T_44 : _GEN_6871; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6873 = 6'h19 == _T_800 ? _T_45 : _GEN_6872; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6874 = 6'h1a == _T_800 ? _T_46 : _GEN_6873; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6875 = 6'h1b == _T_800 ? _T_47 : _GEN_6874; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6876 = 6'h1c == _T_800 ? _T_48 : _GEN_6875; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6877 = 6'h1d == _T_800 ? _T_49 : _GEN_6876; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6878 = 6'h1e == _T_800 ? _T_50 : _GEN_6877; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6879 = 6'h1f == _T_800 ? _T_51 : _GEN_6878; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6880 = 6'h20 == _T_800 ? _T_52 : _GEN_6879; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6881 = 6'h21 == _T_800 ? _T_53 : _GEN_6880; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6882 = 6'h22 == _T_800 ? _T_54 : _GEN_6881; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6883 = 6'h23 == _T_800 ? _T_55 : _GEN_6882; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6884 = 6'h24 == _T_800 ? _T_56 : _GEN_6883; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6885 = 6'h25 == _T_800 ? _T_57 : _GEN_6884; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6886 = 6'h26 == _T_800 ? _T_58 : _GEN_6885; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6887 = 6'h27 == _T_800 ? _T_59 : _GEN_6886; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6888 = 6'h28 == _T_800 ? _T_60 : _GEN_6887; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6889 = 6'h29 == _T_800 ? _T_61 : _GEN_6888; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6890 = 6'h2a == _T_800 ? _T_62 : _GEN_6889; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6891 = 6'h2b == _T_800 ? _T_63 : _GEN_6890; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6892 = 6'h2c == _T_800 ? _T_64 : _GEN_6891; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6893 = 6'h2d == _T_800 ? _T_65 : _GEN_6892; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6894 = 6'h2e == _T_800 ? _T_66 : _GEN_6893; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6895 = 6'h2f == _T_800 ? _T_67 : _GEN_6894; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6896 = 6'h30 == _T_800 ? _T_68 : _GEN_6895; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6897 = 6'h31 == _T_800 ? _T_69 : _GEN_6896; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6898 = 6'h32 == _T_800 ? _T_70 : _GEN_6897; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6899 = 6'h33 == _T_800 ? _T_71 : _GEN_6898; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6900 = 6'h34 == _T_800 ? _T_72 : _GEN_6899; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6901 = 6'h35 == _T_800 ? _T_73 : _GEN_6900; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6902 = 6'h36 == _T_800 ? _T_74 : _GEN_6901; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6903 = 6'h37 == _T_800 ? _T_75 : _GEN_6902; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6904 = 6'h38 == _T_800 ? _T_76 : _GEN_6903; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6905 = 6'h39 == _T_800 ? _T_77 : _GEN_6904; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6906 = 6'h3a == _T_800 ? _T_78 : _GEN_6905; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6907 = 6'h3b == _T_800 ? _T_79 : _GEN_6906; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6908 = 6'h3c == _T_800 ? _T_80 : _GEN_6907; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6909 = 6'h3d == _T_800 ? _T_81 : _GEN_6908; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6910 = 6'h3e == _T_800 ? _T_82 : _GEN_6909; // @[execute.scala 79:10:@2228.4]
  assign _GEN_6911 = 6'h3f == _T_800 ? _T_83 : _GEN_6910; // @[execute.scala 79:10:@2228.4]
  assign _T_802 = _T_792 ? _GEN_6847 : _GEN_6911; // @[execute.scala 79:10:@2228.4]
  assign _T_804 = io_amount < 6'ha; // @[execute.scala 79:15:@2229.4]
  assign _T_806 = io_amount - 6'ha; // @[execute.scala 79:37:@2230.4]
  assign _T_807 = $unsigned(_T_806); // @[execute.scala 79:37:@2231.4]
  assign _T_808 = _T_807[5:0]; // @[execute.scala 79:37:@2232.4]
  assign _T_811 = 6'h36 + io_amount; // @[execute.scala 79:60:@2233.4]
  assign _T_812 = 6'h36 + io_amount; // @[execute.scala 79:60:@2234.4]
  assign _GEN_6913 = 6'h1 == _T_808 ? _T_21 : _T_20; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6914 = 6'h2 == _T_808 ? _T_22 : _GEN_6913; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6915 = 6'h3 == _T_808 ? _T_23 : _GEN_6914; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6916 = 6'h4 == _T_808 ? _T_24 : _GEN_6915; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6917 = 6'h5 == _T_808 ? _T_25 : _GEN_6916; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6918 = 6'h6 == _T_808 ? _T_26 : _GEN_6917; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6919 = 6'h7 == _T_808 ? _T_27 : _GEN_6918; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6920 = 6'h8 == _T_808 ? _T_28 : _GEN_6919; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6921 = 6'h9 == _T_808 ? _T_29 : _GEN_6920; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6922 = 6'ha == _T_808 ? _T_30 : _GEN_6921; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6923 = 6'hb == _T_808 ? _T_31 : _GEN_6922; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6924 = 6'hc == _T_808 ? _T_32 : _GEN_6923; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6925 = 6'hd == _T_808 ? _T_33 : _GEN_6924; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6926 = 6'he == _T_808 ? _T_34 : _GEN_6925; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6927 = 6'hf == _T_808 ? _T_35 : _GEN_6926; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6928 = 6'h10 == _T_808 ? _T_36 : _GEN_6927; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6929 = 6'h11 == _T_808 ? _T_37 : _GEN_6928; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6930 = 6'h12 == _T_808 ? _T_38 : _GEN_6929; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6931 = 6'h13 == _T_808 ? _T_39 : _GEN_6930; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6932 = 6'h14 == _T_808 ? _T_40 : _GEN_6931; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6933 = 6'h15 == _T_808 ? _T_41 : _GEN_6932; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6934 = 6'h16 == _T_808 ? _T_42 : _GEN_6933; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6935 = 6'h17 == _T_808 ? _T_43 : _GEN_6934; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6936 = 6'h18 == _T_808 ? _T_44 : _GEN_6935; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6937 = 6'h19 == _T_808 ? _T_45 : _GEN_6936; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6938 = 6'h1a == _T_808 ? _T_46 : _GEN_6937; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6939 = 6'h1b == _T_808 ? _T_47 : _GEN_6938; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6940 = 6'h1c == _T_808 ? _T_48 : _GEN_6939; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6941 = 6'h1d == _T_808 ? _T_49 : _GEN_6940; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6942 = 6'h1e == _T_808 ? _T_50 : _GEN_6941; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6943 = 6'h1f == _T_808 ? _T_51 : _GEN_6942; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6944 = 6'h20 == _T_808 ? _T_52 : _GEN_6943; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6945 = 6'h21 == _T_808 ? _T_53 : _GEN_6944; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6946 = 6'h22 == _T_808 ? _T_54 : _GEN_6945; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6947 = 6'h23 == _T_808 ? _T_55 : _GEN_6946; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6948 = 6'h24 == _T_808 ? _T_56 : _GEN_6947; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6949 = 6'h25 == _T_808 ? _T_57 : _GEN_6948; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6950 = 6'h26 == _T_808 ? _T_58 : _GEN_6949; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6951 = 6'h27 == _T_808 ? _T_59 : _GEN_6950; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6952 = 6'h28 == _T_808 ? _T_60 : _GEN_6951; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6953 = 6'h29 == _T_808 ? _T_61 : _GEN_6952; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6954 = 6'h2a == _T_808 ? _T_62 : _GEN_6953; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6955 = 6'h2b == _T_808 ? _T_63 : _GEN_6954; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6956 = 6'h2c == _T_808 ? _T_64 : _GEN_6955; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6957 = 6'h2d == _T_808 ? _T_65 : _GEN_6956; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6958 = 6'h2e == _T_808 ? _T_66 : _GEN_6957; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6959 = 6'h2f == _T_808 ? _T_67 : _GEN_6958; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6960 = 6'h30 == _T_808 ? _T_68 : _GEN_6959; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6961 = 6'h31 == _T_808 ? _T_69 : _GEN_6960; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6962 = 6'h32 == _T_808 ? _T_70 : _GEN_6961; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6963 = 6'h33 == _T_808 ? _T_71 : _GEN_6962; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6964 = 6'h34 == _T_808 ? _T_72 : _GEN_6963; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6965 = 6'h35 == _T_808 ? _T_73 : _GEN_6964; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6966 = 6'h36 == _T_808 ? _T_74 : _GEN_6965; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6967 = 6'h37 == _T_808 ? _T_75 : _GEN_6966; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6968 = 6'h38 == _T_808 ? _T_76 : _GEN_6967; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6969 = 6'h39 == _T_808 ? _T_77 : _GEN_6968; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6970 = 6'h3a == _T_808 ? _T_78 : _GEN_6969; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6971 = 6'h3b == _T_808 ? _T_79 : _GEN_6970; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6972 = 6'h3c == _T_808 ? _T_80 : _GEN_6971; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6973 = 6'h3d == _T_808 ? _T_81 : _GEN_6972; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6974 = 6'h3e == _T_808 ? _T_82 : _GEN_6973; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6975 = 6'h3f == _T_808 ? _T_83 : _GEN_6974; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6977 = 6'h1 == _T_812 ? _T_21 : _T_20; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6978 = 6'h2 == _T_812 ? _T_22 : _GEN_6977; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6979 = 6'h3 == _T_812 ? _T_23 : _GEN_6978; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6980 = 6'h4 == _T_812 ? _T_24 : _GEN_6979; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6981 = 6'h5 == _T_812 ? _T_25 : _GEN_6980; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6982 = 6'h6 == _T_812 ? _T_26 : _GEN_6981; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6983 = 6'h7 == _T_812 ? _T_27 : _GEN_6982; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6984 = 6'h8 == _T_812 ? _T_28 : _GEN_6983; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6985 = 6'h9 == _T_812 ? _T_29 : _GEN_6984; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6986 = 6'ha == _T_812 ? _T_30 : _GEN_6985; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6987 = 6'hb == _T_812 ? _T_31 : _GEN_6986; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6988 = 6'hc == _T_812 ? _T_32 : _GEN_6987; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6989 = 6'hd == _T_812 ? _T_33 : _GEN_6988; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6990 = 6'he == _T_812 ? _T_34 : _GEN_6989; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6991 = 6'hf == _T_812 ? _T_35 : _GEN_6990; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6992 = 6'h10 == _T_812 ? _T_36 : _GEN_6991; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6993 = 6'h11 == _T_812 ? _T_37 : _GEN_6992; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6994 = 6'h12 == _T_812 ? _T_38 : _GEN_6993; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6995 = 6'h13 == _T_812 ? _T_39 : _GEN_6994; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6996 = 6'h14 == _T_812 ? _T_40 : _GEN_6995; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6997 = 6'h15 == _T_812 ? _T_41 : _GEN_6996; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6998 = 6'h16 == _T_812 ? _T_42 : _GEN_6997; // @[execute.scala 79:10:@2235.4]
  assign _GEN_6999 = 6'h17 == _T_812 ? _T_43 : _GEN_6998; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7000 = 6'h18 == _T_812 ? _T_44 : _GEN_6999; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7001 = 6'h19 == _T_812 ? _T_45 : _GEN_7000; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7002 = 6'h1a == _T_812 ? _T_46 : _GEN_7001; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7003 = 6'h1b == _T_812 ? _T_47 : _GEN_7002; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7004 = 6'h1c == _T_812 ? _T_48 : _GEN_7003; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7005 = 6'h1d == _T_812 ? _T_49 : _GEN_7004; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7006 = 6'h1e == _T_812 ? _T_50 : _GEN_7005; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7007 = 6'h1f == _T_812 ? _T_51 : _GEN_7006; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7008 = 6'h20 == _T_812 ? _T_52 : _GEN_7007; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7009 = 6'h21 == _T_812 ? _T_53 : _GEN_7008; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7010 = 6'h22 == _T_812 ? _T_54 : _GEN_7009; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7011 = 6'h23 == _T_812 ? _T_55 : _GEN_7010; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7012 = 6'h24 == _T_812 ? _T_56 : _GEN_7011; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7013 = 6'h25 == _T_812 ? _T_57 : _GEN_7012; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7014 = 6'h26 == _T_812 ? _T_58 : _GEN_7013; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7015 = 6'h27 == _T_812 ? _T_59 : _GEN_7014; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7016 = 6'h28 == _T_812 ? _T_60 : _GEN_7015; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7017 = 6'h29 == _T_812 ? _T_61 : _GEN_7016; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7018 = 6'h2a == _T_812 ? _T_62 : _GEN_7017; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7019 = 6'h2b == _T_812 ? _T_63 : _GEN_7018; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7020 = 6'h2c == _T_812 ? _T_64 : _GEN_7019; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7021 = 6'h2d == _T_812 ? _T_65 : _GEN_7020; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7022 = 6'h2e == _T_812 ? _T_66 : _GEN_7021; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7023 = 6'h2f == _T_812 ? _T_67 : _GEN_7022; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7024 = 6'h30 == _T_812 ? _T_68 : _GEN_7023; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7025 = 6'h31 == _T_812 ? _T_69 : _GEN_7024; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7026 = 6'h32 == _T_812 ? _T_70 : _GEN_7025; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7027 = 6'h33 == _T_812 ? _T_71 : _GEN_7026; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7028 = 6'h34 == _T_812 ? _T_72 : _GEN_7027; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7029 = 6'h35 == _T_812 ? _T_73 : _GEN_7028; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7030 = 6'h36 == _T_812 ? _T_74 : _GEN_7029; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7031 = 6'h37 == _T_812 ? _T_75 : _GEN_7030; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7032 = 6'h38 == _T_812 ? _T_76 : _GEN_7031; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7033 = 6'h39 == _T_812 ? _T_77 : _GEN_7032; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7034 = 6'h3a == _T_812 ? _T_78 : _GEN_7033; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7035 = 6'h3b == _T_812 ? _T_79 : _GEN_7034; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7036 = 6'h3c == _T_812 ? _T_80 : _GEN_7035; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7037 = 6'h3d == _T_812 ? _T_81 : _GEN_7036; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7038 = 6'h3e == _T_812 ? _T_82 : _GEN_7037; // @[execute.scala 79:10:@2235.4]
  assign _GEN_7039 = 6'h3f == _T_812 ? _T_83 : _GEN_7038; // @[execute.scala 79:10:@2235.4]
  assign _T_814 = _T_804 ? _GEN_6975 : _GEN_7039; // @[execute.scala 79:10:@2235.4]
  assign _T_816 = io_amount < 6'h9; // @[execute.scala 79:15:@2236.4]
  assign _T_818 = io_amount - 6'h9; // @[execute.scala 79:37:@2237.4]
  assign _T_819 = $unsigned(_T_818); // @[execute.scala 79:37:@2238.4]
  assign _T_820 = _T_819[5:0]; // @[execute.scala 79:37:@2239.4]
  assign _T_823 = 6'h37 + io_amount; // @[execute.scala 79:60:@2240.4]
  assign _T_824 = 6'h37 + io_amount; // @[execute.scala 79:60:@2241.4]
  assign _GEN_7041 = 6'h1 == _T_820 ? _T_21 : _T_20; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7042 = 6'h2 == _T_820 ? _T_22 : _GEN_7041; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7043 = 6'h3 == _T_820 ? _T_23 : _GEN_7042; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7044 = 6'h4 == _T_820 ? _T_24 : _GEN_7043; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7045 = 6'h5 == _T_820 ? _T_25 : _GEN_7044; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7046 = 6'h6 == _T_820 ? _T_26 : _GEN_7045; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7047 = 6'h7 == _T_820 ? _T_27 : _GEN_7046; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7048 = 6'h8 == _T_820 ? _T_28 : _GEN_7047; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7049 = 6'h9 == _T_820 ? _T_29 : _GEN_7048; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7050 = 6'ha == _T_820 ? _T_30 : _GEN_7049; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7051 = 6'hb == _T_820 ? _T_31 : _GEN_7050; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7052 = 6'hc == _T_820 ? _T_32 : _GEN_7051; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7053 = 6'hd == _T_820 ? _T_33 : _GEN_7052; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7054 = 6'he == _T_820 ? _T_34 : _GEN_7053; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7055 = 6'hf == _T_820 ? _T_35 : _GEN_7054; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7056 = 6'h10 == _T_820 ? _T_36 : _GEN_7055; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7057 = 6'h11 == _T_820 ? _T_37 : _GEN_7056; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7058 = 6'h12 == _T_820 ? _T_38 : _GEN_7057; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7059 = 6'h13 == _T_820 ? _T_39 : _GEN_7058; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7060 = 6'h14 == _T_820 ? _T_40 : _GEN_7059; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7061 = 6'h15 == _T_820 ? _T_41 : _GEN_7060; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7062 = 6'h16 == _T_820 ? _T_42 : _GEN_7061; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7063 = 6'h17 == _T_820 ? _T_43 : _GEN_7062; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7064 = 6'h18 == _T_820 ? _T_44 : _GEN_7063; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7065 = 6'h19 == _T_820 ? _T_45 : _GEN_7064; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7066 = 6'h1a == _T_820 ? _T_46 : _GEN_7065; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7067 = 6'h1b == _T_820 ? _T_47 : _GEN_7066; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7068 = 6'h1c == _T_820 ? _T_48 : _GEN_7067; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7069 = 6'h1d == _T_820 ? _T_49 : _GEN_7068; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7070 = 6'h1e == _T_820 ? _T_50 : _GEN_7069; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7071 = 6'h1f == _T_820 ? _T_51 : _GEN_7070; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7072 = 6'h20 == _T_820 ? _T_52 : _GEN_7071; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7073 = 6'h21 == _T_820 ? _T_53 : _GEN_7072; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7074 = 6'h22 == _T_820 ? _T_54 : _GEN_7073; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7075 = 6'h23 == _T_820 ? _T_55 : _GEN_7074; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7076 = 6'h24 == _T_820 ? _T_56 : _GEN_7075; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7077 = 6'h25 == _T_820 ? _T_57 : _GEN_7076; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7078 = 6'h26 == _T_820 ? _T_58 : _GEN_7077; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7079 = 6'h27 == _T_820 ? _T_59 : _GEN_7078; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7080 = 6'h28 == _T_820 ? _T_60 : _GEN_7079; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7081 = 6'h29 == _T_820 ? _T_61 : _GEN_7080; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7082 = 6'h2a == _T_820 ? _T_62 : _GEN_7081; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7083 = 6'h2b == _T_820 ? _T_63 : _GEN_7082; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7084 = 6'h2c == _T_820 ? _T_64 : _GEN_7083; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7085 = 6'h2d == _T_820 ? _T_65 : _GEN_7084; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7086 = 6'h2e == _T_820 ? _T_66 : _GEN_7085; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7087 = 6'h2f == _T_820 ? _T_67 : _GEN_7086; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7088 = 6'h30 == _T_820 ? _T_68 : _GEN_7087; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7089 = 6'h31 == _T_820 ? _T_69 : _GEN_7088; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7090 = 6'h32 == _T_820 ? _T_70 : _GEN_7089; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7091 = 6'h33 == _T_820 ? _T_71 : _GEN_7090; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7092 = 6'h34 == _T_820 ? _T_72 : _GEN_7091; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7093 = 6'h35 == _T_820 ? _T_73 : _GEN_7092; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7094 = 6'h36 == _T_820 ? _T_74 : _GEN_7093; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7095 = 6'h37 == _T_820 ? _T_75 : _GEN_7094; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7096 = 6'h38 == _T_820 ? _T_76 : _GEN_7095; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7097 = 6'h39 == _T_820 ? _T_77 : _GEN_7096; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7098 = 6'h3a == _T_820 ? _T_78 : _GEN_7097; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7099 = 6'h3b == _T_820 ? _T_79 : _GEN_7098; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7100 = 6'h3c == _T_820 ? _T_80 : _GEN_7099; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7101 = 6'h3d == _T_820 ? _T_81 : _GEN_7100; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7102 = 6'h3e == _T_820 ? _T_82 : _GEN_7101; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7103 = 6'h3f == _T_820 ? _T_83 : _GEN_7102; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7105 = 6'h1 == _T_824 ? _T_21 : _T_20; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7106 = 6'h2 == _T_824 ? _T_22 : _GEN_7105; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7107 = 6'h3 == _T_824 ? _T_23 : _GEN_7106; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7108 = 6'h4 == _T_824 ? _T_24 : _GEN_7107; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7109 = 6'h5 == _T_824 ? _T_25 : _GEN_7108; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7110 = 6'h6 == _T_824 ? _T_26 : _GEN_7109; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7111 = 6'h7 == _T_824 ? _T_27 : _GEN_7110; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7112 = 6'h8 == _T_824 ? _T_28 : _GEN_7111; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7113 = 6'h9 == _T_824 ? _T_29 : _GEN_7112; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7114 = 6'ha == _T_824 ? _T_30 : _GEN_7113; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7115 = 6'hb == _T_824 ? _T_31 : _GEN_7114; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7116 = 6'hc == _T_824 ? _T_32 : _GEN_7115; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7117 = 6'hd == _T_824 ? _T_33 : _GEN_7116; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7118 = 6'he == _T_824 ? _T_34 : _GEN_7117; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7119 = 6'hf == _T_824 ? _T_35 : _GEN_7118; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7120 = 6'h10 == _T_824 ? _T_36 : _GEN_7119; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7121 = 6'h11 == _T_824 ? _T_37 : _GEN_7120; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7122 = 6'h12 == _T_824 ? _T_38 : _GEN_7121; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7123 = 6'h13 == _T_824 ? _T_39 : _GEN_7122; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7124 = 6'h14 == _T_824 ? _T_40 : _GEN_7123; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7125 = 6'h15 == _T_824 ? _T_41 : _GEN_7124; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7126 = 6'h16 == _T_824 ? _T_42 : _GEN_7125; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7127 = 6'h17 == _T_824 ? _T_43 : _GEN_7126; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7128 = 6'h18 == _T_824 ? _T_44 : _GEN_7127; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7129 = 6'h19 == _T_824 ? _T_45 : _GEN_7128; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7130 = 6'h1a == _T_824 ? _T_46 : _GEN_7129; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7131 = 6'h1b == _T_824 ? _T_47 : _GEN_7130; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7132 = 6'h1c == _T_824 ? _T_48 : _GEN_7131; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7133 = 6'h1d == _T_824 ? _T_49 : _GEN_7132; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7134 = 6'h1e == _T_824 ? _T_50 : _GEN_7133; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7135 = 6'h1f == _T_824 ? _T_51 : _GEN_7134; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7136 = 6'h20 == _T_824 ? _T_52 : _GEN_7135; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7137 = 6'h21 == _T_824 ? _T_53 : _GEN_7136; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7138 = 6'h22 == _T_824 ? _T_54 : _GEN_7137; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7139 = 6'h23 == _T_824 ? _T_55 : _GEN_7138; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7140 = 6'h24 == _T_824 ? _T_56 : _GEN_7139; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7141 = 6'h25 == _T_824 ? _T_57 : _GEN_7140; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7142 = 6'h26 == _T_824 ? _T_58 : _GEN_7141; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7143 = 6'h27 == _T_824 ? _T_59 : _GEN_7142; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7144 = 6'h28 == _T_824 ? _T_60 : _GEN_7143; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7145 = 6'h29 == _T_824 ? _T_61 : _GEN_7144; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7146 = 6'h2a == _T_824 ? _T_62 : _GEN_7145; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7147 = 6'h2b == _T_824 ? _T_63 : _GEN_7146; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7148 = 6'h2c == _T_824 ? _T_64 : _GEN_7147; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7149 = 6'h2d == _T_824 ? _T_65 : _GEN_7148; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7150 = 6'h2e == _T_824 ? _T_66 : _GEN_7149; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7151 = 6'h2f == _T_824 ? _T_67 : _GEN_7150; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7152 = 6'h30 == _T_824 ? _T_68 : _GEN_7151; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7153 = 6'h31 == _T_824 ? _T_69 : _GEN_7152; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7154 = 6'h32 == _T_824 ? _T_70 : _GEN_7153; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7155 = 6'h33 == _T_824 ? _T_71 : _GEN_7154; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7156 = 6'h34 == _T_824 ? _T_72 : _GEN_7155; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7157 = 6'h35 == _T_824 ? _T_73 : _GEN_7156; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7158 = 6'h36 == _T_824 ? _T_74 : _GEN_7157; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7159 = 6'h37 == _T_824 ? _T_75 : _GEN_7158; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7160 = 6'h38 == _T_824 ? _T_76 : _GEN_7159; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7161 = 6'h39 == _T_824 ? _T_77 : _GEN_7160; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7162 = 6'h3a == _T_824 ? _T_78 : _GEN_7161; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7163 = 6'h3b == _T_824 ? _T_79 : _GEN_7162; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7164 = 6'h3c == _T_824 ? _T_80 : _GEN_7163; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7165 = 6'h3d == _T_824 ? _T_81 : _GEN_7164; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7166 = 6'h3e == _T_824 ? _T_82 : _GEN_7165; // @[execute.scala 79:10:@2242.4]
  assign _GEN_7167 = 6'h3f == _T_824 ? _T_83 : _GEN_7166; // @[execute.scala 79:10:@2242.4]
  assign _T_826 = _T_816 ? _GEN_7103 : _GEN_7167; // @[execute.scala 79:10:@2242.4]
  assign _T_828 = io_amount < 6'h8; // @[execute.scala 79:15:@2243.4]
  assign _T_830 = io_amount - 6'h8; // @[execute.scala 79:37:@2244.4]
  assign _T_831 = $unsigned(_T_830); // @[execute.scala 79:37:@2245.4]
  assign _T_832 = _T_831[5:0]; // @[execute.scala 79:37:@2246.4]
  assign _T_835 = 6'h38 + io_amount; // @[execute.scala 79:60:@2247.4]
  assign _T_836 = 6'h38 + io_amount; // @[execute.scala 79:60:@2248.4]
  assign _GEN_7169 = 6'h1 == _T_832 ? _T_21 : _T_20; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7170 = 6'h2 == _T_832 ? _T_22 : _GEN_7169; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7171 = 6'h3 == _T_832 ? _T_23 : _GEN_7170; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7172 = 6'h4 == _T_832 ? _T_24 : _GEN_7171; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7173 = 6'h5 == _T_832 ? _T_25 : _GEN_7172; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7174 = 6'h6 == _T_832 ? _T_26 : _GEN_7173; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7175 = 6'h7 == _T_832 ? _T_27 : _GEN_7174; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7176 = 6'h8 == _T_832 ? _T_28 : _GEN_7175; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7177 = 6'h9 == _T_832 ? _T_29 : _GEN_7176; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7178 = 6'ha == _T_832 ? _T_30 : _GEN_7177; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7179 = 6'hb == _T_832 ? _T_31 : _GEN_7178; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7180 = 6'hc == _T_832 ? _T_32 : _GEN_7179; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7181 = 6'hd == _T_832 ? _T_33 : _GEN_7180; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7182 = 6'he == _T_832 ? _T_34 : _GEN_7181; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7183 = 6'hf == _T_832 ? _T_35 : _GEN_7182; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7184 = 6'h10 == _T_832 ? _T_36 : _GEN_7183; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7185 = 6'h11 == _T_832 ? _T_37 : _GEN_7184; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7186 = 6'h12 == _T_832 ? _T_38 : _GEN_7185; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7187 = 6'h13 == _T_832 ? _T_39 : _GEN_7186; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7188 = 6'h14 == _T_832 ? _T_40 : _GEN_7187; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7189 = 6'h15 == _T_832 ? _T_41 : _GEN_7188; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7190 = 6'h16 == _T_832 ? _T_42 : _GEN_7189; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7191 = 6'h17 == _T_832 ? _T_43 : _GEN_7190; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7192 = 6'h18 == _T_832 ? _T_44 : _GEN_7191; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7193 = 6'h19 == _T_832 ? _T_45 : _GEN_7192; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7194 = 6'h1a == _T_832 ? _T_46 : _GEN_7193; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7195 = 6'h1b == _T_832 ? _T_47 : _GEN_7194; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7196 = 6'h1c == _T_832 ? _T_48 : _GEN_7195; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7197 = 6'h1d == _T_832 ? _T_49 : _GEN_7196; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7198 = 6'h1e == _T_832 ? _T_50 : _GEN_7197; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7199 = 6'h1f == _T_832 ? _T_51 : _GEN_7198; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7200 = 6'h20 == _T_832 ? _T_52 : _GEN_7199; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7201 = 6'h21 == _T_832 ? _T_53 : _GEN_7200; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7202 = 6'h22 == _T_832 ? _T_54 : _GEN_7201; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7203 = 6'h23 == _T_832 ? _T_55 : _GEN_7202; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7204 = 6'h24 == _T_832 ? _T_56 : _GEN_7203; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7205 = 6'h25 == _T_832 ? _T_57 : _GEN_7204; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7206 = 6'h26 == _T_832 ? _T_58 : _GEN_7205; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7207 = 6'h27 == _T_832 ? _T_59 : _GEN_7206; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7208 = 6'h28 == _T_832 ? _T_60 : _GEN_7207; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7209 = 6'h29 == _T_832 ? _T_61 : _GEN_7208; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7210 = 6'h2a == _T_832 ? _T_62 : _GEN_7209; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7211 = 6'h2b == _T_832 ? _T_63 : _GEN_7210; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7212 = 6'h2c == _T_832 ? _T_64 : _GEN_7211; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7213 = 6'h2d == _T_832 ? _T_65 : _GEN_7212; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7214 = 6'h2e == _T_832 ? _T_66 : _GEN_7213; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7215 = 6'h2f == _T_832 ? _T_67 : _GEN_7214; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7216 = 6'h30 == _T_832 ? _T_68 : _GEN_7215; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7217 = 6'h31 == _T_832 ? _T_69 : _GEN_7216; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7218 = 6'h32 == _T_832 ? _T_70 : _GEN_7217; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7219 = 6'h33 == _T_832 ? _T_71 : _GEN_7218; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7220 = 6'h34 == _T_832 ? _T_72 : _GEN_7219; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7221 = 6'h35 == _T_832 ? _T_73 : _GEN_7220; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7222 = 6'h36 == _T_832 ? _T_74 : _GEN_7221; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7223 = 6'h37 == _T_832 ? _T_75 : _GEN_7222; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7224 = 6'h38 == _T_832 ? _T_76 : _GEN_7223; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7225 = 6'h39 == _T_832 ? _T_77 : _GEN_7224; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7226 = 6'h3a == _T_832 ? _T_78 : _GEN_7225; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7227 = 6'h3b == _T_832 ? _T_79 : _GEN_7226; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7228 = 6'h3c == _T_832 ? _T_80 : _GEN_7227; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7229 = 6'h3d == _T_832 ? _T_81 : _GEN_7228; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7230 = 6'h3e == _T_832 ? _T_82 : _GEN_7229; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7231 = 6'h3f == _T_832 ? _T_83 : _GEN_7230; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7233 = 6'h1 == _T_836 ? _T_21 : _T_20; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7234 = 6'h2 == _T_836 ? _T_22 : _GEN_7233; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7235 = 6'h3 == _T_836 ? _T_23 : _GEN_7234; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7236 = 6'h4 == _T_836 ? _T_24 : _GEN_7235; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7237 = 6'h5 == _T_836 ? _T_25 : _GEN_7236; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7238 = 6'h6 == _T_836 ? _T_26 : _GEN_7237; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7239 = 6'h7 == _T_836 ? _T_27 : _GEN_7238; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7240 = 6'h8 == _T_836 ? _T_28 : _GEN_7239; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7241 = 6'h9 == _T_836 ? _T_29 : _GEN_7240; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7242 = 6'ha == _T_836 ? _T_30 : _GEN_7241; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7243 = 6'hb == _T_836 ? _T_31 : _GEN_7242; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7244 = 6'hc == _T_836 ? _T_32 : _GEN_7243; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7245 = 6'hd == _T_836 ? _T_33 : _GEN_7244; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7246 = 6'he == _T_836 ? _T_34 : _GEN_7245; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7247 = 6'hf == _T_836 ? _T_35 : _GEN_7246; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7248 = 6'h10 == _T_836 ? _T_36 : _GEN_7247; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7249 = 6'h11 == _T_836 ? _T_37 : _GEN_7248; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7250 = 6'h12 == _T_836 ? _T_38 : _GEN_7249; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7251 = 6'h13 == _T_836 ? _T_39 : _GEN_7250; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7252 = 6'h14 == _T_836 ? _T_40 : _GEN_7251; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7253 = 6'h15 == _T_836 ? _T_41 : _GEN_7252; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7254 = 6'h16 == _T_836 ? _T_42 : _GEN_7253; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7255 = 6'h17 == _T_836 ? _T_43 : _GEN_7254; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7256 = 6'h18 == _T_836 ? _T_44 : _GEN_7255; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7257 = 6'h19 == _T_836 ? _T_45 : _GEN_7256; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7258 = 6'h1a == _T_836 ? _T_46 : _GEN_7257; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7259 = 6'h1b == _T_836 ? _T_47 : _GEN_7258; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7260 = 6'h1c == _T_836 ? _T_48 : _GEN_7259; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7261 = 6'h1d == _T_836 ? _T_49 : _GEN_7260; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7262 = 6'h1e == _T_836 ? _T_50 : _GEN_7261; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7263 = 6'h1f == _T_836 ? _T_51 : _GEN_7262; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7264 = 6'h20 == _T_836 ? _T_52 : _GEN_7263; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7265 = 6'h21 == _T_836 ? _T_53 : _GEN_7264; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7266 = 6'h22 == _T_836 ? _T_54 : _GEN_7265; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7267 = 6'h23 == _T_836 ? _T_55 : _GEN_7266; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7268 = 6'h24 == _T_836 ? _T_56 : _GEN_7267; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7269 = 6'h25 == _T_836 ? _T_57 : _GEN_7268; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7270 = 6'h26 == _T_836 ? _T_58 : _GEN_7269; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7271 = 6'h27 == _T_836 ? _T_59 : _GEN_7270; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7272 = 6'h28 == _T_836 ? _T_60 : _GEN_7271; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7273 = 6'h29 == _T_836 ? _T_61 : _GEN_7272; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7274 = 6'h2a == _T_836 ? _T_62 : _GEN_7273; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7275 = 6'h2b == _T_836 ? _T_63 : _GEN_7274; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7276 = 6'h2c == _T_836 ? _T_64 : _GEN_7275; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7277 = 6'h2d == _T_836 ? _T_65 : _GEN_7276; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7278 = 6'h2e == _T_836 ? _T_66 : _GEN_7277; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7279 = 6'h2f == _T_836 ? _T_67 : _GEN_7278; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7280 = 6'h30 == _T_836 ? _T_68 : _GEN_7279; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7281 = 6'h31 == _T_836 ? _T_69 : _GEN_7280; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7282 = 6'h32 == _T_836 ? _T_70 : _GEN_7281; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7283 = 6'h33 == _T_836 ? _T_71 : _GEN_7282; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7284 = 6'h34 == _T_836 ? _T_72 : _GEN_7283; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7285 = 6'h35 == _T_836 ? _T_73 : _GEN_7284; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7286 = 6'h36 == _T_836 ? _T_74 : _GEN_7285; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7287 = 6'h37 == _T_836 ? _T_75 : _GEN_7286; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7288 = 6'h38 == _T_836 ? _T_76 : _GEN_7287; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7289 = 6'h39 == _T_836 ? _T_77 : _GEN_7288; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7290 = 6'h3a == _T_836 ? _T_78 : _GEN_7289; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7291 = 6'h3b == _T_836 ? _T_79 : _GEN_7290; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7292 = 6'h3c == _T_836 ? _T_80 : _GEN_7291; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7293 = 6'h3d == _T_836 ? _T_81 : _GEN_7292; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7294 = 6'h3e == _T_836 ? _T_82 : _GEN_7293; // @[execute.scala 79:10:@2249.4]
  assign _GEN_7295 = 6'h3f == _T_836 ? _T_83 : _GEN_7294; // @[execute.scala 79:10:@2249.4]
  assign _T_838 = _T_828 ? _GEN_7231 : _GEN_7295; // @[execute.scala 79:10:@2249.4]
  assign _T_840 = io_amount < 6'h7; // @[execute.scala 79:15:@2250.4]
  assign _T_842 = io_amount - 6'h7; // @[execute.scala 79:37:@2251.4]
  assign _T_843 = $unsigned(_T_842); // @[execute.scala 79:37:@2252.4]
  assign _T_844 = _T_843[5:0]; // @[execute.scala 79:37:@2253.4]
  assign _T_847 = 6'h39 + io_amount; // @[execute.scala 79:60:@2254.4]
  assign _T_848 = 6'h39 + io_amount; // @[execute.scala 79:60:@2255.4]
  assign _GEN_7297 = 6'h1 == _T_844 ? _T_21 : _T_20; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7298 = 6'h2 == _T_844 ? _T_22 : _GEN_7297; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7299 = 6'h3 == _T_844 ? _T_23 : _GEN_7298; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7300 = 6'h4 == _T_844 ? _T_24 : _GEN_7299; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7301 = 6'h5 == _T_844 ? _T_25 : _GEN_7300; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7302 = 6'h6 == _T_844 ? _T_26 : _GEN_7301; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7303 = 6'h7 == _T_844 ? _T_27 : _GEN_7302; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7304 = 6'h8 == _T_844 ? _T_28 : _GEN_7303; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7305 = 6'h9 == _T_844 ? _T_29 : _GEN_7304; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7306 = 6'ha == _T_844 ? _T_30 : _GEN_7305; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7307 = 6'hb == _T_844 ? _T_31 : _GEN_7306; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7308 = 6'hc == _T_844 ? _T_32 : _GEN_7307; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7309 = 6'hd == _T_844 ? _T_33 : _GEN_7308; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7310 = 6'he == _T_844 ? _T_34 : _GEN_7309; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7311 = 6'hf == _T_844 ? _T_35 : _GEN_7310; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7312 = 6'h10 == _T_844 ? _T_36 : _GEN_7311; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7313 = 6'h11 == _T_844 ? _T_37 : _GEN_7312; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7314 = 6'h12 == _T_844 ? _T_38 : _GEN_7313; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7315 = 6'h13 == _T_844 ? _T_39 : _GEN_7314; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7316 = 6'h14 == _T_844 ? _T_40 : _GEN_7315; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7317 = 6'h15 == _T_844 ? _T_41 : _GEN_7316; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7318 = 6'h16 == _T_844 ? _T_42 : _GEN_7317; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7319 = 6'h17 == _T_844 ? _T_43 : _GEN_7318; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7320 = 6'h18 == _T_844 ? _T_44 : _GEN_7319; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7321 = 6'h19 == _T_844 ? _T_45 : _GEN_7320; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7322 = 6'h1a == _T_844 ? _T_46 : _GEN_7321; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7323 = 6'h1b == _T_844 ? _T_47 : _GEN_7322; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7324 = 6'h1c == _T_844 ? _T_48 : _GEN_7323; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7325 = 6'h1d == _T_844 ? _T_49 : _GEN_7324; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7326 = 6'h1e == _T_844 ? _T_50 : _GEN_7325; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7327 = 6'h1f == _T_844 ? _T_51 : _GEN_7326; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7328 = 6'h20 == _T_844 ? _T_52 : _GEN_7327; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7329 = 6'h21 == _T_844 ? _T_53 : _GEN_7328; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7330 = 6'h22 == _T_844 ? _T_54 : _GEN_7329; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7331 = 6'h23 == _T_844 ? _T_55 : _GEN_7330; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7332 = 6'h24 == _T_844 ? _T_56 : _GEN_7331; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7333 = 6'h25 == _T_844 ? _T_57 : _GEN_7332; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7334 = 6'h26 == _T_844 ? _T_58 : _GEN_7333; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7335 = 6'h27 == _T_844 ? _T_59 : _GEN_7334; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7336 = 6'h28 == _T_844 ? _T_60 : _GEN_7335; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7337 = 6'h29 == _T_844 ? _T_61 : _GEN_7336; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7338 = 6'h2a == _T_844 ? _T_62 : _GEN_7337; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7339 = 6'h2b == _T_844 ? _T_63 : _GEN_7338; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7340 = 6'h2c == _T_844 ? _T_64 : _GEN_7339; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7341 = 6'h2d == _T_844 ? _T_65 : _GEN_7340; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7342 = 6'h2e == _T_844 ? _T_66 : _GEN_7341; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7343 = 6'h2f == _T_844 ? _T_67 : _GEN_7342; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7344 = 6'h30 == _T_844 ? _T_68 : _GEN_7343; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7345 = 6'h31 == _T_844 ? _T_69 : _GEN_7344; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7346 = 6'h32 == _T_844 ? _T_70 : _GEN_7345; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7347 = 6'h33 == _T_844 ? _T_71 : _GEN_7346; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7348 = 6'h34 == _T_844 ? _T_72 : _GEN_7347; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7349 = 6'h35 == _T_844 ? _T_73 : _GEN_7348; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7350 = 6'h36 == _T_844 ? _T_74 : _GEN_7349; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7351 = 6'h37 == _T_844 ? _T_75 : _GEN_7350; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7352 = 6'h38 == _T_844 ? _T_76 : _GEN_7351; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7353 = 6'h39 == _T_844 ? _T_77 : _GEN_7352; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7354 = 6'h3a == _T_844 ? _T_78 : _GEN_7353; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7355 = 6'h3b == _T_844 ? _T_79 : _GEN_7354; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7356 = 6'h3c == _T_844 ? _T_80 : _GEN_7355; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7357 = 6'h3d == _T_844 ? _T_81 : _GEN_7356; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7358 = 6'h3e == _T_844 ? _T_82 : _GEN_7357; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7359 = 6'h3f == _T_844 ? _T_83 : _GEN_7358; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7361 = 6'h1 == _T_848 ? _T_21 : _T_20; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7362 = 6'h2 == _T_848 ? _T_22 : _GEN_7361; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7363 = 6'h3 == _T_848 ? _T_23 : _GEN_7362; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7364 = 6'h4 == _T_848 ? _T_24 : _GEN_7363; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7365 = 6'h5 == _T_848 ? _T_25 : _GEN_7364; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7366 = 6'h6 == _T_848 ? _T_26 : _GEN_7365; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7367 = 6'h7 == _T_848 ? _T_27 : _GEN_7366; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7368 = 6'h8 == _T_848 ? _T_28 : _GEN_7367; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7369 = 6'h9 == _T_848 ? _T_29 : _GEN_7368; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7370 = 6'ha == _T_848 ? _T_30 : _GEN_7369; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7371 = 6'hb == _T_848 ? _T_31 : _GEN_7370; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7372 = 6'hc == _T_848 ? _T_32 : _GEN_7371; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7373 = 6'hd == _T_848 ? _T_33 : _GEN_7372; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7374 = 6'he == _T_848 ? _T_34 : _GEN_7373; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7375 = 6'hf == _T_848 ? _T_35 : _GEN_7374; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7376 = 6'h10 == _T_848 ? _T_36 : _GEN_7375; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7377 = 6'h11 == _T_848 ? _T_37 : _GEN_7376; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7378 = 6'h12 == _T_848 ? _T_38 : _GEN_7377; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7379 = 6'h13 == _T_848 ? _T_39 : _GEN_7378; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7380 = 6'h14 == _T_848 ? _T_40 : _GEN_7379; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7381 = 6'h15 == _T_848 ? _T_41 : _GEN_7380; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7382 = 6'h16 == _T_848 ? _T_42 : _GEN_7381; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7383 = 6'h17 == _T_848 ? _T_43 : _GEN_7382; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7384 = 6'h18 == _T_848 ? _T_44 : _GEN_7383; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7385 = 6'h19 == _T_848 ? _T_45 : _GEN_7384; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7386 = 6'h1a == _T_848 ? _T_46 : _GEN_7385; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7387 = 6'h1b == _T_848 ? _T_47 : _GEN_7386; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7388 = 6'h1c == _T_848 ? _T_48 : _GEN_7387; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7389 = 6'h1d == _T_848 ? _T_49 : _GEN_7388; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7390 = 6'h1e == _T_848 ? _T_50 : _GEN_7389; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7391 = 6'h1f == _T_848 ? _T_51 : _GEN_7390; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7392 = 6'h20 == _T_848 ? _T_52 : _GEN_7391; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7393 = 6'h21 == _T_848 ? _T_53 : _GEN_7392; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7394 = 6'h22 == _T_848 ? _T_54 : _GEN_7393; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7395 = 6'h23 == _T_848 ? _T_55 : _GEN_7394; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7396 = 6'h24 == _T_848 ? _T_56 : _GEN_7395; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7397 = 6'h25 == _T_848 ? _T_57 : _GEN_7396; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7398 = 6'h26 == _T_848 ? _T_58 : _GEN_7397; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7399 = 6'h27 == _T_848 ? _T_59 : _GEN_7398; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7400 = 6'h28 == _T_848 ? _T_60 : _GEN_7399; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7401 = 6'h29 == _T_848 ? _T_61 : _GEN_7400; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7402 = 6'h2a == _T_848 ? _T_62 : _GEN_7401; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7403 = 6'h2b == _T_848 ? _T_63 : _GEN_7402; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7404 = 6'h2c == _T_848 ? _T_64 : _GEN_7403; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7405 = 6'h2d == _T_848 ? _T_65 : _GEN_7404; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7406 = 6'h2e == _T_848 ? _T_66 : _GEN_7405; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7407 = 6'h2f == _T_848 ? _T_67 : _GEN_7406; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7408 = 6'h30 == _T_848 ? _T_68 : _GEN_7407; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7409 = 6'h31 == _T_848 ? _T_69 : _GEN_7408; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7410 = 6'h32 == _T_848 ? _T_70 : _GEN_7409; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7411 = 6'h33 == _T_848 ? _T_71 : _GEN_7410; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7412 = 6'h34 == _T_848 ? _T_72 : _GEN_7411; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7413 = 6'h35 == _T_848 ? _T_73 : _GEN_7412; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7414 = 6'h36 == _T_848 ? _T_74 : _GEN_7413; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7415 = 6'h37 == _T_848 ? _T_75 : _GEN_7414; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7416 = 6'h38 == _T_848 ? _T_76 : _GEN_7415; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7417 = 6'h39 == _T_848 ? _T_77 : _GEN_7416; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7418 = 6'h3a == _T_848 ? _T_78 : _GEN_7417; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7419 = 6'h3b == _T_848 ? _T_79 : _GEN_7418; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7420 = 6'h3c == _T_848 ? _T_80 : _GEN_7419; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7421 = 6'h3d == _T_848 ? _T_81 : _GEN_7420; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7422 = 6'h3e == _T_848 ? _T_82 : _GEN_7421; // @[execute.scala 79:10:@2256.4]
  assign _GEN_7423 = 6'h3f == _T_848 ? _T_83 : _GEN_7422; // @[execute.scala 79:10:@2256.4]
  assign _T_850 = _T_840 ? _GEN_7359 : _GEN_7423; // @[execute.scala 79:10:@2256.4]
  assign _T_852 = io_amount < 6'h6; // @[execute.scala 79:15:@2257.4]
  assign _T_854 = io_amount - 6'h6; // @[execute.scala 79:37:@2258.4]
  assign _T_855 = $unsigned(_T_854); // @[execute.scala 79:37:@2259.4]
  assign _T_856 = _T_855[5:0]; // @[execute.scala 79:37:@2260.4]
  assign _T_859 = 6'h3a + io_amount; // @[execute.scala 79:60:@2261.4]
  assign _T_860 = 6'h3a + io_amount; // @[execute.scala 79:60:@2262.4]
  assign _GEN_7425 = 6'h1 == _T_856 ? _T_21 : _T_20; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7426 = 6'h2 == _T_856 ? _T_22 : _GEN_7425; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7427 = 6'h3 == _T_856 ? _T_23 : _GEN_7426; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7428 = 6'h4 == _T_856 ? _T_24 : _GEN_7427; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7429 = 6'h5 == _T_856 ? _T_25 : _GEN_7428; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7430 = 6'h6 == _T_856 ? _T_26 : _GEN_7429; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7431 = 6'h7 == _T_856 ? _T_27 : _GEN_7430; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7432 = 6'h8 == _T_856 ? _T_28 : _GEN_7431; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7433 = 6'h9 == _T_856 ? _T_29 : _GEN_7432; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7434 = 6'ha == _T_856 ? _T_30 : _GEN_7433; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7435 = 6'hb == _T_856 ? _T_31 : _GEN_7434; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7436 = 6'hc == _T_856 ? _T_32 : _GEN_7435; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7437 = 6'hd == _T_856 ? _T_33 : _GEN_7436; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7438 = 6'he == _T_856 ? _T_34 : _GEN_7437; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7439 = 6'hf == _T_856 ? _T_35 : _GEN_7438; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7440 = 6'h10 == _T_856 ? _T_36 : _GEN_7439; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7441 = 6'h11 == _T_856 ? _T_37 : _GEN_7440; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7442 = 6'h12 == _T_856 ? _T_38 : _GEN_7441; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7443 = 6'h13 == _T_856 ? _T_39 : _GEN_7442; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7444 = 6'h14 == _T_856 ? _T_40 : _GEN_7443; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7445 = 6'h15 == _T_856 ? _T_41 : _GEN_7444; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7446 = 6'h16 == _T_856 ? _T_42 : _GEN_7445; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7447 = 6'h17 == _T_856 ? _T_43 : _GEN_7446; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7448 = 6'h18 == _T_856 ? _T_44 : _GEN_7447; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7449 = 6'h19 == _T_856 ? _T_45 : _GEN_7448; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7450 = 6'h1a == _T_856 ? _T_46 : _GEN_7449; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7451 = 6'h1b == _T_856 ? _T_47 : _GEN_7450; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7452 = 6'h1c == _T_856 ? _T_48 : _GEN_7451; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7453 = 6'h1d == _T_856 ? _T_49 : _GEN_7452; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7454 = 6'h1e == _T_856 ? _T_50 : _GEN_7453; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7455 = 6'h1f == _T_856 ? _T_51 : _GEN_7454; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7456 = 6'h20 == _T_856 ? _T_52 : _GEN_7455; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7457 = 6'h21 == _T_856 ? _T_53 : _GEN_7456; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7458 = 6'h22 == _T_856 ? _T_54 : _GEN_7457; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7459 = 6'h23 == _T_856 ? _T_55 : _GEN_7458; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7460 = 6'h24 == _T_856 ? _T_56 : _GEN_7459; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7461 = 6'h25 == _T_856 ? _T_57 : _GEN_7460; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7462 = 6'h26 == _T_856 ? _T_58 : _GEN_7461; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7463 = 6'h27 == _T_856 ? _T_59 : _GEN_7462; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7464 = 6'h28 == _T_856 ? _T_60 : _GEN_7463; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7465 = 6'h29 == _T_856 ? _T_61 : _GEN_7464; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7466 = 6'h2a == _T_856 ? _T_62 : _GEN_7465; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7467 = 6'h2b == _T_856 ? _T_63 : _GEN_7466; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7468 = 6'h2c == _T_856 ? _T_64 : _GEN_7467; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7469 = 6'h2d == _T_856 ? _T_65 : _GEN_7468; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7470 = 6'h2e == _T_856 ? _T_66 : _GEN_7469; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7471 = 6'h2f == _T_856 ? _T_67 : _GEN_7470; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7472 = 6'h30 == _T_856 ? _T_68 : _GEN_7471; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7473 = 6'h31 == _T_856 ? _T_69 : _GEN_7472; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7474 = 6'h32 == _T_856 ? _T_70 : _GEN_7473; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7475 = 6'h33 == _T_856 ? _T_71 : _GEN_7474; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7476 = 6'h34 == _T_856 ? _T_72 : _GEN_7475; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7477 = 6'h35 == _T_856 ? _T_73 : _GEN_7476; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7478 = 6'h36 == _T_856 ? _T_74 : _GEN_7477; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7479 = 6'h37 == _T_856 ? _T_75 : _GEN_7478; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7480 = 6'h38 == _T_856 ? _T_76 : _GEN_7479; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7481 = 6'h39 == _T_856 ? _T_77 : _GEN_7480; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7482 = 6'h3a == _T_856 ? _T_78 : _GEN_7481; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7483 = 6'h3b == _T_856 ? _T_79 : _GEN_7482; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7484 = 6'h3c == _T_856 ? _T_80 : _GEN_7483; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7485 = 6'h3d == _T_856 ? _T_81 : _GEN_7484; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7486 = 6'h3e == _T_856 ? _T_82 : _GEN_7485; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7487 = 6'h3f == _T_856 ? _T_83 : _GEN_7486; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7489 = 6'h1 == _T_860 ? _T_21 : _T_20; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7490 = 6'h2 == _T_860 ? _T_22 : _GEN_7489; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7491 = 6'h3 == _T_860 ? _T_23 : _GEN_7490; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7492 = 6'h4 == _T_860 ? _T_24 : _GEN_7491; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7493 = 6'h5 == _T_860 ? _T_25 : _GEN_7492; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7494 = 6'h6 == _T_860 ? _T_26 : _GEN_7493; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7495 = 6'h7 == _T_860 ? _T_27 : _GEN_7494; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7496 = 6'h8 == _T_860 ? _T_28 : _GEN_7495; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7497 = 6'h9 == _T_860 ? _T_29 : _GEN_7496; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7498 = 6'ha == _T_860 ? _T_30 : _GEN_7497; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7499 = 6'hb == _T_860 ? _T_31 : _GEN_7498; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7500 = 6'hc == _T_860 ? _T_32 : _GEN_7499; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7501 = 6'hd == _T_860 ? _T_33 : _GEN_7500; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7502 = 6'he == _T_860 ? _T_34 : _GEN_7501; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7503 = 6'hf == _T_860 ? _T_35 : _GEN_7502; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7504 = 6'h10 == _T_860 ? _T_36 : _GEN_7503; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7505 = 6'h11 == _T_860 ? _T_37 : _GEN_7504; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7506 = 6'h12 == _T_860 ? _T_38 : _GEN_7505; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7507 = 6'h13 == _T_860 ? _T_39 : _GEN_7506; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7508 = 6'h14 == _T_860 ? _T_40 : _GEN_7507; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7509 = 6'h15 == _T_860 ? _T_41 : _GEN_7508; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7510 = 6'h16 == _T_860 ? _T_42 : _GEN_7509; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7511 = 6'h17 == _T_860 ? _T_43 : _GEN_7510; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7512 = 6'h18 == _T_860 ? _T_44 : _GEN_7511; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7513 = 6'h19 == _T_860 ? _T_45 : _GEN_7512; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7514 = 6'h1a == _T_860 ? _T_46 : _GEN_7513; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7515 = 6'h1b == _T_860 ? _T_47 : _GEN_7514; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7516 = 6'h1c == _T_860 ? _T_48 : _GEN_7515; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7517 = 6'h1d == _T_860 ? _T_49 : _GEN_7516; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7518 = 6'h1e == _T_860 ? _T_50 : _GEN_7517; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7519 = 6'h1f == _T_860 ? _T_51 : _GEN_7518; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7520 = 6'h20 == _T_860 ? _T_52 : _GEN_7519; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7521 = 6'h21 == _T_860 ? _T_53 : _GEN_7520; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7522 = 6'h22 == _T_860 ? _T_54 : _GEN_7521; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7523 = 6'h23 == _T_860 ? _T_55 : _GEN_7522; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7524 = 6'h24 == _T_860 ? _T_56 : _GEN_7523; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7525 = 6'h25 == _T_860 ? _T_57 : _GEN_7524; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7526 = 6'h26 == _T_860 ? _T_58 : _GEN_7525; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7527 = 6'h27 == _T_860 ? _T_59 : _GEN_7526; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7528 = 6'h28 == _T_860 ? _T_60 : _GEN_7527; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7529 = 6'h29 == _T_860 ? _T_61 : _GEN_7528; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7530 = 6'h2a == _T_860 ? _T_62 : _GEN_7529; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7531 = 6'h2b == _T_860 ? _T_63 : _GEN_7530; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7532 = 6'h2c == _T_860 ? _T_64 : _GEN_7531; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7533 = 6'h2d == _T_860 ? _T_65 : _GEN_7532; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7534 = 6'h2e == _T_860 ? _T_66 : _GEN_7533; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7535 = 6'h2f == _T_860 ? _T_67 : _GEN_7534; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7536 = 6'h30 == _T_860 ? _T_68 : _GEN_7535; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7537 = 6'h31 == _T_860 ? _T_69 : _GEN_7536; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7538 = 6'h32 == _T_860 ? _T_70 : _GEN_7537; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7539 = 6'h33 == _T_860 ? _T_71 : _GEN_7538; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7540 = 6'h34 == _T_860 ? _T_72 : _GEN_7539; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7541 = 6'h35 == _T_860 ? _T_73 : _GEN_7540; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7542 = 6'h36 == _T_860 ? _T_74 : _GEN_7541; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7543 = 6'h37 == _T_860 ? _T_75 : _GEN_7542; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7544 = 6'h38 == _T_860 ? _T_76 : _GEN_7543; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7545 = 6'h39 == _T_860 ? _T_77 : _GEN_7544; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7546 = 6'h3a == _T_860 ? _T_78 : _GEN_7545; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7547 = 6'h3b == _T_860 ? _T_79 : _GEN_7546; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7548 = 6'h3c == _T_860 ? _T_80 : _GEN_7547; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7549 = 6'h3d == _T_860 ? _T_81 : _GEN_7548; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7550 = 6'h3e == _T_860 ? _T_82 : _GEN_7549; // @[execute.scala 79:10:@2263.4]
  assign _GEN_7551 = 6'h3f == _T_860 ? _T_83 : _GEN_7550; // @[execute.scala 79:10:@2263.4]
  assign _T_862 = _T_852 ? _GEN_7487 : _GEN_7551; // @[execute.scala 79:10:@2263.4]
  assign _T_864 = io_amount < 6'h5; // @[execute.scala 79:15:@2264.4]
  assign _T_866 = io_amount - 6'h5; // @[execute.scala 79:37:@2265.4]
  assign _T_867 = $unsigned(_T_866); // @[execute.scala 79:37:@2266.4]
  assign _T_868 = _T_867[5:0]; // @[execute.scala 79:37:@2267.4]
  assign _T_871 = 6'h3b + io_amount; // @[execute.scala 79:60:@2268.4]
  assign _T_872 = 6'h3b + io_amount; // @[execute.scala 79:60:@2269.4]
  assign _GEN_7553 = 6'h1 == _T_868 ? _T_21 : _T_20; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7554 = 6'h2 == _T_868 ? _T_22 : _GEN_7553; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7555 = 6'h3 == _T_868 ? _T_23 : _GEN_7554; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7556 = 6'h4 == _T_868 ? _T_24 : _GEN_7555; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7557 = 6'h5 == _T_868 ? _T_25 : _GEN_7556; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7558 = 6'h6 == _T_868 ? _T_26 : _GEN_7557; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7559 = 6'h7 == _T_868 ? _T_27 : _GEN_7558; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7560 = 6'h8 == _T_868 ? _T_28 : _GEN_7559; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7561 = 6'h9 == _T_868 ? _T_29 : _GEN_7560; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7562 = 6'ha == _T_868 ? _T_30 : _GEN_7561; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7563 = 6'hb == _T_868 ? _T_31 : _GEN_7562; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7564 = 6'hc == _T_868 ? _T_32 : _GEN_7563; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7565 = 6'hd == _T_868 ? _T_33 : _GEN_7564; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7566 = 6'he == _T_868 ? _T_34 : _GEN_7565; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7567 = 6'hf == _T_868 ? _T_35 : _GEN_7566; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7568 = 6'h10 == _T_868 ? _T_36 : _GEN_7567; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7569 = 6'h11 == _T_868 ? _T_37 : _GEN_7568; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7570 = 6'h12 == _T_868 ? _T_38 : _GEN_7569; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7571 = 6'h13 == _T_868 ? _T_39 : _GEN_7570; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7572 = 6'h14 == _T_868 ? _T_40 : _GEN_7571; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7573 = 6'h15 == _T_868 ? _T_41 : _GEN_7572; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7574 = 6'h16 == _T_868 ? _T_42 : _GEN_7573; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7575 = 6'h17 == _T_868 ? _T_43 : _GEN_7574; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7576 = 6'h18 == _T_868 ? _T_44 : _GEN_7575; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7577 = 6'h19 == _T_868 ? _T_45 : _GEN_7576; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7578 = 6'h1a == _T_868 ? _T_46 : _GEN_7577; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7579 = 6'h1b == _T_868 ? _T_47 : _GEN_7578; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7580 = 6'h1c == _T_868 ? _T_48 : _GEN_7579; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7581 = 6'h1d == _T_868 ? _T_49 : _GEN_7580; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7582 = 6'h1e == _T_868 ? _T_50 : _GEN_7581; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7583 = 6'h1f == _T_868 ? _T_51 : _GEN_7582; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7584 = 6'h20 == _T_868 ? _T_52 : _GEN_7583; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7585 = 6'h21 == _T_868 ? _T_53 : _GEN_7584; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7586 = 6'h22 == _T_868 ? _T_54 : _GEN_7585; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7587 = 6'h23 == _T_868 ? _T_55 : _GEN_7586; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7588 = 6'h24 == _T_868 ? _T_56 : _GEN_7587; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7589 = 6'h25 == _T_868 ? _T_57 : _GEN_7588; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7590 = 6'h26 == _T_868 ? _T_58 : _GEN_7589; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7591 = 6'h27 == _T_868 ? _T_59 : _GEN_7590; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7592 = 6'h28 == _T_868 ? _T_60 : _GEN_7591; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7593 = 6'h29 == _T_868 ? _T_61 : _GEN_7592; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7594 = 6'h2a == _T_868 ? _T_62 : _GEN_7593; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7595 = 6'h2b == _T_868 ? _T_63 : _GEN_7594; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7596 = 6'h2c == _T_868 ? _T_64 : _GEN_7595; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7597 = 6'h2d == _T_868 ? _T_65 : _GEN_7596; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7598 = 6'h2e == _T_868 ? _T_66 : _GEN_7597; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7599 = 6'h2f == _T_868 ? _T_67 : _GEN_7598; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7600 = 6'h30 == _T_868 ? _T_68 : _GEN_7599; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7601 = 6'h31 == _T_868 ? _T_69 : _GEN_7600; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7602 = 6'h32 == _T_868 ? _T_70 : _GEN_7601; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7603 = 6'h33 == _T_868 ? _T_71 : _GEN_7602; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7604 = 6'h34 == _T_868 ? _T_72 : _GEN_7603; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7605 = 6'h35 == _T_868 ? _T_73 : _GEN_7604; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7606 = 6'h36 == _T_868 ? _T_74 : _GEN_7605; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7607 = 6'h37 == _T_868 ? _T_75 : _GEN_7606; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7608 = 6'h38 == _T_868 ? _T_76 : _GEN_7607; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7609 = 6'h39 == _T_868 ? _T_77 : _GEN_7608; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7610 = 6'h3a == _T_868 ? _T_78 : _GEN_7609; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7611 = 6'h3b == _T_868 ? _T_79 : _GEN_7610; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7612 = 6'h3c == _T_868 ? _T_80 : _GEN_7611; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7613 = 6'h3d == _T_868 ? _T_81 : _GEN_7612; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7614 = 6'h3e == _T_868 ? _T_82 : _GEN_7613; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7615 = 6'h3f == _T_868 ? _T_83 : _GEN_7614; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7617 = 6'h1 == _T_872 ? _T_21 : _T_20; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7618 = 6'h2 == _T_872 ? _T_22 : _GEN_7617; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7619 = 6'h3 == _T_872 ? _T_23 : _GEN_7618; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7620 = 6'h4 == _T_872 ? _T_24 : _GEN_7619; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7621 = 6'h5 == _T_872 ? _T_25 : _GEN_7620; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7622 = 6'h6 == _T_872 ? _T_26 : _GEN_7621; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7623 = 6'h7 == _T_872 ? _T_27 : _GEN_7622; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7624 = 6'h8 == _T_872 ? _T_28 : _GEN_7623; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7625 = 6'h9 == _T_872 ? _T_29 : _GEN_7624; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7626 = 6'ha == _T_872 ? _T_30 : _GEN_7625; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7627 = 6'hb == _T_872 ? _T_31 : _GEN_7626; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7628 = 6'hc == _T_872 ? _T_32 : _GEN_7627; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7629 = 6'hd == _T_872 ? _T_33 : _GEN_7628; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7630 = 6'he == _T_872 ? _T_34 : _GEN_7629; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7631 = 6'hf == _T_872 ? _T_35 : _GEN_7630; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7632 = 6'h10 == _T_872 ? _T_36 : _GEN_7631; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7633 = 6'h11 == _T_872 ? _T_37 : _GEN_7632; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7634 = 6'h12 == _T_872 ? _T_38 : _GEN_7633; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7635 = 6'h13 == _T_872 ? _T_39 : _GEN_7634; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7636 = 6'h14 == _T_872 ? _T_40 : _GEN_7635; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7637 = 6'h15 == _T_872 ? _T_41 : _GEN_7636; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7638 = 6'h16 == _T_872 ? _T_42 : _GEN_7637; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7639 = 6'h17 == _T_872 ? _T_43 : _GEN_7638; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7640 = 6'h18 == _T_872 ? _T_44 : _GEN_7639; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7641 = 6'h19 == _T_872 ? _T_45 : _GEN_7640; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7642 = 6'h1a == _T_872 ? _T_46 : _GEN_7641; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7643 = 6'h1b == _T_872 ? _T_47 : _GEN_7642; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7644 = 6'h1c == _T_872 ? _T_48 : _GEN_7643; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7645 = 6'h1d == _T_872 ? _T_49 : _GEN_7644; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7646 = 6'h1e == _T_872 ? _T_50 : _GEN_7645; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7647 = 6'h1f == _T_872 ? _T_51 : _GEN_7646; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7648 = 6'h20 == _T_872 ? _T_52 : _GEN_7647; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7649 = 6'h21 == _T_872 ? _T_53 : _GEN_7648; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7650 = 6'h22 == _T_872 ? _T_54 : _GEN_7649; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7651 = 6'h23 == _T_872 ? _T_55 : _GEN_7650; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7652 = 6'h24 == _T_872 ? _T_56 : _GEN_7651; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7653 = 6'h25 == _T_872 ? _T_57 : _GEN_7652; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7654 = 6'h26 == _T_872 ? _T_58 : _GEN_7653; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7655 = 6'h27 == _T_872 ? _T_59 : _GEN_7654; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7656 = 6'h28 == _T_872 ? _T_60 : _GEN_7655; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7657 = 6'h29 == _T_872 ? _T_61 : _GEN_7656; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7658 = 6'h2a == _T_872 ? _T_62 : _GEN_7657; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7659 = 6'h2b == _T_872 ? _T_63 : _GEN_7658; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7660 = 6'h2c == _T_872 ? _T_64 : _GEN_7659; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7661 = 6'h2d == _T_872 ? _T_65 : _GEN_7660; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7662 = 6'h2e == _T_872 ? _T_66 : _GEN_7661; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7663 = 6'h2f == _T_872 ? _T_67 : _GEN_7662; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7664 = 6'h30 == _T_872 ? _T_68 : _GEN_7663; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7665 = 6'h31 == _T_872 ? _T_69 : _GEN_7664; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7666 = 6'h32 == _T_872 ? _T_70 : _GEN_7665; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7667 = 6'h33 == _T_872 ? _T_71 : _GEN_7666; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7668 = 6'h34 == _T_872 ? _T_72 : _GEN_7667; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7669 = 6'h35 == _T_872 ? _T_73 : _GEN_7668; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7670 = 6'h36 == _T_872 ? _T_74 : _GEN_7669; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7671 = 6'h37 == _T_872 ? _T_75 : _GEN_7670; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7672 = 6'h38 == _T_872 ? _T_76 : _GEN_7671; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7673 = 6'h39 == _T_872 ? _T_77 : _GEN_7672; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7674 = 6'h3a == _T_872 ? _T_78 : _GEN_7673; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7675 = 6'h3b == _T_872 ? _T_79 : _GEN_7674; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7676 = 6'h3c == _T_872 ? _T_80 : _GEN_7675; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7677 = 6'h3d == _T_872 ? _T_81 : _GEN_7676; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7678 = 6'h3e == _T_872 ? _T_82 : _GEN_7677; // @[execute.scala 79:10:@2270.4]
  assign _GEN_7679 = 6'h3f == _T_872 ? _T_83 : _GEN_7678; // @[execute.scala 79:10:@2270.4]
  assign _T_874 = _T_864 ? _GEN_7615 : _GEN_7679; // @[execute.scala 79:10:@2270.4]
  assign _T_876 = io_amount < 6'h4; // @[execute.scala 79:15:@2271.4]
  assign _T_878 = io_amount - 6'h4; // @[execute.scala 79:37:@2272.4]
  assign _T_879 = $unsigned(_T_878); // @[execute.scala 79:37:@2273.4]
  assign _T_880 = _T_879[5:0]; // @[execute.scala 79:37:@2274.4]
  assign _T_883 = 6'h3c + io_amount; // @[execute.scala 79:60:@2275.4]
  assign _T_884 = 6'h3c + io_amount; // @[execute.scala 79:60:@2276.4]
  assign _GEN_7681 = 6'h1 == _T_880 ? _T_21 : _T_20; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7682 = 6'h2 == _T_880 ? _T_22 : _GEN_7681; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7683 = 6'h3 == _T_880 ? _T_23 : _GEN_7682; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7684 = 6'h4 == _T_880 ? _T_24 : _GEN_7683; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7685 = 6'h5 == _T_880 ? _T_25 : _GEN_7684; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7686 = 6'h6 == _T_880 ? _T_26 : _GEN_7685; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7687 = 6'h7 == _T_880 ? _T_27 : _GEN_7686; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7688 = 6'h8 == _T_880 ? _T_28 : _GEN_7687; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7689 = 6'h9 == _T_880 ? _T_29 : _GEN_7688; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7690 = 6'ha == _T_880 ? _T_30 : _GEN_7689; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7691 = 6'hb == _T_880 ? _T_31 : _GEN_7690; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7692 = 6'hc == _T_880 ? _T_32 : _GEN_7691; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7693 = 6'hd == _T_880 ? _T_33 : _GEN_7692; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7694 = 6'he == _T_880 ? _T_34 : _GEN_7693; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7695 = 6'hf == _T_880 ? _T_35 : _GEN_7694; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7696 = 6'h10 == _T_880 ? _T_36 : _GEN_7695; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7697 = 6'h11 == _T_880 ? _T_37 : _GEN_7696; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7698 = 6'h12 == _T_880 ? _T_38 : _GEN_7697; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7699 = 6'h13 == _T_880 ? _T_39 : _GEN_7698; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7700 = 6'h14 == _T_880 ? _T_40 : _GEN_7699; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7701 = 6'h15 == _T_880 ? _T_41 : _GEN_7700; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7702 = 6'h16 == _T_880 ? _T_42 : _GEN_7701; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7703 = 6'h17 == _T_880 ? _T_43 : _GEN_7702; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7704 = 6'h18 == _T_880 ? _T_44 : _GEN_7703; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7705 = 6'h19 == _T_880 ? _T_45 : _GEN_7704; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7706 = 6'h1a == _T_880 ? _T_46 : _GEN_7705; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7707 = 6'h1b == _T_880 ? _T_47 : _GEN_7706; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7708 = 6'h1c == _T_880 ? _T_48 : _GEN_7707; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7709 = 6'h1d == _T_880 ? _T_49 : _GEN_7708; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7710 = 6'h1e == _T_880 ? _T_50 : _GEN_7709; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7711 = 6'h1f == _T_880 ? _T_51 : _GEN_7710; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7712 = 6'h20 == _T_880 ? _T_52 : _GEN_7711; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7713 = 6'h21 == _T_880 ? _T_53 : _GEN_7712; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7714 = 6'h22 == _T_880 ? _T_54 : _GEN_7713; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7715 = 6'h23 == _T_880 ? _T_55 : _GEN_7714; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7716 = 6'h24 == _T_880 ? _T_56 : _GEN_7715; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7717 = 6'h25 == _T_880 ? _T_57 : _GEN_7716; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7718 = 6'h26 == _T_880 ? _T_58 : _GEN_7717; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7719 = 6'h27 == _T_880 ? _T_59 : _GEN_7718; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7720 = 6'h28 == _T_880 ? _T_60 : _GEN_7719; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7721 = 6'h29 == _T_880 ? _T_61 : _GEN_7720; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7722 = 6'h2a == _T_880 ? _T_62 : _GEN_7721; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7723 = 6'h2b == _T_880 ? _T_63 : _GEN_7722; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7724 = 6'h2c == _T_880 ? _T_64 : _GEN_7723; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7725 = 6'h2d == _T_880 ? _T_65 : _GEN_7724; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7726 = 6'h2e == _T_880 ? _T_66 : _GEN_7725; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7727 = 6'h2f == _T_880 ? _T_67 : _GEN_7726; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7728 = 6'h30 == _T_880 ? _T_68 : _GEN_7727; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7729 = 6'h31 == _T_880 ? _T_69 : _GEN_7728; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7730 = 6'h32 == _T_880 ? _T_70 : _GEN_7729; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7731 = 6'h33 == _T_880 ? _T_71 : _GEN_7730; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7732 = 6'h34 == _T_880 ? _T_72 : _GEN_7731; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7733 = 6'h35 == _T_880 ? _T_73 : _GEN_7732; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7734 = 6'h36 == _T_880 ? _T_74 : _GEN_7733; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7735 = 6'h37 == _T_880 ? _T_75 : _GEN_7734; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7736 = 6'h38 == _T_880 ? _T_76 : _GEN_7735; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7737 = 6'h39 == _T_880 ? _T_77 : _GEN_7736; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7738 = 6'h3a == _T_880 ? _T_78 : _GEN_7737; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7739 = 6'h3b == _T_880 ? _T_79 : _GEN_7738; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7740 = 6'h3c == _T_880 ? _T_80 : _GEN_7739; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7741 = 6'h3d == _T_880 ? _T_81 : _GEN_7740; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7742 = 6'h3e == _T_880 ? _T_82 : _GEN_7741; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7743 = 6'h3f == _T_880 ? _T_83 : _GEN_7742; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7745 = 6'h1 == _T_884 ? _T_21 : _T_20; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7746 = 6'h2 == _T_884 ? _T_22 : _GEN_7745; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7747 = 6'h3 == _T_884 ? _T_23 : _GEN_7746; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7748 = 6'h4 == _T_884 ? _T_24 : _GEN_7747; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7749 = 6'h5 == _T_884 ? _T_25 : _GEN_7748; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7750 = 6'h6 == _T_884 ? _T_26 : _GEN_7749; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7751 = 6'h7 == _T_884 ? _T_27 : _GEN_7750; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7752 = 6'h8 == _T_884 ? _T_28 : _GEN_7751; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7753 = 6'h9 == _T_884 ? _T_29 : _GEN_7752; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7754 = 6'ha == _T_884 ? _T_30 : _GEN_7753; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7755 = 6'hb == _T_884 ? _T_31 : _GEN_7754; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7756 = 6'hc == _T_884 ? _T_32 : _GEN_7755; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7757 = 6'hd == _T_884 ? _T_33 : _GEN_7756; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7758 = 6'he == _T_884 ? _T_34 : _GEN_7757; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7759 = 6'hf == _T_884 ? _T_35 : _GEN_7758; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7760 = 6'h10 == _T_884 ? _T_36 : _GEN_7759; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7761 = 6'h11 == _T_884 ? _T_37 : _GEN_7760; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7762 = 6'h12 == _T_884 ? _T_38 : _GEN_7761; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7763 = 6'h13 == _T_884 ? _T_39 : _GEN_7762; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7764 = 6'h14 == _T_884 ? _T_40 : _GEN_7763; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7765 = 6'h15 == _T_884 ? _T_41 : _GEN_7764; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7766 = 6'h16 == _T_884 ? _T_42 : _GEN_7765; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7767 = 6'h17 == _T_884 ? _T_43 : _GEN_7766; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7768 = 6'h18 == _T_884 ? _T_44 : _GEN_7767; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7769 = 6'h19 == _T_884 ? _T_45 : _GEN_7768; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7770 = 6'h1a == _T_884 ? _T_46 : _GEN_7769; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7771 = 6'h1b == _T_884 ? _T_47 : _GEN_7770; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7772 = 6'h1c == _T_884 ? _T_48 : _GEN_7771; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7773 = 6'h1d == _T_884 ? _T_49 : _GEN_7772; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7774 = 6'h1e == _T_884 ? _T_50 : _GEN_7773; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7775 = 6'h1f == _T_884 ? _T_51 : _GEN_7774; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7776 = 6'h20 == _T_884 ? _T_52 : _GEN_7775; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7777 = 6'h21 == _T_884 ? _T_53 : _GEN_7776; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7778 = 6'h22 == _T_884 ? _T_54 : _GEN_7777; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7779 = 6'h23 == _T_884 ? _T_55 : _GEN_7778; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7780 = 6'h24 == _T_884 ? _T_56 : _GEN_7779; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7781 = 6'h25 == _T_884 ? _T_57 : _GEN_7780; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7782 = 6'h26 == _T_884 ? _T_58 : _GEN_7781; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7783 = 6'h27 == _T_884 ? _T_59 : _GEN_7782; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7784 = 6'h28 == _T_884 ? _T_60 : _GEN_7783; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7785 = 6'h29 == _T_884 ? _T_61 : _GEN_7784; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7786 = 6'h2a == _T_884 ? _T_62 : _GEN_7785; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7787 = 6'h2b == _T_884 ? _T_63 : _GEN_7786; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7788 = 6'h2c == _T_884 ? _T_64 : _GEN_7787; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7789 = 6'h2d == _T_884 ? _T_65 : _GEN_7788; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7790 = 6'h2e == _T_884 ? _T_66 : _GEN_7789; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7791 = 6'h2f == _T_884 ? _T_67 : _GEN_7790; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7792 = 6'h30 == _T_884 ? _T_68 : _GEN_7791; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7793 = 6'h31 == _T_884 ? _T_69 : _GEN_7792; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7794 = 6'h32 == _T_884 ? _T_70 : _GEN_7793; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7795 = 6'h33 == _T_884 ? _T_71 : _GEN_7794; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7796 = 6'h34 == _T_884 ? _T_72 : _GEN_7795; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7797 = 6'h35 == _T_884 ? _T_73 : _GEN_7796; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7798 = 6'h36 == _T_884 ? _T_74 : _GEN_7797; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7799 = 6'h37 == _T_884 ? _T_75 : _GEN_7798; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7800 = 6'h38 == _T_884 ? _T_76 : _GEN_7799; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7801 = 6'h39 == _T_884 ? _T_77 : _GEN_7800; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7802 = 6'h3a == _T_884 ? _T_78 : _GEN_7801; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7803 = 6'h3b == _T_884 ? _T_79 : _GEN_7802; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7804 = 6'h3c == _T_884 ? _T_80 : _GEN_7803; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7805 = 6'h3d == _T_884 ? _T_81 : _GEN_7804; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7806 = 6'h3e == _T_884 ? _T_82 : _GEN_7805; // @[execute.scala 79:10:@2277.4]
  assign _GEN_7807 = 6'h3f == _T_884 ? _T_83 : _GEN_7806; // @[execute.scala 79:10:@2277.4]
  assign _T_886 = _T_876 ? _GEN_7743 : _GEN_7807; // @[execute.scala 79:10:@2277.4]
  assign _T_888 = io_amount < 6'h3; // @[execute.scala 79:15:@2278.4]
  assign _T_890 = io_amount - 6'h3; // @[execute.scala 79:37:@2279.4]
  assign _T_891 = $unsigned(_T_890); // @[execute.scala 79:37:@2280.4]
  assign _T_892 = _T_891[5:0]; // @[execute.scala 79:37:@2281.4]
  assign _T_895 = 6'h3d + io_amount; // @[execute.scala 79:60:@2282.4]
  assign _T_896 = 6'h3d + io_amount; // @[execute.scala 79:60:@2283.4]
  assign _GEN_7809 = 6'h1 == _T_892 ? _T_21 : _T_20; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7810 = 6'h2 == _T_892 ? _T_22 : _GEN_7809; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7811 = 6'h3 == _T_892 ? _T_23 : _GEN_7810; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7812 = 6'h4 == _T_892 ? _T_24 : _GEN_7811; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7813 = 6'h5 == _T_892 ? _T_25 : _GEN_7812; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7814 = 6'h6 == _T_892 ? _T_26 : _GEN_7813; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7815 = 6'h7 == _T_892 ? _T_27 : _GEN_7814; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7816 = 6'h8 == _T_892 ? _T_28 : _GEN_7815; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7817 = 6'h9 == _T_892 ? _T_29 : _GEN_7816; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7818 = 6'ha == _T_892 ? _T_30 : _GEN_7817; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7819 = 6'hb == _T_892 ? _T_31 : _GEN_7818; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7820 = 6'hc == _T_892 ? _T_32 : _GEN_7819; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7821 = 6'hd == _T_892 ? _T_33 : _GEN_7820; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7822 = 6'he == _T_892 ? _T_34 : _GEN_7821; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7823 = 6'hf == _T_892 ? _T_35 : _GEN_7822; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7824 = 6'h10 == _T_892 ? _T_36 : _GEN_7823; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7825 = 6'h11 == _T_892 ? _T_37 : _GEN_7824; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7826 = 6'h12 == _T_892 ? _T_38 : _GEN_7825; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7827 = 6'h13 == _T_892 ? _T_39 : _GEN_7826; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7828 = 6'h14 == _T_892 ? _T_40 : _GEN_7827; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7829 = 6'h15 == _T_892 ? _T_41 : _GEN_7828; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7830 = 6'h16 == _T_892 ? _T_42 : _GEN_7829; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7831 = 6'h17 == _T_892 ? _T_43 : _GEN_7830; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7832 = 6'h18 == _T_892 ? _T_44 : _GEN_7831; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7833 = 6'h19 == _T_892 ? _T_45 : _GEN_7832; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7834 = 6'h1a == _T_892 ? _T_46 : _GEN_7833; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7835 = 6'h1b == _T_892 ? _T_47 : _GEN_7834; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7836 = 6'h1c == _T_892 ? _T_48 : _GEN_7835; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7837 = 6'h1d == _T_892 ? _T_49 : _GEN_7836; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7838 = 6'h1e == _T_892 ? _T_50 : _GEN_7837; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7839 = 6'h1f == _T_892 ? _T_51 : _GEN_7838; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7840 = 6'h20 == _T_892 ? _T_52 : _GEN_7839; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7841 = 6'h21 == _T_892 ? _T_53 : _GEN_7840; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7842 = 6'h22 == _T_892 ? _T_54 : _GEN_7841; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7843 = 6'h23 == _T_892 ? _T_55 : _GEN_7842; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7844 = 6'h24 == _T_892 ? _T_56 : _GEN_7843; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7845 = 6'h25 == _T_892 ? _T_57 : _GEN_7844; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7846 = 6'h26 == _T_892 ? _T_58 : _GEN_7845; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7847 = 6'h27 == _T_892 ? _T_59 : _GEN_7846; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7848 = 6'h28 == _T_892 ? _T_60 : _GEN_7847; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7849 = 6'h29 == _T_892 ? _T_61 : _GEN_7848; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7850 = 6'h2a == _T_892 ? _T_62 : _GEN_7849; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7851 = 6'h2b == _T_892 ? _T_63 : _GEN_7850; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7852 = 6'h2c == _T_892 ? _T_64 : _GEN_7851; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7853 = 6'h2d == _T_892 ? _T_65 : _GEN_7852; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7854 = 6'h2e == _T_892 ? _T_66 : _GEN_7853; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7855 = 6'h2f == _T_892 ? _T_67 : _GEN_7854; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7856 = 6'h30 == _T_892 ? _T_68 : _GEN_7855; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7857 = 6'h31 == _T_892 ? _T_69 : _GEN_7856; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7858 = 6'h32 == _T_892 ? _T_70 : _GEN_7857; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7859 = 6'h33 == _T_892 ? _T_71 : _GEN_7858; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7860 = 6'h34 == _T_892 ? _T_72 : _GEN_7859; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7861 = 6'h35 == _T_892 ? _T_73 : _GEN_7860; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7862 = 6'h36 == _T_892 ? _T_74 : _GEN_7861; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7863 = 6'h37 == _T_892 ? _T_75 : _GEN_7862; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7864 = 6'h38 == _T_892 ? _T_76 : _GEN_7863; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7865 = 6'h39 == _T_892 ? _T_77 : _GEN_7864; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7866 = 6'h3a == _T_892 ? _T_78 : _GEN_7865; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7867 = 6'h3b == _T_892 ? _T_79 : _GEN_7866; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7868 = 6'h3c == _T_892 ? _T_80 : _GEN_7867; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7869 = 6'h3d == _T_892 ? _T_81 : _GEN_7868; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7870 = 6'h3e == _T_892 ? _T_82 : _GEN_7869; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7871 = 6'h3f == _T_892 ? _T_83 : _GEN_7870; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7873 = 6'h1 == _T_896 ? _T_21 : _T_20; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7874 = 6'h2 == _T_896 ? _T_22 : _GEN_7873; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7875 = 6'h3 == _T_896 ? _T_23 : _GEN_7874; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7876 = 6'h4 == _T_896 ? _T_24 : _GEN_7875; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7877 = 6'h5 == _T_896 ? _T_25 : _GEN_7876; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7878 = 6'h6 == _T_896 ? _T_26 : _GEN_7877; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7879 = 6'h7 == _T_896 ? _T_27 : _GEN_7878; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7880 = 6'h8 == _T_896 ? _T_28 : _GEN_7879; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7881 = 6'h9 == _T_896 ? _T_29 : _GEN_7880; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7882 = 6'ha == _T_896 ? _T_30 : _GEN_7881; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7883 = 6'hb == _T_896 ? _T_31 : _GEN_7882; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7884 = 6'hc == _T_896 ? _T_32 : _GEN_7883; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7885 = 6'hd == _T_896 ? _T_33 : _GEN_7884; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7886 = 6'he == _T_896 ? _T_34 : _GEN_7885; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7887 = 6'hf == _T_896 ? _T_35 : _GEN_7886; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7888 = 6'h10 == _T_896 ? _T_36 : _GEN_7887; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7889 = 6'h11 == _T_896 ? _T_37 : _GEN_7888; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7890 = 6'h12 == _T_896 ? _T_38 : _GEN_7889; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7891 = 6'h13 == _T_896 ? _T_39 : _GEN_7890; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7892 = 6'h14 == _T_896 ? _T_40 : _GEN_7891; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7893 = 6'h15 == _T_896 ? _T_41 : _GEN_7892; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7894 = 6'h16 == _T_896 ? _T_42 : _GEN_7893; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7895 = 6'h17 == _T_896 ? _T_43 : _GEN_7894; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7896 = 6'h18 == _T_896 ? _T_44 : _GEN_7895; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7897 = 6'h19 == _T_896 ? _T_45 : _GEN_7896; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7898 = 6'h1a == _T_896 ? _T_46 : _GEN_7897; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7899 = 6'h1b == _T_896 ? _T_47 : _GEN_7898; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7900 = 6'h1c == _T_896 ? _T_48 : _GEN_7899; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7901 = 6'h1d == _T_896 ? _T_49 : _GEN_7900; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7902 = 6'h1e == _T_896 ? _T_50 : _GEN_7901; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7903 = 6'h1f == _T_896 ? _T_51 : _GEN_7902; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7904 = 6'h20 == _T_896 ? _T_52 : _GEN_7903; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7905 = 6'h21 == _T_896 ? _T_53 : _GEN_7904; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7906 = 6'h22 == _T_896 ? _T_54 : _GEN_7905; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7907 = 6'h23 == _T_896 ? _T_55 : _GEN_7906; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7908 = 6'h24 == _T_896 ? _T_56 : _GEN_7907; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7909 = 6'h25 == _T_896 ? _T_57 : _GEN_7908; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7910 = 6'h26 == _T_896 ? _T_58 : _GEN_7909; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7911 = 6'h27 == _T_896 ? _T_59 : _GEN_7910; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7912 = 6'h28 == _T_896 ? _T_60 : _GEN_7911; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7913 = 6'h29 == _T_896 ? _T_61 : _GEN_7912; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7914 = 6'h2a == _T_896 ? _T_62 : _GEN_7913; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7915 = 6'h2b == _T_896 ? _T_63 : _GEN_7914; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7916 = 6'h2c == _T_896 ? _T_64 : _GEN_7915; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7917 = 6'h2d == _T_896 ? _T_65 : _GEN_7916; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7918 = 6'h2e == _T_896 ? _T_66 : _GEN_7917; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7919 = 6'h2f == _T_896 ? _T_67 : _GEN_7918; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7920 = 6'h30 == _T_896 ? _T_68 : _GEN_7919; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7921 = 6'h31 == _T_896 ? _T_69 : _GEN_7920; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7922 = 6'h32 == _T_896 ? _T_70 : _GEN_7921; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7923 = 6'h33 == _T_896 ? _T_71 : _GEN_7922; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7924 = 6'h34 == _T_896 ? _T_72 : _GEN_7923; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7925 = 6'h35 == _T_896 ? _T_73 : _GEN_7924; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7926 = 6'h36 == _T_896 ? _T_74 : _GEN_7925; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7927 = 6'h37 == _T_896 ? _T_75 : _GEN_7926; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7928 = 6'h38 == _T_896 ? _T_76 : _GEN_7927; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7929 = 6'h39 == _T_896 ? _T_77 : _GEN_7928; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7930 = 6'h3a == _T_896 ? _T_78 : _GEN_7929; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7931 = 6'h3b == _T_896 ? _T_79 : _GEN_7930; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7932 = 6'h3c == _T_896 ? _T_80 : _GEN_7931; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7933 = 6'h3d == _T_896 ? _T_81 : _GEN_7932; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7934 = 6'h3e == _T_896 ? _T_82 : _GEN_7933; // @[execute.scala 79:10:@2284.4]
  assign _GEN_7935 = 6'h3f == _T_896 ? _T_83 : _GEN_7934; // @[execute.scala 79:10:@2284.4]
  assign _T_898 = _T_888 ? _GEN_7871 : _GEN_7935; // @[execute.scala 79:10:@2284.4]
  assign _T_900 = io_amount < 6'h2; // @[execute.scala 79:15:@2285.4]
  assign _T_902 = io_amount - 6'h2; // @[execute.scala 79:37:@2286.4]
  assign _T_903 = $unsigned(_T_902); // @[execute.scala 79:37:@2287.4]
  assign _T_904 = _T_903[5:0]; // @[execute.scala 79:37:@2288.4]
  assign _T_907 = 6'h3e + io_amount; // @[execute.scala 79:60:@2289.4]
  assign _T_908 = 6'h3e + io_amount; // @[execute.scala 79:60:@2290.4]
  assign _GEN_7937 = 6'h1 == _T_904 ? _T_21 : _T_20; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7938 = 6'h2 == _T_904 ? _T_22 : _GEN_7937; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7939 = 6'h3 == _T_904 ? _T_23 : _GEN_7938; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7940 = 6'h4 == _T_904 ? _T_24 : _GEN_7939; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7941 = 6'h5 == _T_904 ? _T_25 : _GEN_7940; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7942 = 6'h6 == _T_904 ? _T_26 : _GEN_7941; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7943 = 6'h7 == _T_904 ? _T_27 : _GEN_7942; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7944 = 6'h8 == _T_904 ? _T_28 : _GEN_7943; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7945 = 6'h9 == _T_904 ? _T_29 : _GEN_7944; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7946 = 6'ha == _T_904 ? _T_30 : _GEN_7945; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7947 = 6'hb == _T_904 ? _T_31 : _GEN_7946; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7948 = 6'hc == _T_904 ? _T_32 : _GEN_7947; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7949 = 6'hd == _T_904 ? _T_33 : _GEN_7948; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7950 = 6'he == _T_904 ? _T_34 : _GEN_7949; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7951 = 6'hf == _T_904 ? _T_35 : _GEN_7950; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7952 = 6'h10 == _T_904 ? _T_36 : _GEN_7951; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7953 = 6'h11 == _T_904 ? _T_37 : _GEN_7952; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7954 = 6'h12 == _T_904 ? _T_38 : _GEN_7953; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7955 = 6'h13 == _T_904 ? _T_39 : _GEN_7954; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7956 = 6'h14 == _T_904 ? _T_40 : _GEN_7955; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7957 = 6'h15 == _T_904 ? _T_41 : _GEN_7956; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7958 = 6'h16 == _T_904 ? _T_42 : _GEN_7957; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7959 = 6'h17 == _T_904 ? _T_43 : _GEN_7958; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7960 = 6'h18 == _T_904 ? _T_44 : _GEN_7959; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7961 = 6'h19 == _T_904 ? _T_45 : _GEN_7960; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7962 = 6'h1a == _T_904 ? _T_46 : _GEN_7961; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7963 = 6'h1b == _T_904 ? _T_47 : _GEN_7962; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7964 = 6'h1c == _T_904 ? _T_48 : _GEN_7963; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7965 = 6'h1d == _T_904 ? _T_49 : _GEN_7964; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7966 = 6'h1e == _T_904 ? _T_50 : _GEN_7965; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7967 = 6'h1f == _T_904 ? _T_51 : _GEN_7966; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7968 = 6'h20 == _T_904 ? _T_52 : _GEN_7967; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7969 = 6'h21 == _T_904 ? _T_53 : _GEN_7968; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7970 = 6'h22 == _T_904 ? _T_54 : _GEN_7969; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7971 = 6'h23 == _T_904 ? _T_55 : _GEN_7970; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7972 = 6'h24 == _T_904 ? _T_56 : _GEN_7971; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7973 = 6'h25 == _T_904 ? _T_57 : _GEN_7972; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7974 = 6'h26 == _T_904 ? _T_58 : _GEN_7973; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7975 = 6'h27 == _T_904 ? _T_59 : _GEN_7974; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7976 = 6'h28 == _T_904 ? _T_60 : _GEN_7975; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7977 = 6'h29 == _T_904 ? _T_61 : _GEN_7976; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7978 = 6'h2a == _T_904 ? _T_62 : _GEN_7977; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7979 = 6'h2b == _T_904 ? _T_63 : _GEN_7978; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7980 = 6'h2c == _T_904 ? _T_64 : _GEN_7979; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7981 = 6'h2d == _T_904 ? _T_65 : _GEN_7980; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7982 = 6'h2e == _T_904 ? _T_66 : _GEN_7981; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7983 = 6'h2f == _T_904 ? _T_67 : _GEN_7982; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7984 = 6'h30 == _T_904 ? _T_68 : _GEN_7983; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7985 = 6'h31 == _T_904 ? _T_69 : _GEN_7984; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7986 = 6'h32 == _T_904 ? _T_70 : _GEN_7985; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7987 = 6'h33 == _T_904 ? _T_71 : _GEN_7986; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7988 = 6'h34 == _T_904 ? _T_72 : _GEN_7987; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7989 = 6'h35 == _T_904 ? _T_73 : _GEN_7988; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7990 = 6'h36 == _T_904 ? _T_74 : _GEN_7989; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7991 = 6'h37 == _T_904 ? _T_75 : _GEN_7990; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7992 = 6'h38 == _T_904 ? _T_76 : _GEN_7991; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7993 = 6'h39 == _T_904 ? _T_77 : _GEN_7992; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7994 = 6'h3a == _T_904 ? _T_78 : _GEN_7993; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7995 = 6'h3b == _T_904 ? _T_79 : _GEN_7994; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7996 = 6'h3c == _T_904 ? _T_80 : _GEN_7995; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7997 = 6'h3d == _T_904 ? _T_81 : _GEN_7996; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7998 = 6'h3e == _T_904 ? _T_82 : _GEN_7997; // @[execute.scala 79:10:@2291.4]
  assign _GEN_7999 = 6'h3f == _T_904 ? _T_83 : _GEN_7998; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8001 = 6'h1 == _T_908 ? _T_21 : _T_20; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8002 = 6'h2 == _T_908 ? _T_22 : _GEN_8001; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8003 = 6'h3 == _T_908 ? _T_23 : _GEN_8002; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8004 = 6'h4 == _T_908 ? _T_24 : _GEN_8003; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8005 = 6'h5 == _T_908 ? _T_25 : _GEN_8004; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8006 = 6'h6 == _T_908 ? _T_26 : _GEN_8005; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8007 = 6'h7 == _T_908 ? _T_27 : _GEN_8006; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8008 = 6'h8 == _T_908 ? _T_28 : _GEN_8007; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8009 = 6'h9 == _T_908 ? _T_29 : _GEN_8008; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8010 = 6'ha == _T_908 ? _T_30 : _GEN_8009; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8011 = 6'hb == _T_908 ? _T_31 : _GEN_8010; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8012 = 6'hc == _T_908 ? _T_32 : _GEN_8011; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8013 = 6'hd == _T_908 ? _T_33 : _GEN_8012; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8014 = 6'he == _T_908 ? _T_34 : _GEN_8013; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8015 = 6'hf == _T_908 ? _T_35 : _GEN_8014; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8016 = 6'h10 == _T_908 ? _T_36 : _GEN_8015; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8017 = 6'h11 == _T_908 ? _T_37 : _GEN_8016; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8018 = 6'h12 == _T_908 ? _T_38 : _GEN_8017; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8019 = 6'h13 == _T_908 ? _T_39 : _GEN_8018; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8020 = 6'h14 == _T_908 ? _T_40 : _GEN_8019; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8021 = 6'h15 == _T_908 ? _T_41 : _GEN_8020; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8022 = 6'h16 == _T_908 ? _T_42 : _GEN_8021; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8023 = 6'h17 == _T_908 ? _T_43 : _GEN_8022; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8024 = 6'h18 == _T_908 ? _T_44 : _GEN_8023; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8025 = 6'h19 == _T_908 ? _T_45 : _GEN_8024; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8026 = 6'h1a == _T_908 ? _T_46 : _GEN_8025; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8027 = 6'h1b == _T_908 ? _T_47 : _GEN_8026; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8028 = 6'h1c == _T_908 ? _T_48 : _GEN_8027; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8029 = 6'h1d == _T_908 ? _T_49 : _GEN_8028; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8030 = 6'h1e == _T_908 ? _T_50 : _GEN_8029; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8031 = 6'h1f == _T_908 ? _T_51 : _GEN_8030; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8032 = 6'h20 == _T_908 ? _T_52 : _GEN_8031; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8033 = 6'h21 == _T_908 ? _T_53 : _GEN_8032; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8034 = 6'h22 == _T_908 ? _T_54 : _GEN_8033; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8035 = 6'h23 == _T_908 ? _T_55 : _GEN_8034; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8036 = 6'h24 == _T_908 ? _T_56 : _GEN_8035; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8037 = 6'h25 == _T_908 ? _T_57 : _GEN_8036; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8038 = 6'h26 == _T_908 ? _T_58 : _GEN_8037; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8039 = 6'h27 == _T_908 ? _T_59 : _GEN_8038; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8040 = 6'h28 == _T_908 ? _T_60 : _GEN_8039; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8041 = 6'h29 == _T_908 ? _T_61 : _GEN_8040; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8042 = 6'h2a == _T_908 ? _T_62 : _GEN_8041; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8043 = 6'h2b == _T_908 ? _T_63 : _GEN_8042; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8044 = 6'h2c == _T_908 ? _T_64 : _GEN_8043; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8045 = 6'h2d == _T_908 ? _T_65 : _GEN_8044; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8046 = 6'h2e == _T_908 ? _T_66 : _GEN_8045; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8047 = 6'h2f == _T_908 ? _T_67 : _GEN_8046; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8048 = 6'h30 == _T_908 ? _T_68 : _GEN_8047; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8049 = 6'h31 == _T_908 ? _T_69 : _GEN_8048; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8050 = 6'h32 == _T_908 ? _T_70 : _GEN_8049; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8051 = 6'h33 == _T_908 ? _T_71 : _GEN_8050; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8052 = 6'h34 == _T_908 ? _T_72 : _GEN_8051; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8053 = 6'h35 == _T_908 ? _T_73 : _GEN_8052; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8054 = 6'h36 == _T_908 ? _T_74 : _GEN_8053; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8055 = 6'h37 == _T_908 ? _T_75 : _GEN_8054; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8056 = 6'h38 == _T_908 ? _T_76 : _GEN_8055; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8057 = 6'h39 == _T_908 ? _T_77 : _GEN_8056; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8058 = 6'h3a == _T_908 ? _T_78 : _GEN_8057; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8059 = 6'h3b == _T_908 ? _T_79 : _GEN_8058; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8060 = 6'h3c == _T_908 ? _T_80 : _GEN_8059; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8061 = 6'h3d == _T_908 ? _T_81 : _GEN_8060; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8062 = 6'h3e == _T_908 ? _T_82 : _GEN_8061; // @[execute.scala 79:10:@2291.4]
  assign _GEN_8063 = 6'h3f == _T_908 ? _T_83 : _GEN_8062; // @[execute.scala 79:10:@2291.4]
  assign _T_910 = _T_900 ? _GEN_7999 : _GEN_8063; // @[execute.scala 79:10:@2291.4]
  assign _T_912 = io_amount < 6'h1; // @[execute.scala 79:15:@2292.4]
  assign _T_914 = io_amount - 6'h1; // @[execute.scala 79:37:@2293.4]
  assign _T_915 = $unsigned(_T_914); // @[execute.scala 79:37:@2294.4]
  assign _T_916 = _T_915[5:0]; // @[execute.scala 79:37:@2295.4]
  assign _T_919 = 6'h3f + io_amount; // @[execute.scala 79:60:@2296.4]
  assign _T_920 = 6'h3f + io_amount; // @[execute.scala 79:60:@2297.4]
  assign _GEN_8065 = 6'h1 == _T_916 ? _T_21 : _T_20; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8066 = 6'h2 == _T_916 ? _T_22 : _GEN_8065; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8067 = 6'h3 == _T_916 ? _T_23 : _GEN_8066; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8068 = 6'h4 == _T_916 ? _T_24 : _GEN_8067; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8069 = 6'h5 == _T_916 ? _T_25 : _GEN_8068; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8070 = 6'h6 == _T_916 ? _T_26 : _GEN_8069; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8071 = 6'h7 == _T_916 ? _T_27 : _GEN_8070; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8072 = 6'h8 == _T_916 ? _T_28 : _GEN_8071; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8073 = 6'h9 == _T_916 ? _T_29 : _GEN_8072; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8074 = 6'ha == _T_916 ? _T_30 : _GEN_8073; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8075 = 6'hb == _T_916 ? _T_31 : _GEN_8074; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8076 = 6'hc == _T_916 ? _T_32 : _GEN_8075; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8077 = 6'hd == _T_916 ? _T_33 : _GEN_8076; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8078 = 6'he == _T_916 ? _T_34 : _GEN_8077; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8079 = 6'hf == _T_916 ? _T_35 : _GEN_8078; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8080 = 6'h10 == _T_916 ? _T_36 : _GEN_8079; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8081 = 6'h11 == _T_916 ? _T_37 : _GEN_8080; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8082 = 6'h12 == _T_916 ? _T_38 : _GEN_8081; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8083 = 6'h13 == _T_916 ? _T_39 : _GEN_8082; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8084 = 6'h14 == _T_916 ? _T_40 : _GEN_8083; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8085 = 6'h15 == _T_916 ? _T_41 : _GEN_8084; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8086 = 6'h16 == _T_916 ? _T_42 : _GEN_8085; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8087 = 6'h17 == _T_916 ? _T_43 : _GEN_8086; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8088 = 6'h18 == _T_916 ? _T_44 : _GEN_8087; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8089 = 6'h19 == _T_916 ? _T_45 : _GEN_8088; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8090 = 6'h1a == _T_916 ? _T_46 : _GEN_8089; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8091 = 6'h1b == _T_916 ? _T_47 : _GEN_8090; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8092 = 6'h1c == _T_916 ? _T_48 : _GEN_8091; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8093 = 6'h1d == _T_916 ? _T_49 : _GEN_8092; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8094 = 6'h1e == _T_916 ? _T_50 : _GEN_8093; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8095 = 6'h1f == _T_916 ? _T_51 : _GEN_8094; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8096 = 6'h20 == _T_916 ? _T_52 : _GEN_8095; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8097 = 6'h21 == _T_916 ? _T_53 : _GEN_8096; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8098 = 6'h22 == _T_916 ? _T_54 : _GEN_8097; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8099 = 6'h23 == _T_916 ? _T_55 : _GEN_8098; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8100 = 6'h24 == _T_916 ? _T_56 : _GEN_8099; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8101 = 6'h25 == _T_916 ? _T_57 : _GEN_8100; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8102 = 6'h26 == _T_916 ? _T_58 : _GEN_8101; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8103 = 6'h27 == _T_916 ? _T_59 : _GEN_8102; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8104 = 6'h28 == _T_916 ? _T_60 : _GEN_8103; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8105 = 6'h29 == _T_916 ? _T_61 : _GEN_8104; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8106 = 6'h2a == _T_916 ? _T_62 : _GEN_8105; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8107 = 6'h2b == _T_916 ? _T_63 : _GEN_8106; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8108 = 6'h2c == _T_916 ? _T_64 : _GEN_8107; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8109 = 6'h2d == _T_916 ? _T_65 : _GEN_8108; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8110 = 6'h2e == _T_916 ? _T_66 : _GEN_8109; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8111 = 6'h2f == _T_916 ? _T_67 : _GEN_8110; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8112 = 6'h30 == _T_916 ? _T_68 : _GEN_8111; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8113 = 6'h31 == _T_916 ? _T_69 : _GEN_8112; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8114 = 6'h32 == _T_916 ? _T_70 : _GEN_8113; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8115 = 6'h33 == _T_916 ? _T_71 : _GEN_8114; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8116 = 6'h34 == _T_916 ? _T_72 : _GEN_8115; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8117 = 6'h35 == _T_916 ? _T_73 : _GEN_8116; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8118 = 6'h36 == _T_916 ? _T_74 : _GEN_8117; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8119 = 6'h37 == _T_916 ? _T_75 : _GEN_8118; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8120 = 6'h38 == _T_916 ? _T_76 : _GEN_8119; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8121 = 6'h39 == _T_916 ? _T_77 : _GEN_8120; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8122 = 6'h3a == _T_916 ? _T_78 : _GEN_8121; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8123 = 6'h3b == _T_916 ? _T_79 : _GEN_8122; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8124 = 6'h3c == _T_916 ? _T_80 : _GEN_8123; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8125 = 6'h3d == _T_916 ? _T_81 : _GEN_8124; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8126 = 6'h3e == _T_916 ? _T_82 : _GEN_8125; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8127 = 6'h3f == _T_916 ? _T_83 : _GEN_8126; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8129 = 6'h1 == _T_920 ? _T_21 : _T_20; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8130 = 6'h2 == _T_920 ? _T_22 : _GEN_8129; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8131 = 6'h3 == _T_920 ? _T_23 : _GEN_8130; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8132 = 6'h4 == _T_920 ? _T_24 : _GEN_8131; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8133 = 6'h5 == _T_920 ? _T_25 : _GEN_8132; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8134 = 6'h6 == _T_920 ? _T_26 : _GEN_8133; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8135 = 6'h7 == _T_920 ? _T_27 : _GEN_8134; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8136 = 6'h8 == _T_920 ? _T_28 : _GEN_8135; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8137 = 6'h9 == _T_920 ? _T_29 : _GEN_8136; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8138 = 6'ha == _T_920 ? _T_30 : _GEN_8137; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8139 = 6'hb == _T_920 ? _T_31 : _GEN_8138; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8140 = 6'hc == _T_920 ? _T_32 : _GEN_8139; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8141 = 6'hd == _T_920 ? _T_33 : _GEN_8140; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8142 = 6'he == _T_920 ? _T_34 : _GEN_8141; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8143 = 6'hf == _T_920 ? _T_35 : _GEN_8142; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8144 = 6'h10 == _T_920 ? _T_36 : _GEN_8143; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8145 = 6'h11 == _T_920 ? _T_37 : _GEN_8144; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8146 = 6'h12 == _T_920 ? _T_38 : _GEN_8145; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8147 = 6'h13 == _T_920 ? _T_39 : _GEN_8146; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8148 = 6'h14 == _T_920 ? _T_40 : _GEN_8147; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8149 = 6'h15 == _T_920 ? _T_41 : _GEN_8148; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8150 = 6'h16 == _T_920 ? _T_42 : _GEN_8149; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8151 = 6'h17 == _T_920 ? _T_43 : _GEN_8150; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8152 = 6'h18 == _T_920 ? _T_44 : _GEN_8151; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8153 = 6'h19 == _T_920 ? _T_45 : _GEN_8152; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8154 = 6'h1a == _T_920 ? _T_46 : _GEN_8153; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8155 = 6'h1b == _T_920 ? _T_47 : _GEN_8154; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8156 = 6'h1c == _T_920 ? _T_48 : _GEN_8155; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8157 = 6'h1d == _T_920 ? _T_49 : _GEN_8156; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8158 = 6'h1e == _T_920 ? _T_50 : _GEN_8157; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8159 = 6'h1f == _T_920 ? _T_51 : _GEN_8158; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8160 = 6'h20 == _T_920 ? _T_52 : _GEN_8159; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8161 = 6'h21 == _T_920 ? _T_53 : _GEN_8160; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8162 = 6'h22 == _T_920 ? _T_54 : _GEN_8161; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8163 = 6'h23 == _T_920 ? _T_55 : _GEN_8162; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8164 = 6'h24 == _T_920 ? _T_56 : _GEN_8163; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8165 = 6'h25 == _T_920 ? _T_57 : _GEN_8164; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8166 = 6'h26 == _T_920 ? _T_58 : _GEN_8165; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8167 = 6'h27 == _T_920 ? _T_59 : _GEN_8166; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8168 = 6'h28 == _T_920 ? _T_60 : _GEN_8167; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8169 = 6'h29 == _T_920 ? _T_61 : _GEN_8168; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8170 = 6'h2a == _T_920 ? _T_62 : _GEN_8169; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8171 = 6'h2b == _T_920 ? _T_63 : _GEN_8170; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8172 = 6'h2c == _T_920 ? _T_64 : _GEN_8171; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8173 = 6'h2d == _T_920 ? _T_65 : _GEN_8172; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8174 = 6'h2e == _T_920 ? _T_66 : _GEN_8173; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8175 = 6'h2f == _T_920 ? _T_67 : _GEN_8174; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8176 = 6'h30 == _T_920 ? _T_68 : _GEN_8175; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8177 = 6'h31 == _T_920 ? _T_69 : _GEN_8176; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8178 = 6'h32 == _T_920 ? _T_70 : _GEN_8177; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8179 = 6'h33 == _T_920 ? _T_71 : _GEN_8178; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8180 = 6'h34 == _T_920 ? _T_72 : _GEN_8179; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8181 = 6'h35 == _T_920 ? _T_73 : _GEN_8180; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8182 = 6'h36 == _T_920 ? _T_74 : _GEN_8181; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8183 = 6'h37 == _T_920 ? _T_75 : _GEN_8182; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8184 = 6'h38 == _T_920 ? _T_76 : _GEN_8183; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8185 = 6'h39 == _T_920 ? _T_77 : _GEN_8184; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8186 = 6'h3a == _T_920 ? _T_78 : _GEN_8185; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8187 = 6'h3b == _T_920 ? _T_79 : _GEN_8186; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8188 = 6'h3c == _T_920 ? _T_80 : _GEN_8187; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8189 = 6'h3d == _T_920 ? _T_81 : _GEN_8188; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8190 = 6'h3e == _T_920 ? _T_82 : _GEN_8189; // @[execute.scala 79:10:@2298.4]
  assign _GEN_8191 = 6'h3f == _T_920 ? _T_83 : _GEN_8190; // @[execute.scala 79:10:@2298.4]
  assign _T_922 = _T_912 ? _GEN_8127 : _GEN_8191; // @[execute.scala 79:10:@2298.4]
  assign _T_999 = {_T_250,_T_238,_T_226,_T_214,_T_202,_T_190,_T_178,_GEN_63}; // @[execute.scala 89:73:@2370.4]
  assign _T_1007 = {_T_346,_T_334,_T_322,_T_310,_T_298,_T_286,_T_274,_T_262,_T_999}; // @[execute.scala 89:73:@2378.4]
  assign _T_1014 = {_T_442,_T_430,_T_418,_T_406,_T_394,_T_382,_T_370,_T_358}; // @[execute.scala 89:73:@2385.4]
  assign _T_1023 = {_T_538,_T_526,_T_514,_T_502,_T_490,_T_478,_T_466,_T_454,_T_1014,_T_1007}; // @[execute.scala 89:73:@2394.4]
  assign _T_1030 = {_T_634,_T_622,_T_610,_T_598,_T_586,_T_574,_T_562,_T_550}; // @[execute.scala 89:73:@2401.4]
  assign _T_1038 = {_T_730,_T_718,_T_706,_T_694,_T_682,_T_670,_T_658,_T_646,_T_1030}; // @[execute.scala 89:73:@2409.4]
  assign _T_1045 = {_T_826,_T_814,_T_802,_T_790,_T_778,_T_766,_T_754,_T_742}; // @[execute.scala 89:73:@2416.4]
  assign _T_1054 = {_T_922,_T_910,_T_898,_T_886,_T_874,_T_862,_T_850,_T_838,_T_1045,_T_1038}; // @[execute.scala 89:73:@2425.4]
  assign _T_1055 = {_T_1054,_T_1023}; // @[execute.scala 89:73:@2426.4]
  assign _T_1056 = 2'h3 == io_opcode; // @[Mux.scala 46:19:@2427.4]
  assign _T_1057 = _T_1056 ? _T_1055 : io_word; // @[Mux.scala 46:16:@2428.4]
  assign _T_1058 = 2'h2 == io_opcode; // @[Mux.scala 46:19:@2429.4]
  assign _T_1059 = _T_1058 ? _T_19 : _T_1057; // @[Mux.scala 46:16:@2430.4]
  assign _T_1060 = 2'h1 == io_opcode; // @[Mux.scala 46:19:@2431.4]
  assign _T_1061 = _T_1060 ? _T_16 : _T_1059; // @[Mux.scala 46:16:@2432.4]
  assign _T_1062 = 2'h0 == io_opcode; // @[Mux.scala 46:19:@2433.4]
  assign res = _T_1062 ? _T_15 : {{63'd0}, _T_1061}; // @[Mux.scala 46:16:@2434.4]
  assign io_res = res[63:0]; // @[execute.scala 93:10:@2438.4]
endmodule
