module DecodeUnit( // @[:@625.2]
  input  [31:0] io_finst_inst, // @[:@628.4]
  input         io_finst_tag, // @[:@628.4]
  input  [63:0] io_finst_pc, // @[:@628.4]
  output        io_dinst_rd_valid, // @[:@628.4]
  output [4:0]  io_dinst_rd_bits, // @[:@628.4]
  output [4:0]  io_dinst_rs1_bits, // @[:@628.4]
  output        io_dinst_rs2_valid, // @[:@628.4]
  output [4:0]  io_dinst_rs2_bits, // @[:@628.4]
  output [25:0] io_dinst_imm_bits, // @[:@628.4]
  output        io_dinst_shift_val_valid, // @[:@628.4]
  output [5:0]  io_dinst_shift_val_bits, // @[:@628.4]
  output [1:0]  io_dinst_shift_type, // @[:@628.4]
  output [3:0]  io_dinst_cond_bits, // @[:@628.4]
  output [2:0]  io_dinst_itype, // @[:@628.4]
  output [2:0]  io_dinst_op, // @[:@628.4]
  output        io_dinst_nzcv_en, // @[:@628.4]
  output        io_dinst_tag, // @[:@628.4]
  output [63:0] io_dinst_pc // @[:@628.4]
);
  wire [7:0] _T_117; // @[decode.scala 121:33:@630.4]
  wire [7:0] _T_118; // @[decode.scala 121:44:@631.4]
  wire [7:0] _T_119; // @[decode.scala 121:56:@632.4]
  wire [7:0] _T_120; // @[decode.scala 121:69:@633.4]
  wire [31:0] instBE; // @[Cat.scala 30:58:@636.4]
  wire [31:0] _T_210; // @[Lookup.scala 9:38:@681.4]
  wire  _T_211; // @[Lookup.scala 9:38:@682.4]
  wire  _T_215; // @[Lookup.scala 9:38:@684.4]
  wire  _T_219; // @[Lookup.scala 9:38:@686.4]
  wire  _T_223; // @[Lookup.scala 9:38:@688.4]
  wire  _T_227; // @[Lookup.scala 9:38:@690.4]
  wire  _T_231; // @[Lookup.scala 9:38:@692.4]
  wire  _T_235; // @[Lookup.scala 9:38:@694.4]
  wire  _T_239; // @[Lookup.scala 9:38:@696.4]
  wire [31:0] _T_242; // @[Lookup.scala 9:38:@697.4]
  wire  _T_243; // @[Lookup.scala 9:38:@698.4]
  wire  _T_247; // @[Lookup.scala 9:38:@700.4]
  wire [31:0] _T_250; // @[Lookup.scala 9:38:@701.4]
  wire  _T_251; // @[Lookup.scala 9:38:@702.4]
  wire [31:0] _T_254; // @[Lookup.scala 9:38:@703.4]
  wire  _T_255; // @[Lookup.scala 9:38:@704.4]
  wire  _T_259; // @[Lookup.scala 9:38:@706.4]
  wire  _T_263; // @[Lookup.scala 9:38:@708.4]
  wire  _T_267; // @[Lookup.scala 9:38:@710.4]
  wire [31:0] _T_270; // @[Lookup.scala 9:38:@711.4]
  wire  _T_271; // @[Lookup.scala 9:38:@712.4]
  wire [2:0] _T_272; // @[Lookup.scala 11:37:@713.4]
  wire [2:0] _T_273; // @[Lookup.scala 11:37:@714.4]
  wire [2:0] _T_274; // @[Lookup.scala 11:37:@715.4]
  wire [2:0] _T_275; // @[Lookup.scala 11:37:@716.4]
  wire [2:0] _T_276; // @[Lookup.scala 11:37:@717.4]
  wire [2:0] _T_277; // @[Lookup.scala 11:37:@718.4]
  wire [2:0] _T_278; // @[Lookup.scala 11:37:@719.4]
  wire [2:0] _T_279; // @[Lookup.scala 11:37:@720.4]
  wire [2:0] _T_280; // @[Lookup.scala 11:37:@721.4]
  wire [2:0] _T_281; // @[Lookup.scala 11:37:@722.4]
  wire [2:0] _T_282; // @[Lookup.scala 11:37:@723.4]
  wire [2:0] _T_283; // @[Lookup.scala 11:37:@724.4]
  wire [2:0] _T_284; // @[Lookup.scala 11:37:@725.4]
  wire [2:0] _T_285; // @[Lookup.scala 11:37:@726.4]
  wire [2:0] _T_286; // @[Lookup.scala 11:37:@727.4]
  wire [2:0] dinst_itype; // @[Lookup.scala 11:37:@728.4]
  wire [2:0] _T_289; // @[Lookup.scala 11:37:@730.4]
  wire [2:0] _T_290; // @[Lookup.scala 11:37:@731.4]
  wire [2:0] _T_291; // @[Lookup.scala 11:37:@732.4]
  wire [2:0] _T_292; // @[Lookup.scala 11:37:@733.4]
  wire [2:0] _T_293; // @[Lookup.scala 11:37:@734.4]
  wire [2:0] _T_294; // @[Lookup.scala 11:37:@735.4]
  wire [2:0] _T_295; // @[Lookup.scala 11:37:@736.4]
  wire [2:0] _T_296; // @[Lookup.scala 11:37:@737.4]
  wire [2:0] _T_297; // @[Lookup.scala 11:37:@738.4]
  wire [2:0] _T_298; // @[Lookup.scala 11:37:@739.4]
  wire [2:0] _T_299; // @[Lookup.scala 11:37:@740.4]
  wire [2:0] _T_300; // @[Lookup.scala 11:37:@741.4]
  wire [2:0] _T_301; // @[Lookup.scala 11:37:@742.4]
  wire [2:0] _T_302; // @[Lookup.scala 11:37:@743.4]
  wire  _T_305; // @[Lookup.scala 11:37:@746.4]
  wire  _T_306; // @[Lookup.scala 11:37:@747.4]
  wire  _T_307; // @[Lookup.scala 11:37:@748.4]
  wire  _T_308; // @[Lookup.scala 11:37:@749.4]
  wire  _T_309; // @[Lookup.scala 11:37:@750.4]
  wire  _T_310; // @[Lookup.scala 11:37:@751.4]
  wire  _T_311; // @[Lookup.scala 11:37:@752.4]
  wire  _T_312; // @[Lookup.scala 11:37:@753.4]
  wire  _T_313; // @[Lookup.scala 11:37:@754.4]
  wire  _T_314; // @[Lookup.scala 11:37:@755.4]
  wire  _T_315; // @[Lookup.scala 11:37:@756.4]
  wire  _T_316; // @[Lookup.scala 11:37:@757.4]
  wire  _T_317; // @[Lookup.scala 11:37:@758.4]
  wire  _T_318; // @[Lookup.scala 11:37:@759.4]
  wire  _T_322; // @[Lookup.scala 11:37:@763.4]
  wire  _T_323; // @[Lookup.scala 11:37:@764.4]
  wire  _T_324; // @[Lookup.scala 11:37:@765.4]
  wire  _T_325; // @[Lookup.scala 11:37:@766.4]
  wire  _T_326; // @[Lookup.scala 11:37:@767.4]
  wire  _T_327; // @[Lookup.scala 11:37:@768.4]
  wire  _T_328; // @[Lookup.scala 11:37:@769.4]
  wire  _T_329; // @[Lookup.scala 11:37:@770.4]
  wire  _T_330; // @[Lookup.scala 11:37:@771.4]
  wire  _T_331; // @[Lookup.scala 11:37:@772.4]
  wire  _T_332; // @[Lookup.scala 11:37:@773.4]
  wire  _T_333; // @[Lookup.scala 11:37:@774.4]
  wire  _T_334; // @[Lookup.scala 11:37:@775.4]
  wire  _T_345; // @[Lookup.scala 11:37:@786.4]
  wire  _T_346; // @[Lookup.scala 11:37:@787.4]
  wire  _T_347; // @[Lookup.scala 11:37:@788.4]
  wire  _T_348; // @[Lookup.scala 11:37:@789.4]
  wire  _T_349; // @[Lookup.scala 11:37:@790.4]
  wire  _T_350; // @[Lookup.scala 11:37:@791.4]
  wire  _T_402; // @[Lookup.scala 11:37:@843.4]
  wire  _T_403; // @[Lookup.scala 11:37:@844.4]
  wire  _T_404; // @[Lookup.scala 11:37:@845.4]
  wire  _T_405; // @[Lookup.scala 11:37:@846.4]
  wire  _T_406; // @[Lookup.scala 11:37:@847.4]
  wire  _T_407; // @[Lookup.scala 11:37:@848.4]
  wire  _T_408; // @[Lookup.scala 11:37:@849.4]
  wire  _T_409; // @[Lookup.scala 11:37:@850.4]
  wire  _T_410; // @[Lookup.scala 11:37:@851.4]
  wire  _T_411; // @[Lookup.scala 11:37:@852.4]
  wire  _T_412; // @[Lookup.scala 11:37:@853.4]
  wire  _T_413; // @[Lookup.scala 11:37:@854.4]
  wire  _T_414; // @[Lookup.scala 11:37:@855.4]
  wire [4:0] _T_432; // @[decode.scala 39:64:@873.4]
  wire  _T_435; // @[Mux.scala 46:19:@876.4]
  wire [4:0] _T_436; // @[Mux.scala 46:16:@877.4]
  wire  _T_437; // @[Mux.scala 46:19:@878.4]
  wire [4:0] _T_438; // @[Mux.scala 46:16:@879.4]
  wire  _T_439; // @[Mux.scala 46:19:@880.4]
  wire [4:0] _T_441; // @[decode.scala 42:65:@883.4]
  wire [4:0] _T_444; // @[Mux.scala 46:16:@886.4]
  wire [4:0] _T_447; // @[decode.scala 44:65:@890.4]
  wire [5:0] _T_450; // @[decode.scala 45:65:@894.4]
  wire [25:0] _T_451; // @[decode.scala 46:62:@895.4]
  wire [18:0] _T_452; // @[decode.scala 47:62:@896.4]
  wire [11:0] _T_453; // @[decode.scala 48:62:@897.4]
  wire [25:0] _T_456; // @[Mux.scala 46:16:@900.4]
  wire [25:0] _T_458; // @[Mux.scala 46:16:@902.4]
  wire  _T_459; // @[Mux.scala 46:19:@903.4]
  wire [25:0] _T_460; // @[Mux.scala 46:16:@904.4]
  wire  _T_461; // @[Mux.scala 46:19:@905.4]
  wire [25:0] _T_462; // @[Mux.scala 46:16:@906.4]
  wire [25:0] dinst_imm_bits; // @[Mux.scala 46:16:@908.4]
  wire  _T_465; // @[decode.scala 51:54:@910.4]
  wire [3:0] _T_468; // @[decode.scala 51:49:@911.4]
  wire [25:0] _T_470; // @[Mux.scala 46:16:@913.4]
  wire [25:0] _T_472; // @[Mux.scala 46:16:@915.4]
  wire [1:0] _T_473; // @[decode.scala 53:72:@917.4]
  wire [1:0] _T_476; // @[Mux.scala 46:16:@920.4]
  wire [3:0] _T_479; // @[decode.scala 55:66:@924.4]
  assign _T_117 = io_finst_inst[7:0]; // @[decode.scala 121:33:@630.4]
  assign _T_118 = io_finst_inst[15:8]; // @[decode.scala 121:44:@631.4]
  assign _T_119 = io_finst_inst[23:16]; // @[decode.scala 121:56:@632.4]
  assign _T_120 = io_finst_inst[31:24]; // @[decode.scala 121:69:@633.4]
  assign instBE = {_T_117,_T_118,_T_119,_T_120}; // @[Cat.scala 30:58:@636.4]
  assign _T_210 = instBE & 32'hff200000; // @[Lookup.scala 9:38:@681.4]
  assign _T_211 = 32'h8a000000 == _T_210; // @[Lookup.scala 9:38:@682.4]
  assign _T_215 = 32'h8a200000 == _T_210; // @[Lookup.scala 9:38:@684.4]
  assign _T_219 = 32'haa000000 == _T_210; // @[Lookup.scala 9:38:@686.4]
  assign _T_223 = 32'haa200000 == _T_210; // @[Lookup.scala 9:38:@688.4]
  assign _T_227 = 32'hca000000 == _T_210; // @[Lookup.scala 9:38:@690.4]
  assign _T_231 = 32'hca200000 == _T_210; // @[Lookup.scala 9:38:@692.4]
  assign _T_235 = 32'hea000000 == _T_210; // @[Lookup.scala 9:38:@694.4]
  assign _T_239 = 32'hea200000 == _T_210; // @[Lookup.scala 9:38:@696.4]
  assign _T_242 = instBE & 32'hfc000000; // @[Lookup.scala 9:38:@697.4]
  assign _T_243 = 32'h14000000 == _T_242; // @[Lookup.scala 9:38:@698.4]
  assign _T_247 = 32'h94000000 == _T_242; // @[Lookup.scala 9:38:@700.4]
  assign _T_250 = instBE & 32'hff000010; // @[Lookup.scala 9:38:@701.4]
  assign _T_251 = 32'h54000000 == _T_250; // @[Lookup.scala 9:38:@702.4]
  assign _T_254 = instBE & 32'hff800000; // @[Lookup.scala 9:38:@703.4]
  assign _T_255 = 32'h91000000 == _T_254; // @[Lookup.scala 9:38:@704.4]
  assign _T_259 = 32'hb1000000 == _T_254; // @[Lookup.scala 9:38:@706.4]
  assign _T_263 = 32'hd1000000 == _T_254; // @[Lookup.scala 9:38:@708.4]
  assign _T_267 = 32'hf1000000 == _T_254; // @[Lookup.scala 9:38:@710.4]
  assign _T_270 = instBE & 32'hff000000; // @[Lookup.scala 9:38:@711.4]
  assign _T_271 = 32'h58000000 == _T_270; // @[Lookup.scala 9:38:@712.4]
  assign _T_272 = _T_271 ? 3'h5 : 3'h0; // @[Lookup.scala 11:37:@713.4]
  assign _T_273 = _T_267 ? 3'h4 : _T_272; // @[Lookup.scala 11:37:@714.4]
  assign _T_274 = _T_263 ? 3'h4 : _T_273; // @[Lookup.scala 11:37:@715.4]
  assign _T_275 = _T_259 ? 3'h4 : _T_274; // @[Lookup.scala 11:37:@716.4]
  assign _T_276 = _T_255 ? 3'h4 : _T_275; // @[Lookup.scala 11:37:@717.4]
  assign _T_277 = _T_251 ? 3'h3 : _T_276; // @[Lookup.scala 11:37:@718.4]
  assign _T_278 = _T_247 ? 3'h2 : _T_277; // @[Lookup.scala 11:37:@719.4]
  assign _T_279 = _T_243 ? 3'h2 : _T_278; // @[Lookup.scala 11:37:@720.4]
  assign _T_280 = _T_239 ? 3'h1 : _T_279; // @[Lookup.scala 11:37:@721.4]
  assign _T_281 = _T_235 ? 3'h1 : _T_280; // @[Lookup.scala 11:37:@722.4]
  assign _T_282 = _T_231 ? 3'h1 : _T_281; // @[Lookup.scala 11:37:@723.4]
  assign _T_283 = _T_227 ? 3'h1 : _T_282; // @[Lookup.scala 11:37:@724.4]
  assign _T_284 = _T_223 ? 3'h1 : _T_283; // @[Lookup.scala 11:37:@725.4]
  assign _T_285 = _T_219 ? 3'h1 : _T_284; // @[Lookup.scala 11:37:@726.4]
  assign _T_286 = _T_215 ? 3'h1 : _T_285; // @[Lookup.scala 11:37:@727.4]
  assign dinst_itype = _T_211 ? 3'h1 : _T_286; // @[Lookup.scala 11:37:@728.4]
  assign _T_289 = _T_267 ? 3'h7 : 3'h0; // @[Lookup.scala 11:37:@730.4]
  assign _T_290 = _T_263 ? 3'h7 : _T_289; // @[Lookup.scala 11:37:@731.4]
  assign _T_291 = _T_259 ? 3'h6 : _T_290; // @[Lookup.scala 11:37:@732.4]
  assign _T_292 = _T_255 ? 3'h6 : _T_291; // @[Lookup.scala 11:37:@733.4]
  assign _T_293 = _T_251 ? 3'h1 : _T_292; // @[Lookup.scala 11:37:@734.4]
  assign _T_294 = _T_247 ? 3'h0 : _T_293; // @[Lookup.scala 11:37:@735.4]
  assign _T_295 = _T_243 ? 3'h0 : _T_294; // @[Lookup.scala 11:37:@736.4]
  assign _T_296 = _T_239 ? 3'h1 : _T_295; // @[Lookup.scala 11:37:@737.4]
  assign _T_297 = _T_235 ? 3'h0 : _T_296; // @[Lookup.scala 11:37:@738.4]
  assign _T_298 = _T_231 ? 3'h5 : _T_297; // @[Lookup.scala 11:37:@739.4]
  assign _T_299 = _T_227 ? 3'h4 : _T_298; // @[Lookup.scala 11:37:@740.4]
  assign _T_300 = _T_223 ? 3'h3 : _T_299; // @[Lookup.scala 11:37:@741.4]
  assign _T_301 = _T_219 ? 3'h2 : _T_300; // @[Lookup.scala 11:37:@742.4]
  assign _T_302 = _T_215 ? 3'h1 : _T_301; // @[Lookup.scala 11:37:@743.4]
  assign _T_305 = _T_267 ? 1'h1 : _T_271; // @[Lookup.scala 11:37:@746.4]
  assign _T_306 = _T_263 ? 1'h1 : _T_305; // @[Lookup.scala 11:37:@747.4]
  assign _T_307 = _T_259 ? 1'h1 : _T_306; // @[Lookup.scala 11:37:@748.4]
  assign _T_308 = _T_255 ? 1'h1 : _T_307; // @[Lookup.scala 11:37:@749.4]
  assign _T_309 = _T_251 ? 1'h0 : _T_308; // @[Lookup.scala 11:37:@750.4]
  assign _T_310 = _T_247 ? 1'h0 : _T_309; // @[Lookup.scala 11:37:@751.4]
  assign _T_311 = _T_243 ? 1'h0 : _T_310; // @[Lookup.scala 11:37:@752.4]
  assign _T_312 = _T_239 ? 1'h1 : _T_311; // @[Lookup.scala 11:37:@753.4]
  assign _T_313 = _T_235 ? 1'h1 : _T_312; // @[Lookup.scala 11:37:@754.4]
  assign _T_314 = _T_231 ? 1'h1 : _T_313; // @[Lookup.scala 11:37:@755.4]
  assign _T_315 = _T_227 ? 1'h1 : _T_314; // @[Lookup.scala 11:37:@756.4]
  assign _T_316 = _T_223 ? 1'h1 : _T_315; // @[Lookup.scala 11:37:@757.4]
  assign _T_317 = _T_219 ? 1'h1 : _T_316; // @[Lookup.scala 11:37:@758.4]
  assign _T_318 = _T_215 ? 1'h1 : _T_317; // @[Lookup.scala 11:37:@759.4]
  assign _T_322 = _T_263 ? 1'h1 : _T_267; // @[Lookup.scala 11:37:@763.4]
  assign _T_323 = _T_259 ? 1'h1 : _T_322; // @[Lookup.scala 11:37:@764.4]
  assign _T_324 = _T_255 ? 1'h1 : _T_323; // @[Lookup.scala 11:37:@765.4]
  assign _T_325 = _T_251 ? 1'h0 : _T_324; // @[Lookup.scala 11:37:@766.4]
  assign _T_326 = _T_247 ? 1'h0 : _T_325; // @[Lookup.scala 11:37:@767.4]
  assign _T_327 = _T_243 ? 1'h0 : _T_326; // @[Lookup.scala 11:37:@768.4]
  assign _T_328 = _T_239 ? 1'h1 : _T_327; // @[Lookup.scala 11:37:@769.4]
  assign _T_329 = _T_235 ? 1'h1 : _T_328; // @[Lookup.scala 11:37:@770.4]
  assign _T_330 = _T_231 ? 1'h1 : _T_329; // @[Lookup.scala 11:37:@771.4]
  assign _T_331 = _T_227 ? 1'h1 : _T_330; // @[Lookup.scala 11:37:@772.4]
  assign _T_332 = _T_223 ? 1'h1 : _T_331; // @[Lookup.scala 11:37:@773.4]
  assign _T_333 = _T_219 ? 1'h1 : _T_332; // @[Lookup.scala 11:37:@774.4]
  assign _T_334 = _T_215 ? 1'h1 : _T_333; // @[Lookup.scala 11:37:@775.4]
  assign _T_345 = _T_235 ? 1'h1 : _T_239; // @[Lookup.scala 11:37:@786.4]
  assign _T_346 = _T_231 ? 1'h1 : _T_345; // @[Lookup.scala 11:37:@787.4]
  assign _T_347 = _T_227 ? 1'h1 : _T_346; // @[Lookup.scala 11:37:@788.4]
  assign _T_348 = _T_223 ? 1'h1 : _T_347; // @[Lookup.scala 11:37:@789.4]
  assign _T_349 = _T_219 ? 1'h1 : _T_348; // @[Lookup.scala 11:37:@790.4]
  assign _T_350 = _T_215 ? 1'h1 : _T_349; // @[Lookup.scala 11:37:@791.4]
  assign _T_402 = _T_263 ? 1'h0 : _T_267; // @[Lookup.scala 11:37:@843.4]
  assign _T_403 = _T_259 ? 1'h1 : _T_402; // @[Lookup.scala 11:37:@844.4]
  assign _T_404 = _T_255 ? 1'h0 : _T_403; // @[Lookup.scala 11:37:@845.4]
  assign _T_405 = _T_251 ? 1'h0 : _T_404; // @[Lookup.scala 11:37:@846.4]
  assign _T_406 = _T_247 ? 1'h0 : _T_405; // @[Lookup.scala 11:37:@847.4]
  assign _T_407 = _T_243 ? 1'h0 : _T_406; // @[Lookup.scala 11:37:@848.4]
  assign _T_408 = _T_239 ? 1'h1 : _T_407; // @[Lookup.scala 11:37:@849.4]
  assign _T_409 = _T_235 ? 1'h1 : _T_408; // @[Lookup.scala 11:37:@850.4]
  assign _T_410 = _T_231 ? 1'h0 : _T_409; // @[Lookup.scala 11:37:@851.4]
  assign _T_411 = _T_227 ? 1'h0 : _T_410; // @[Lookup.scala 11:37:@852.4]
  assign _T_412 = _T_223 ? 1'h0 : _T_411; // @[Lookup.scala 11:37:@853.4]
  assign _T_413 = _T_219 ? 1'h0 : _T_412; // @[Lookup.scala 11:37:@854.4]
  assign _T_414 = _T_215 ? 1'h0 : _T_413; // @[Lookup.scala 11:37:@855.4]
  assign _T_432 = instBE[4:0]; // @[decode.scala 39:64:@873.4]
  assign _T_435 = 3'h5 == dinst_itype; // @[Mux.scala 46:19:@876.4]
  assign _T_436 = _T_435 ? _T_432 : 5'h0; // @[Mux.scala 46:16:@877.4]
  assign _T_437 = 3'h4 == dinst_itype; // @[Mux.scala 46:19:@878.4]
  assign _T_438 = _T_437 ? _T_432 : _T_436; // @[Mux.scala 46:16:@879.4]
  assign _T_439 = 3'h1 == dinst_itype; // @[Mux.scala 46:19:@880.4]
  assign _T_441 = instBE[9:5]; // @[decode.scala 42:65:@883.4]
  assign _T_444 = _T_437 ? _T_441 : 5'h0; // @[Mux.scala 46:16:@886.4]
  assign _T_447 = instBE[20:16]; // @[decode.scala 44:65:@890.4]
  assign _T_450 = instBE[15:10]; // @[decode.scala 45:65:@894.4]
  assign _T_451 = instBE[25:0]; // @[decode.scala 46:62:@895.4]
  assign _T_452 = instBE[23:5]; // @[decode.scala 47:62:@896.4]
  assign _T_453 = instBE[21:10]; // @[decode.scala 48:62:@897.4]
  assign _T_456 = _T_435 ? {{7'd0}, _T_452} : 26'h0; // @[Mux.scala 46:16:@900.4]
  assign _T_458 = _T_437 ? {{14'd0}, _T_453} : _T_456; // @[Mux.scala 46:16:@902.4]
  assign _T_459 = 3'h3 == dinst_itype; // @[Mux.scala 46:19:@903.4]
  assign _T_460 = _T_459 ? {{7'd0}, _T_452} : _T_458; // @[Mux.scala 46:16:@904.4]
  assign _T_461 = 3'h2 == dinst_itype; // @[Mux.scala 46:19:@905.4]
  assign _T_462 = _T_461 ? _T_451 : _T_460; // @[Mux.scala 46:16:@906.4]
  assign dinst_imm_bits = _T_439 ? {{20'd0}, _T_450} : _T_462; // @[Mux.scala 46:16:@908.4]
  assign _T_465 = instBE[22]; // @[decode.scala 51:54:@910.4]
  assign _T_468 = _T_465 ? 4'hc : 4'h0; // @[decode.scala 51:49:@911.4]
  assign _T_470 = _T_439 ? dinst_imm_bits : 26'h0; // @[Mux.scala 46:16:@913.4]
  assign _T_472 = _T_437 ? {{22'd0}, _T_468} : _T_470; // @[Mux.scala 46:16:@915.4]
  assign _T_473 = instBE[23:22]; // @[decode.scala 53:72:@917.4]
  assign _T_476 = _T_437 ? _T_473 : 2'h0; // @[Mux.scala 46:16:@920.4]
  assign _T_479 = instBE[3:0]; // @[decode.scala 55:66:@924.4]
  assign io_dinst_rd_valid = _T_211 ? 1'h1 : _T_318; // @[decode.scala 125:12:@960.4]
  assign io_dinst_rd_bits = _T_439 ? _T_432 : _T_438; // @[decode.scala 125:12:@959.4]
  assign io_dinst_rs1_bits = _T_439 ? _T_441 : _T_444; // @[decode.scala 125:12:@957.4]
  assign io_dinst_rs2_valid = _T_211 ? 1'h1 : _T_350; // @[decode.scala 125:12:@956.4]
  assign io_dinst_rs2_bits = _T_439 ? _T_447 : 5'h0; // @[decode.scala 125:12:@955.4]
  assign io_dinst_imm_bits = _T_439 ? {{20'd0}, _T_450} : _T_462; // @[decode.scala 125:12:@953.4]
  assign io_dinst_shift_val_valid = _T_211 ? 1'h1 : _T_334; // @[decode.scala 125:12:@952.4]
  assign io_dinst_shift_val_bits = _T_472[5:0]; // @[decode.scala 125:12:@951.4]
  assign io_dinst_shift_type = _T_439 ? _T_473 : _T_476; // @[decode.scala 125:12:@950.4]
  assign io_dinst_cond_bits = _T_459 ? _T_479 : 4'h0; // @[decode.scala 125:12:@948.4]
  assign io_dinst_itype = _T_211 ? 3'h1 : _T_286; // @[decode.scala 125:12:@947.4]
  assign io_dinst_op = _T_211 ? 3'h0 : _T_302; // @[decode.scala 125:12:@946.4]
  assign io_dinst_nzcv_en = _T_211 ? 1'h0 : _T_414; // @[decode.scala 125:12:@945.4]
  assign io_dinst_tag = io_finst_tag; // @[decode.scala 125:12:@944.4]
  assign io_dinst_pc = io_finst_pc; // @[decode.scala 125:12:@941.4]
endmodule
