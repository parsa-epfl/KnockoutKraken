module ExtendReg(
  input  [63:0] io_value,
  input  [2:0]  io_option,
  input  [1:0]  io_shift,
  output [63:0] io_res
);
  wire  isSigned; // @[LoadStore.scala 52:27]
  wire [1:0] size; // @[LoadStore.scala 53:23]
  wire [7:0] _T_2; // @[LoadStore.scala 55:57]
  wire [63:0] _T_3; // @[LoadStore.scala 55:67]
  wire [15:0] _T_5; // @[LoadStore.scala 56:57]
  wire [63:0] _T_6; // @[LoadStore.scala 56:67]
  wire [31:0] _T_8; // @[LoadStore.scala 57:57]
  wire [63:0] _T_9; // @[LoadStore.scala 57:67]
  wire  _T_11; // @[Mux.scala 80:60]
  wire [63:0] _T_12; // @[Mux.scala 80:57]
  wire  _T_13; // @[Mux.scala 80:60]
  wire [63:0] _T_14; // @[Mux.scala 80:57]
  wire  _T_15; // @[Mux.scala 80:60]
  wire [63:0] _T_18; // @[LoadStore.scala 61:60]
  wire [63:0] _T_20; // @[LoadStore.scala 62:60]
  wire [63:0] _T_22; // @[LoadStore.scala 63:60]
  wire [63:0] _T_24; // @[Mux.scala 80:57]
  wire [63:0] _T_26; // @[Mux.scala 80:57]
  wire [63:0] valUExt; // @[Mux.scala 80:57]
  wire [63:0] _T_29; // @[LoadStore.scala 66:44]
  wire [63:0] res; // @[LoadStore.scala 66:25]
  wire [66:0] _GEN_0; // @[LoadStore.scala 67:17]
  wire [66:0] _T_31; // @[LoadStore.scala 67:17]
  assign isSigned = io_option[2]; // @[LoadStore.scala 52:27]
  assign size = io_option[1:0]; // @[LoadStore.scala 53:23]
  assign _T_2 = io_value[7:0]; // @[LoadStore.scala 55:57]
  assign _T_3 = {{56{_T_2[7]}},_T_2}; // @[LoadStore.scala 55:67]
  assign _T_5 = io_value[15:0]; // @[LoadStore.scala 56:57]
  assign _T_6 = {{48{_T_5[15]}},_T_5}; // @[LoadStore.scala 56:67]
  assign _T_8 = io_value[31:0]; // @[LoadStore.scala 57:57]
  assign _T_9 = {{32{_T_8[31]}},_T_8}; // @[LoadStore.scala 57:67]
  assign _T_11 = 2'h1 == size; // @[Mux.scala 80:60]
  assign _T_12 = _T_11 ? $signed(_T_6) : $signed(_T_3); // @[Mux.scala 80:57]
  assign _T_13 = 2'h2 == size; // @[Mux.scala 80:60]
  assign _T_14 = _T_13 ? $signed(_T_9) : $signed(_T_12); // @[Mux.scala 80:57]
  assign _T_15 = 2'h3 == size; // @[Mux.scala 80:60]
  assign _T_18 = {{56'd0}, io_value[7:0]}; // @[LoadStore.scala 61:60]
  assign _T_20 = {{48'd0}, io_value[15:0]}; // @[LoadStore.scala 62:60]
  assign _T_22 = {{32'd0}, io_value[31:0]}; // @[LoadStore.scala 63:60]
  assign _T_24 = _T_11 ? _T_20 : _T_18; // @[Mux.scala 80:57]
  assign _T_26 = _T_13 ? _T_22 : _T_24; // @[Mux.scala 80:57]
  assign valUExt = _T_15 ? io_value : _T_26; // @[Mux.scala 80:57]
  assign _T_29 = _T_15 ? $signed(io_value) : $signed(_T_14); // @[LoadStore.scala 66:44]
  assign res = isSigned ? _T_29 : valUExt; // @[LoadStore.scala 66:25]
  assign _GEN_0 = {{3'd0}, res}; // @[LoadStore.scala 67:17]
  assign _T_31 = _GEN_0 << io_shift; // @[LoadStore.scala 67:17]
  assign io_res = _T_31[63:0]; // @[LoadStore.scala 67:10]
endmodule
