module BasicALU( // @[:@2656.2]
  input  [63:0] io_a, // @[:@2659.4]
  input  [63:0] io_b, // @[:@2659.4]
  input  [2:0]  io_opcode, // @[:@2659.4]
  output [63:0] io_res, // @[:@2659.4]
  output [3:0]  io_nzcv // @[:@2659.4]
);
  wire [63:0] _T_16; // @[execute.scala 29:34:@2661.4]
  wire [63:0] _T_17; // @[execute.scala 30:36:@2662.4]
  wire [63:0] _T_18; // @[execute.scala 30:34:@2663.4]
  wire [63:0] _T_19; // @[execute.scala 31:34:@2664.4]
  wire [63:0] _T_21; // @[execute.scala 32:34:@2666.4]
  wire [63:0] _T_22; // @[execute.scala 33:34:@2667.4]
  wire [63:0] _T_24; // @[execute.scala 34:34:@2669.4]
  wire [64:0] _T_25; // @[execute.scala 35:34:@2670.4]
  wire [63:0] _T_26; // @[execute.scala 35:34:@2671.4]
  wire [64:0] _T_27; // @[execute.scala 36:34:@2672.4]
  wire [64:0] _T_28; // @[execute.scala 36:34:@2673.4]
  wire [63:0] _T_29; // @[execute.scala 36:34:@2674.4]
  wire  _T_30; // @[Mux.scala 46:19:@2675.4]
  wire [63:0] _T_31; // @[Mux.scala 46:16:@2676.4]
  wire  _T_32; // @[Mux.scala 46:19:@2677.4]
  wire [63:0] _T_33; // @[Mux.scala 46:16:@2678.4]
  wire  _T_34; // @[Mux.scala 46:19:@2679.4]
  wire [63:0] _T_35; // @[Mux.scala 46:16:@2680.4]
  wire  _T_36; // @[Mux.scala 46:19:@2681.4]
  wire [63:0] _T_37; // @[Mux.scala 46:16:@2682.4]
  wire  _T_38; // @[Mux.scala 46:19:@2683.4]
  wire [63:0] _T_39; // @[Mux.scala 46:16:@2684.4]
  wire  _T_40; // @[Mux.scala 46:19:@2685.4]
  wire [63:0] _T_41; // @[Mux.scala 46:16:@2686.4]
  wire  _T_42; // @[Mux.scala 46:19:@2687.4]
  wire [63:0] _T_43; // @[Mux.scala 46:16:@2688.4]
  wire  _T_44; // @[Mux.scala 46:19:@2689.4]
  wire [63:0] res; // @[Mux.scala 46:16:@2690.4]
  wire [63:0] _T_58; // @[execute.scala 43:18:@2696.4]
  wire  nzcv_0; // @[execute.scala 43:25:@2697.4]
  wire  nzcv_1; // @[execute.scala 44:18:@2699.4]
  wire  nzcv_2; // @[execute.scala 46:28:@2702.4]
  wire [63:0] _T_67; // @[execute.scala 48:23:@2705.4]
  wire [63:0] _T_68; // @[execute.scala 48:37:@2706.4]
  wire [64:0] _T_69; // @[execute.scala 48:30:@2707.4]
  wire [63:0] _T_70; // @[execute.scala 48:30:@2708.4]
  wire [63:0] sign_sum; // @[execute.scala 48:30:@2709.4]
  wire  _T_73; // @[execute.scala 49:27:@2711.4]
  wire  _T_76; // @[execute.scala 49:47:@2713.4]
  wire  isPos; // @[execute.scala 49:33:@2714.4]
  wire  _T_79; // @[execute.scala 50:27:@2716.4]
  wire  _T_82; // @[execute.scala 50:47:@2718.4]
  wire  isNeg; // @[execute.scala 50:33:@2719.4]
  wire  _T_84; // @[execute.scala 52:27:@2721.6]
  wire  _T_86; // @[execute.scala 52:16:@2722.6]
  wire  _T_88; // @[execute.scala 54:27:@2727.8]
  wire  _T_90; // @[execute.scala 54:16:@2728.8]
  wire  _GEN_0; // @[execute.scala 53:21:@2726.6]
  wire  nzcv_3; // @[execute.scala 51:15:@2720.4]
  wire [1:0] _T_92; // @[execute.scala 59:19:@2734.4]
  wire [1:0] _T_93; // @[execute.scala 59:19:@2735.4]
  assign _T_16 = io_a & io_b; // @[execute.scala 29:34:@2661.4]
  assign _T_17 = ~ io_b; // @[execute.scala 30:36:@2662.4]
  assign _T_18 = io_a & _T_17; // @[execute.scala 30:34:@2663.4]
  assign _T_19 = io_a | io_b; // @[execute.scala 31:34:@2664.4]
  assign _T_21 = io_a | _T_17; // @[execute.scala 32:34:@2666.4]
  assign _T_22 = io_a ^ io_b; // @[execute.scala 33:34:@2667.4]
  assign _T_24 = io_a ^ _T_17; // @[execute.scala 34:34:@2669.4]
  assign _T_25 = io_a + io_b; // @[execute.scala 35:34:@2670.4]
  assign _T_26 = io_a + io_b; // @[execute.scala 35:34:@2671.4]
  assign _T_27 = io_a - io_b; // @[execute.scala 36:34:@2672.4]
  assign _T_28 = $unsigned(_T_27); // @[execute.scala 36:34:@2673.4]
  assign _T_29 = _T_28[63:0]; // @[execute.scala 36:34:@2674.4]
  assign _T_30 = 3'h7 == io_opcode; // @[Mux.scala 46:19:@2675.4]
  assign _T_31 = _T_30 ? _T_29 : 64'h0; // @[Mux.scala 46:16:@2676.4]
  assign _T_32 = 3'h6 == io_opcode; // @[Mux.scala 46:19:@2677.4]
  assign _T_33 = _T_32 ? _T_26 : _T_31; // @[Mux.scala 46:16:@2678.4]
  assign _T_34 = 3'h5 == io_opcode; // @[Mux.scala 46:19:@2679.4]
  assign _T_35 = _T_34 ? _T_24 : _T_33; // @[Mux.scala 46:16:@2680.4]
  assign _T_36 = 3'h4 == io_opcode; // @[Mux.scala 46:19:@2681.4]
  assign _T_37 = _T_36 ? _T_22 : _T_35; // @[Mux.scala 46:16:@2682.4]
  assign _T_38 = 3'h3 == io_opcode; // @[Mux.scala 46:19:@2683.4]
  assign _T_39 = _T_38 ? _T_21 : _T_37; // @[Mux.scala 46:16:@2684.4]
  assign _T_40 = 3'h2 == io_opcode; // @[Mux.scala 46:19:@2685.4]
  assign _T_41 = _T_40 ? _T_19 : _T_39; // @[Mux.scala 46:16:@2686.4]
  assign _T_42 = 3'h1 == io_opcode; // @[Mux.scala 46:19:@2687.4]
  assign _T_43 = _T_42 ? _T_18 : _T_41; // @[Mux.scala 46:16:@2688.4]
  assign _T_44 = 3'h0 == io_opcode; // @[Mux.scala 46:19:@2689.4]
  assign res = _T_44 ? _T_16 : _T_43; // @[Mux.scala 46:16:@2690.4]
  assign _T_58 = $signed(res); // @[execute.scala 43:18:@2696.4]
  assign nzcv_0 = $signed(_T_58) < $signed(64'sh0); // @[execute.scala 43:25:@2697.4]
  assign nzcv_1 = res == 64'h0; // @[execute.scala 44:18:@2699.4]
  assign nzcv_2 = _T_25[64]; // @[execute.scala 46:28:@2702.4]
  assign _T_67 = $signed(io_a); // @[execute.scala 48:23:@2705.4]
  assign _T_68 = $signed(io_b); // @[execute.scala 48:37:@2706.4]
  assign _T_69 = $signed(_T_67) + $signed(_T_68); // @[execute.scala 48:30:@2707.4]
  assign _T_70 = $signed(_T_67) + $signed(_T_68); // @[execute.scala 48:30:@2708.4]
  assign sign_sum = $signed(_T_70); // @[execute.scala 48:30:@2709.4]
  assign _T_73 = $signed(_T_67) > $signed(64'sh0); // @[execute.scala 49:27:@2711.4]
  assign _T_76 = $signed(_T_68) > $signed(64'sh0); // @[execute.scala 49:47:@2713.4]
  assign isPos = _T_73 & _T_76; // @[execute.scala 49:33:@2714.4]
  assign _T_79 = $signed(_T_67) < $signed(64'sh0); // @[execute.scala 50:27:@2716.4]
  assign _T_82 = $signed(_T_68) < $signed(64'sh0); // @[execute.scala 50:47:@2718.4]
  assign isNeg = _T_79 & _T_82; // @[execute.scala 50:33:@2719.4]
  assign _T_84 = $signed(sign_sum) > $signed(64'sh0); // @[execute.scala 52:27:@2721.6]
  assign _T_86 = _T_84 == 1'h0; // @[execute.scala 52:16:@2722.6]
  assign _T_88 = $signed(sign_sum) < $signed(64'sh0); // @[execute.scala 54:27:@2727.8]
  assign _T_90 = _T_88 == 1'h0; // @[execute.scala 54:16:@2728.8]
  assign _GEN_0 = isNeg ? _T_90 : 1'h0; // @[execute.scala 53:21:@2726.6]
  assign nzcv_3 = isPos ? _T_86 : _GEN_0; // @[execute.scala 51:15:@2720.4]
  assign _T_92 = {nzcv_1,nzcv_0}; // @[execute.scala 59:19:@2734.4]
  assign _T_93 = {nzcv_3,nzcv_2}; // @[execute.scala 59:19:@2735.4]
  assign io_res = _T_44 ? _T_16 : _T_43; // @[execute.scala 61:10:@2738.4]
  assign io_nzcv = {_T_93,_T_92}; // @[execute.scala 59:11:@2737.4]
endmodule
