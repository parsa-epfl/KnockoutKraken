module Move(
  input  [3:0]  io_op,
  input  [1:0]  io_hw,
  input  [15:0] io_imm,
  input  [63:0] io_rd,
  output [63:0] io_res
);
  wire [5:0] pos; // @[Cat.scala 29:58]
  wire  _T_4; // @[Mux.scala 80:60]
  wire [63:0] result; // @[Mux.scala 80:57]
  wire  vecBools_0; // @[Execute.scala 203:33]
  wire  vecBools_1; // @[Execute.scala 203:33]
  wire  vecBools_2; // @[Execute.scala 203:33]
  wire  vecBools_3; // @[Execute.scala 203:33]
  wire  vecBools_4; // @[Execute.scala 203:33]
  wire  vecBools_5; // @[Execute.scala 203:33]
  wire  vecBools_6; // @[Execute.scala 203:33]
  wire  vecBools_7; // @[Execute.scala 203:33]
  wire  vecBools_8; // @[Execute.scala 203:33]
  wire  vecBools_9; // @[Execute.scala 203:33]
  wire  vecBools_10; // @[Execute.scala 203:33]
  wire  vecBools_11; // @[Execute.scala 203:33]
  wire  vecBools_12; // @[Execute.scala 203:33]
  wire  vecBools_13; // @[Execute.scala 203:33]
  wire  vecBools_14; // @[Execute.scala 203:33]
  wire  vecBools_15; // @[Execute.scala 203:33]
  wire  _T_86; // @[Execute.scala 206:14]
  wire  vecResult_0; // @[Execute.scala 206:23]
  wire  _GEN_1; // @[Execute.scala 206:23]
  wire  _GEN_2; // @[Execute.scala 206:23]
  wire  _GEN_3; // @[Execute.scala 206:23]
  wire  _GEN_4; // @[Execute.scala 206:23]
  wire  _GEN_5; // @[Execute.scala 206:23]
  wire  _GEN_6; // @[Execute.scala 206:23]
  wire  _GEN_7; // @[Execute.scala 206:23]
  wire  _GEN_8; // @[Execute.scala 206:23]
  wire  _GEN_9; // @[Execute.scala 206:23]
  wire  _GEN_10; // @[Execute.scala 206:23]
  wire  _GEN_11; // @[Execute.scala 206:23]
  wire  _GEN_12; // @[Execute.scala 206:23]
  wire  _GEN_13; // @[Execute.scala 206:23]
  wire  _GEN_14; // @[Execute.scala 206:23]
  wire  _GEN_15; // @[Execute.scala 206:23]
  wire  _T_87; // @[Execute.scala 206:14]
  wire  vecResult_1; // @[Execute.scala 206:23]
  wire  _GEN_17; // @[Execute.scala 206:23]
  wire  _GEN_18; // @[Execute.scala 206:23]
  wire  _GEN_19; // @[Execute.scala 206:23]
  wire  _GEN_20; // @[Execute.scala 206:23]
  wire  _GEN_21; // @[Execute.scala 206:23]
  wire  _GEN_22; // @[Execute.scala 206:23]
  wire  _GEN_23; // @[Execute.scala 206:23]
  wire  _GEN_24; // @[Execute.scala 206:23]
  wire  _GEN_25; // @[Execute.scala 206:23]
  wire  _GEN_26; // @[Execute.scala 206:23]
  wire  _GEN_27; // @[Execute.scala 206:23]
  wire  _GEN_28; // @[Execute.scala 206:23]
  wire  _GEN_29; // @[Execute.scala 206:23]
  wire  _GEN_30; // @[Execute.scala 206:23]
  wire  _GEN_31; // @[Execute.scala 206:23]
  wire  _T_88; // @[Execute.scala 206:14]
  wire  vecResult_2; // @[Execute.scala 206:23]
  wire  _GEN_33; // @[Execute.scala 206:23]
  wire  _GEN_34; // @[Execute.scala 206:23]
  wire  _GEN_35; // @[Execute.scala 206:23]
  wire  _GEN_36; // @[Execute.scala 206:23]
  wire  _GEN_37; // @[Execute.scala 206:23]
  wire  _GEN_38; // @[Execute.scala 206:23]
  wire  _GEN_39; // @[Execute.scala 206:23]
  wire  _GEN_40; // @[Execute.scala 206:23]
  wire  _GEN_41; // @[Execute.scala 206:23]
  wire  _GEN_42; // @[Execute.scala 206:23]
  wire  _GEN_43; // @[Execute.scala 206:23]
  wire  _GEN_44; // @[Execute.scala 206:23]
  wire  _GEN_45; // @[Execute.scala 206:23]
  wire  _GEN_46; // @[Execute.scala 206:23]
  wire  _GEN_47; // @[Execute.scala 206:23]
  wire  _T_89; // @[Execute.scala 206:14]
  wire  vecResult_3; // @[Execute.scala 206:23]
  wire  _GEN_49; // @[Execute.scala 206:23]
  wire  _GEN_50; // @[Execute.scala 206:23]
  wire  _GEN_51; // @[Execute.scala 206:23]
  wire  _GEN_52; // @[Execute.scala 206:23]
  wire  _GEN_53; // @[Execute.scala 206:23]
  wire  _GEN_54; // @[Execute.scala 206:23]
  wire  _GEN_55; // @[Execute.scala 206:23]
  wire  _GEN_56; // @[Execute.scala 206:23]
  wire  _GEN_57; // @[Execute.scala 206:23]
  wire  _GEN_58; // @[Execute.scala 206:23]
  wire  _GEN_59; // @[Execute.scala 206:23]
  wire  _GEN_60; // @[Execute.scala 206:23]
  wire  _GEN_61; // @[Execute.scala 206:23]
  wire  _GEN_62; // @[Execute.scala 206:23]
  wire  _GEN_63; // @[Execute.scala 206:23]
  wire  _T_90; // @[Execute.scala 206:14]
  wire  vecResult_4; // @[Execute.scala 206:23]
  wire  _GEN_65; // @[Execute.scala 206:23]
  wire  _GEN_66; // @[Execute.scala 206:23]
  wire  _GEN_67; // @[Execute.scala 206:23]
  wire  _GEN_68; // @[Execute.scala 206:23]
  wire  _GEN_69; // @[Execute.scala 206:23]
  wire  _GEN_70; // @[Execute.scala 206:23]
  wire  _GEN_71; // @[Execute.scala 206:23]
  wire  _GEN_72; // @[Execute.scala 206:23]
  wire  _GEN_73; // @[Execute.scala 206:23]
  wire  _GEN_74; // @[Execute.scala 206:23]
  wire  _GEN_75; // @[Execute.scala 206:23]
  wire  _GEN_76; // @[Execute.scala 206:23]
  wire  _GEN_77; // @[Execute.scala 206:23]
  wire  _GEN_78; // @[Execute.scala 206:23]
  wire  _GEN_79; // @[Execute.scala 206:23]
  wire  _T_91; // @[Execute.scala 206:14]
  wire  vecResult_5; // @[Execute.scala 206:23]
  wire  _GEN_81; // @[Execute.scala 206:23]
  wire  _GEN_82; // @[Execute.scala 206:23]
  wire  _GEN_83; // @[Execute.scala 206:23]
  wire  _GEN_84; // @[Execute.scala 206:23]
  wire  _GEN_85; // @[Execute.scala 206:23]
  wire  _GEN_86; // @[Execute.scala 206:23]
  wire  _GEN_87; // @[Execute.scala 206:23]
  wire  _GEN_88; // @[Execute.scala 206:23]
  wire  _GEN_89; // @[Execute.scala 206:23]
  wire  _GEN_90; // @[Execute.scala 206:23]
  wire  _GEN_91; // @[Execute.scala 206:23]
  wire  _GEN_92; // @[Execute.scala 206:23]
  wire  _GEN_93; // @[Execute.scala 206:23]
  wire  _GEN_94; // @[Execute.scala 206:23]
  wire  _GEN_95; // @[Execute.scala 206:23]
  wire  _T_92; // @[Execute.scala 206:14]
  wire  vecResult_6; // @[Execute.scala 206:23]
  wire  _GEN_97; // @[Execute.scala 206:23]
  wire  _GEN_98; // @[Execute.scala 206:23]
  wire  _GEN_99; // @[Execute.scala 206:23]
  wire  _GEN_100; // @[Execute.scala 206:23]
  wire  _GEN_101; // @[Execute.scala 206:23]
  wire  _GEN_102; // @[Execute.scala 206:23]
  wire  _GEN_103; // @[Execute.scala 206:23]
  wire  _GEN_104; // @[Execute.scala 206:23]
  wire  _GEN_105; // @[Execute.scala 206:23]
  wire  _GEN_106; // @[Execute.scala 206:23]
  wire  _GEN_107; // @[Execute.scala 206:23]
  wire  _GEN_108; // @[Execute.scala 206:23]
  wire  _GEN_109; // @[Execute.scala 206:23]
  wire  _GEN_110; // @[Execute.scala 206:23]
  wire  _GEN_111; // @[Execute.scala 206:23]
  wire  _T_93; // @[Execute.scala 206:14]
  wire  vecResult_7; // @[Execute.scala 206:23]
  wire  _GEN_113; // @[Execute.scala 206:23]
  wire  _GEN_114; // @[Execute.scala 206:23]
  wire  _GEN_115; // @[Execute.scala 206:23]
  wire  _GEN_116; // @[Execute.scala 206:23]
  wire  _GEN_117; // @[Execute.scala 206:23]
  wire  _GEN_118; // @[Execute.scala 206:23]
  wire  _GEN_119; // @[Execute.scala 206:23]
  wire  _GEN_120; // @[Execute.scala 206:23]
  wire  _GEN_121; // @[Execute.scala 206:23]
  wire  _GEN_122; // @[Execute.scala 206:23]
  wire  _GEN_123; // @[Execute.scala 206:23]
  wire  _GEN_124; // @[Execute.scala 206:23]
  wire  _GEN_125; // @[Execute.scala 206:23]
  wire  _GEN_126; // @[Execute.scala 206:23]
  wire  _GEN_127; // @[Execute.scala 206:23]
  wire  _T_94; // @[Execute.scala 206:14]
  wire  vecResult_8; // @[Execute.scala 206:23]
  wire  _GEN_129; // @[Execute.scala 206:23]
  wire  _GEN_130; // @[Execute.scala 206:23]
  wire  _GEN_131; // @[Execute.scala 206:23]
  wire  _GEN_132; // @[Execute.scala 206:23]
  wire  _GEN_133; // @[Execute.scala 206:23]
  wire  _GEN_134; // @[Execute.scala 206:23]
  wire  _GEN_135; // @[Execute.scala 206:23]
  wire  _GEN_136; // @[Execute.scala 206:23]
  wire  _GEN_137; // @[Execute.scala 206:23]
  wire  _GEN_138; // @[Execute.scala 206:23]
  wire  _GEN_139; // @[Execute.scala 206:23]
  wire  _GEN_140; // @[Execute.scala 206:23]
  wire  _GEN_141; // @[Execute.scala 206:23]
  wire  _GEN_142; // @[Execute.scala 206:23]
  wire  _GEN_143; // @[Execute.scala 206:23]
  wire  _T_95; // @[Execute.scala 206:14]
  wire  vecResult_9; // @[Execute.scala 206:23]
  wire  _GEN_145; // @[Execute.scala 206:23]
  wire  _GEN_146; // @[Execute.scala 206:23]
  wire  _GEN_147; // @[Execute.scala 206:23]
  wire  _GEN_148; // @[Execute.scala 206:23]
  wire  _GEN_149; // @[Execute.scala 206:23]
  wire  _GEN_150; // @[Execute.scala 206:23]
  wire  _GEN_151; // @[Execute.scala 206:23]
  wire  _GEN_152; // @[Execute.scala 206:23]
  wire  _GEN_153; // @[Execute.scala 206:23]
  wire  _GEN_154; // @[Execute.scala 206:23]
  wire  _GEN_155; // @[Execute.scala 206:23]
  wire  _GEN_156; // @[Execute.scala 206:23]
  wire  _GEN_157; // @[Execute.scala 206:23]
  wire  _GEN_158; // @[Execute.scala 206:23]
  wire  _GEN_159; // @[Execute.scala 206:23]
  wire  _T_96; // @[Execute.scala 206:14]
  wire  vecResult_10; // @[Execute.scala 206:23]
  wire  _GEN_161; // @[Execute.scala 206:23]
  wire  _GEN_162; // @[Execute.scala 206:23]
  wire  _GEN_163; // @[Execute.scala 206:23]
  wire  _GEN_164; // @[Execute.scala 206:23]
  wire  _GEN_165; // @[Execute.scala 206:23]
  wire  _GEN_166; // @[Execute.scala 206:23]
  wire  _GEN_167; // @[Execute.scala 206:23]
  wire  _GEN_168; // @[Execute.scala 206:23]
  wire  _GEN_169; // @[Execute.scala 206:23]
  wire  _GEN_170; // @[Execute.scala 206:23]
  wire  _GEN_171; // @[Execute.scala 206:23]
  wire  _GEN_172; // @[Execute.scala 206:23]
  wire  _GEN_173; // @[Execute.scala 206:23]
  wire  _GEN_174; // @[Execute.scala 206:23]
  wire  _GEN_175; // @[Execute.scala 206:23]
  wire  _T_97; // @[Execute.scala 206:14]
  wire  vecResult_11; // @[Execute.scala 206:23]
  wire  _GEN_177; // @[Execute.scala 206:23]
  wire  _GEN_178; // @[Execute.scala 206:23]
  wire  _GEN_179; // @[Execute.scala 206:23]
  wire  _GEN_180; // @[Execute.scala 206:23]
  wire  _GEN_181; // @[Execute.scala 206:23]
  wire  _GEN_182; // @[Execute.scala 206:23]
  wire  _GEN_183; // @[Execute.scala 206:23]
  wire  _GEN_184; // @[Execute.scala 206:23]
  wire  _GEN_185; // @[Execute.scala 206:23]
  wire  _GEN_186; // @[Execute.scala 206:23]
  wire  _GEN_187; // @[Execute.scala 206:23]
  wire  _GEN_188; // @[Execute.scala 206:23]
  wire  _GEN_189; // @[Execute.scala 206:23]
  wire  _GEN_190; // @[Execute.scala 206:23]
  wire  _GEN_191; // @[Execute.scala 206:23]
  wire  _T_98; // @[Execute.scala 206:14]
  wire  vecResult_12; // @[Execute.scala 206:23]
  wire  _GEN_193; // @[Execute.scala 206:23]
  wire  _GEN_194; // @[Execute.scala 206:23]
  wire  _GEN_195; // @[Execute.scala 206:23]
  wire  _GEN_196; // @[Execute.scala 206:23]
  wire  _GEN_197; // @[Execute.scala 206:23]
  wire  _GEN_198; // @[Execute.scala 206:23]
  wire  _GEN_199; // @[Execute.scala 206:23]
  wire  _GEN_200; // @[Execute.scala 206:23]
  wire  _GEN_201; // @[Execute.scala 206:23]
  wire  _GEN_202; // @[Execute.scala 206:23]
  wire  _GEN_203; // @[Execute.scala 206:23]
  wire  _GEN_204; // @[Execute.scala 206:23]
  wire  _GEN_205; // @[Execute.scala 206:23]
  wire  _GEN_206; // @[Execute.scala 206:23]
  wire  _GEN_207; // @[Execute.scala 206:23]
  wire  _T_99; // @[Execute.scala 206:14]
  wire  vecResult_13; // @[Execute.scala 206:23]
  wire  _GEN_209; // @[Execute.scala 206:23]
  wire  _GEN_210; // @[Execute.scala 206:23]
  wire  _GEN_211; // @[Execute.scala 206:23]
  wire  _GEN_212; // @[Execute.scala 206:23]
  wire  _GEN_213; // @[Execute.scala 206:23]
  wire  _GEN_214; // @[Execute.scala 206:23]
  wire  _GEN_215; // @[Execute.scala 206:23]
  wire  _GEN_216; // @[Execute.scala 206:23]
  wire  _GEN_217; // @[Execute.scala 206:23]
  wire  _GEN_218; // @[Execute.scala 206:23]
  wire  _GEN_219; // @[Execute.scala 206:23]
  wire  _GEN_220; // @[Execute.scala 206:23]
  wire  _GEN_221; // @[Execute.scala 206:23]
  wire  _GEN_222; // @[Execute.scala 206:23]
  wire  _GEN_223; // @[Execute.scala 206:23]
  wire  _T_100; // @[Execute.scala 206:14]
  wire  vecResult_14; // @[Execute.scala 206:23]
  wire  _GEN_225; // @[Execute.scala 206:23]
  wire  _GEN_226; // @[Execute.scala 206:23]
  wire  _GEN_227; // @[Execute.scala 206:23]
  wire  _GEN_228; // @[Execute.scala 206:23]
  wire  _GEN_229; // @[Execute.scala 206:23]
  wire  _GEN_230; // @[Execute.scala 206:23]
  wire  _GEN_231; // @[Execute.scala 206:23]
  wire  _GEN_232; // @[Execute.scala 206:23]
  wire  _GEN_233; // @[Execute.scala 206:23]
  wire  _GEN_234; // @[Execute.scala 206:23]
  wire  _GEN_235; // @[Execute.scala 206:23]
  wire  _GEN_236; // @[Execute.scala 206:23]
  wire  _GEN_237; // @[Execute.scala 206:23]
  wire  _GEN_238; // @[Execute.scala 206:23]
  wire  _GEN_239; // @[Execute.scala 206:23]
  wire  _T_101; // @[Execute.scala 206:14]
  wire  vecResult_15; // @[Execute.scala 206:23]
  wire  _GEN_241; // @[Execute.scala 206:23]
  wire  _GEN_242; // @[Execute.scala 206:23]
  wire  _GEN_243; // @[Execute.scala 206:23]
  wire  _GEN_244; // @[Execute.scala 206:23]
  wire  _GEN_245; // @[Execute.scala 206:23]
  wire  _GEN_246; // @[Execute.scala 206:23]
  wire  _GEN_247; // @[Execute.scala 206:23]
  wire  _GEN_248; // @[Execute.scala 206:23]
  wire  _GEN_249; // @[Execute.scala 206:23]
  wire  _GEN_250; // @[Execute.scala 206:23]
  wire  _GEN_251; // @[Execute.scala 206:23]
  wire  _GEN_252; // @[Execute.scala 206:23]
  wire  _GEN_253; // @[Execute.scala 206:23]
  wire  _GEN_254; // @[Execute.scala 206:23]
  wire  _GEN_255; // @[Execute.scala 206:23]
  wire  _T_102; // @[Execute.scala 206:14]
  wire  vecResult_16; // @[Execute.scala 206:23]
  wire  _GEN_257; // @[Execute.scala 206:23]
  wire  _GEN_258; // @[Execute.scala 206:23]
  wire  _GEN_259; // @[Execute.scala 206:23]
  wire  _GEN_260; // @[Execute.scala 206:23]
  wire  _GEN_261; // @[Execute.scala 206:23]
  wire  _GEN_262; // @[Execute.scala 206:23]
  wire  _GEN_263; // @[Execute.scala 206:23]
  wire  _GEN_264; // @[Execute.scala 206:23]
  wire  _GEN_265; // @[Execute.scala 206:23]
  wire  _GEN_266; // @[Execute.scala 206:23]
  wire  _GEN_267; // @[Execute.scala 206:23]
  wire  _GEN_268; // @[Execute.scala 206:23]
  wire  _GEN_269; // @[Execute.scala 206:23]
  wire  _GEN_270; // @[Execute.scala 206:23]
  wire  _GEN_271; // @[Execute.scala 206:23]
  wire  _T_103; // @[Execute.scala 206:14]
  wire  vecResult_17; // @[Execute.scala 206:23]
  wire  _GEN_273; // @[Execute.scala 206:23]
  wire  _GEN_274; // @[Execute.scala 206:23]
  wire  _GEN_275; // @[Execute.scala 206:23]
  wire  _GEN_276; // @[Execute.scala 206:23]
  wire  _GEN_277; // @[Execute.scala 206:23]
  wire  _GEN_278; // @[Execute.scala 206:23]
  wire  _GEN_279; // @[Execute.scala 206:23]
  wire  _GEN_280; // @[Execute.scala 206:23]
  wire  _GEN_281; // @[Execute.scala 206:23]
  wire  _GEN_282; // @[Execute.scala 206:23]
  wire  _GEN_283; // @[Execute.scala 206:23]
  wire  _GEN_284; // @[Execute.scala 206:23]
  wire  _GEN_285; // @[Execute.scala 206:23]
  wire  _GEN_286; // @[Execute.scala 206:23]
  wire  _GEN_287; // @[Execute.scala 206:23]
  wire  _T_104; // @[Execute.scala 206:14]
  wire  vecResult_18; // @[Execute.scala 206:23]
  wire  _GEN_289; // @[Execute.scala 206:23]
  wire  _GEN_290; // @[Execute.scala 206:23]
  wire  _GEN_291; // @[Execute.scala 206:23]
  wire  _GEN_292; // @[Execute.scala 206:23]
  wire  _GEN_293; // @[Execute.scala 206:23]
  wire  _GEN_294; // @[Execute.scala 206:23]
  wire  _GEN_295; // @[Execute.scala 206:23]
  wire  _GEN_296; // @[Execute.scala 206:23]
  wire  _GEN_297; // @[Execute.scala 206:23]
  wire  _GEN_298; // @[Execute.scala 206:23]
  wire  _GEN_299; // @[Execute.scala 206:23]
  wire  _GEN_300; // @[Execute.scala 206:23]
  wire  _GEN_301; // @[Execute.scala 206:23]
  wire  _GEN_302; // @[Execute.scala 206:23]
  wire  _GEN_303; // @[Execute.scala 206:23]
  wire  _T_105; // @[Execute.scala 206:14]
  wire  vecResult_19; // @[Execute.scala 206:23]
  wire  _GEN_305; // @[Execute.scala 206:23]
  wire  _GEN_306; // @[Execute.scala 206:23]
  wire  _GEN_307; // @[Execute.scala 206:23]
  wire  _GEN_308; // @[Execute.scala 206:23]
  wire  _GEN_309; // @[Execute.scala 206:23]
  wire  _GEN_310; // @[Execute.scala 206:23]
  wire  _GEN_311; // @[Execute.scala 206:23]
  wire  _GEN_312; // @[Execute.scala 206:23]
  wire  _GEN_313; // @[Execute.scala 206:23]
  wire  _GEN_314; // @[Execute.scala 206:23]
  wire  _GEN_315; // @[Execute.scala 206:23]
  wire  _GEN_316; // @[Execute.scala 206:23]
  wire  _GEN_317; // @[Execute.scala 206:23]
  wire  _GEN_318; // @[Execute.scala 206:23]
  wire  _GEN_319; // @[Execute.scala 206:23]
  wire  _T_106; // @[Execute.scala 206:14]
  wire  vecResult_20; // @[Execute.scala 206:23]
  wire  _GEN_321; // @[Execute.scala 206:23]
  wire  _GEN_322; // @[Execute.scala 206:23]
  wire  _GEN_323; // @[Execute.scala 206:23]
  wire  _GEN_324; // @[Execute.scala 206:23]
  wire  _GEN_325; // @[Execute.scala 206:23]
  wire  _GEN_326; // @[Execute.scala 206:23]
  wire  _GEN_327; // @[Execute.scala 206:23]
  wire  _GEN_328; // @[Execute.scala 206:23]
  wire  _GEN_329; // @[Execute.scala 206:23]
  wire  _GEN_330; // @[Execute.scala 206:23]
  wire  _GEN_331; // @[Execute.scala 206:23]
  wire  _GEN_332; // @[Execute.scala 206:23]
  wire  _GEN_333; // @[Execute.scala 206:23]
  wire  _GEN_334; // @[Execute.scala 206:23]
  wire  _GEN_335; // @[Execute.scala 206:23]
  wire  _T_107; // @[Execute.scala 206:14]
  wire  vecResult_21; // @[Execute.scala 206:23]
  wire  _GEN_337; // @[Execute.scala 206:23]
  wire  _GEN_338; // @[Execute.scala 206:23]
  wire  _GEN_339; // @[Execute.scala 206:23]
  wire  _GEN_340; // @[Execute.scala 206:23]
  wire  _GEN_341; // @[Execute.scala 206:23]
  wire  _GEN_342; // @[Execute.scala 206:23]
  wire  _GEN_343; // @[Execute.scala 206:23]
  wire  _GEN_344; // @[Execute.scala 206:23]
  wire  _GEN_345; // @[Execute.scala 206:23]
  wire  _GEN_346; // @[Execute.scala 206:23]
  wire  _GEN_347; // @[Execute.scala 206:23]
  wire  _GEN_348; // @[Execute.scala 206:23]
  wire  _GEN_349; // @[Execute.scala 206:23]
  wire  _GEN_350; // @[Execute.scala 206:23]
  wire  _GEN_351; // @[Execute.scala 206:23]
  wire  _T_108; // @[Execute.scala 206:14]
  wire  vecResult_22; // @[Execute.scala 206:23]
  wire  _GEN_353; // @[Execute.scala 206:23]
  wire  _GEN_354; // @[Execute.scala 206:23]
  wire  _GEN_355; // @[Execute.scala 206:23]
  wire  _GEN_356; // @[Execute.scala 206:23]
  wire  _GEN_357; // @[Execute.scala 206:23]
  wire  _GEN_358; // @[Execute.scala 206:23]
  wire  _GEN_359; // @[Execute.scala 206:23]
  wire  _GEN_360; // @[Execute.scala 206:23]
  wire  _GEN_361; // @[Execute.scala 206:23]
  wire  _GEN_362; // @[Execute.scala 206:23]
  wire  _GEN_363; // @[Execute.scala 206:23]
  wire  _GEN_364; // @[Execute.scala 206:23]
  wire  _GEN_365; // @[Execute.scala 206:23]
  wire  _GEN_366; // @[Execute.scala 206:23]
  wire  _GEN_367; // @[Execute.scala 206:23]
  wire  _T_109; // @[Execute.scala 206:14]
  wire  vecResult_23; // @[Execute.scala 206:23]
  wire  _GEN_369; // @[Execute.scala 206:23]
  wire  _GEN_370; // @[Execute.scala 206:23]
  wire  _GEN_371; // @[Execute.scala 206:23]
  wire  _GEN_372; // @[Execute.scala 206:23]
  wire  _GEN_373; // @[Execute.scala 206:23]
  wire  _GEN_374; // @[Execute.scala 206:23]
  wire  _GEN_375; // @[Execute.scala 206:23]
  wire  _GEN_376; // @[Execute.scala 206:23]
  wire  _GEN_377; // @[Execute.scala 206:23]
  wire  _GEN_378; // @[Execute.scala 206:23]
  wire  _GEN_379; // @[Execute.scala 206:23]
  wire  _GEN_380; // @[Execute.scala 206:23]
  wire  _GEN_381; // @[Execute.scala 206:23]
  wire  _GEN_382; // @[Execute.scala 206:23]
  wire  _GEN_383; // @[Execute.scala 206:23]
  wire  _T_110; // @[Execute.scala 206:14]
  wire  vecResult_24; // @[Execute.scala 206:23]
  wire  _GEN_385; // @[Execute.scala 206:23]
  wire  _GEN_386; // @[Execute.scala 206:23]
  wire  _GEN_387; // @[Execute.scala 206:23]
  wire  _GEN_388; // @[Execute.scala 206:23]
  wire  _GEN_389; // @[Execute.scala 206:23]
  wire  _GEN_390; // @[Execute.scala 206:23]
  wire  _GEN_391; // @[Execute.scala 206:23]
  wire  _GEN_392; // @[Execute.scala 206:23]
  wire  _GEN_393; // @[Execute.scala 206:23]
  wire  _GEN_394; // @[Execute.scala 206:23]
  wire  _GEN_395; // @[Execute.scala 206:23]
  wire  _GEN_396; // @[Execute.scala 206:23]
  wire  _GEN_397; // @[Execute.scala 206:23]
  wire  _GEN_398; // @[Execute.scala 206:23]
  wire  _GEN_399; // @[Execute.scala 206:23]
  wire  _T_111; // @[Execute.scala 206:14]
  wire  vecResult_25; // @[Execute.scala 206:23]
  wire  _GEN_401; // @[Execute.scala 206:23]
  wire  _GEN_402; // @[Execute.scala 206:23]
  wire  _GEN_403; // @[Execute.scala 206:23]
  wire  _GEN_404; // @[Execute.scala 206:23]
  wire  _GEN_405; // @[Execute.scala 206:23]
  wire  _GEN_406; // @[Execute.scala 206:23]
  wire  _GEN_407; // @[Execute.scala 206:23]
  wire  _GEN_408; // @[Execute.scala 206:23]
  wire  _GEN_409; // @[Execute.scala 206:23]
  wire  _GEN_410; // @[Execute.scala 206:23]
  wire  _GEN_411; // @[Execute.scala 206:23]
  wire  _GEN_412; // @[Execute.scala 206:23]
  wire  _GEN_413; // @[Execute.scala 206:23]
  wire  _GEN_414; // @[Execute.scala 206:23]
  wire  _GEN_415; // @[Execute.scala 206:23]
  wire  _T_112; // @[Execute.scala 206:14]
  wire  vecResult_26; // @[Execute.scala 206:23]
  wire  _GEN_417; // @[Execute.scala 206:23]
  wire  _GEN_418; // @[Execute.scala 206:23]
  wire  _GEN_419; // @[Execute.scala 206:23]
  wire  _GEN_420; // @[Execute.scala 206:23]
  wire  _GEN_421; // @[Execute.scala 206:23]
  wire  _GEN_422; // @[Execute.scala 206:23]
  wire  _GEN_423; // @[Execute.scala 206:23]
  wire  _GEN_424; // @[Execute.scala 206:23]
  wire  _GEN_425; // @[Execute.scala 206:23]
  wire  _GEN_426; // @[Execute.scala 206:23]
  wire  _GEN_427; // @[Execute.scala 206:23]
  wire  _GEN_428; // @[Execute.scala 206:23]
  wire  _GEN_429; // @[Execute.scala 206:23]
  wire  _GEN_430; // @[Execute.scala 206:23]
  wire  _GEN_431; // @[Execute.scala 206:23]
  wire  _T_113; // @[Execute.scala 206:14]
  wire  vecResult_27; // @[Execute.scala 206:23]
  wire  _GEN_433; // @[Execute.scala 206:23]
  wire  _GEN_434; // @[Execute.scala 206:23]
  wire  _GEN_435; // @[Execute.scala 206:23]
  wire  _GEN_436; // @[Execute.scala 206:23]
  wire  _GEN_437; // @[Execute.scala 206:23]
  wire  _GEN_438; // @[Execute.scala 206:23]
  wire  _GEN_439; // @[Execute.scala 206:23]
  wire  _GEN_440; // @[Execute.scala 206:23]
  wire  _GEN_441; // @[Execute.scala 206:23]
  wire  _GEN_442; // @[Execute.scala 206:23]
  wire  _GEN_443; // @[Execute.scala 206:23]
  wire  _GEN_444; // @[Execute.scala 206:23]
  wire  _GEN_445; // @[Execute.scala 206:23]
  wire  _GEN_446; // @[Execute.scala 206:23]
  wire  _GEN_447; // @[Execute.scala 206:23]
  wire  _T_114; // @[Execute.scala 206:14]
  wire  vecResult_28; // @[Execute.scala 206:23]
  wire  _GEN_449; // @[Execute.scala 206:23]
  wire  _GEN_450; // @[Execute.scala 206:23]
  wire  _GEN_451; // @[Execute.scala 206:23]
  wire  _GEN_452; // @[Execute.scala 206:23]
  wire  _GEN_453; // @[Execute.scala 206:23]
  wire  _GEN_454; // @[Execute.scala 206:23]
  wire  _GEN_455; // @[Execute.scala 206:23]
  wire  _GEN_456; // @[Execute.scala 206:23]
  wire  _GEN_457; // @[Execute.scala 206:23]
  wire  _GEN_458; // @[Execute.scala 206:23]
  wire  _GEN_459; // @[Execute.scala 206:23]
  wire  _GEN_460; // @[Execute.scala 206:23]
  wire  _GEN_461; // @[Execute.scala 206:23]
  wire  _GEN_462; // @[Execute.scala 206:23]
  wire  _GEN_463; // @[Execute.scala 206:23]
  wire  _T_115; // @[Execute.scala 206:14]
  wire  vecResult_29; // @[Execute.scala 206:23]
  wire  _GEN_465; // @[Execute.scala 206:23]
  wire  _GEN_466; // @[Execute.scala 206:23]
  wire  _GEN_467; // @[Execute.scala 206:23]
  wire  _GEN_468; // @[Execute.scala 206:23]
  wire  _GEN_469; // @[Execute.scala 206:23]
  wire  _GEN_470; // @[Execute.scala 206:23]
  wire  _GEN_471; // @[Execute.scala 206:23]
  wire  _GEN_472; // @[Execute.scala 206:23]
  wire  _GEN_473; // @[Execute.scala 206:23]
  wire  _GEN_474; // @[Execute.scala 206:23]
  wire  _GEN_475; // @[Execute.scala 206:23]
  wire  _GEN_476; // @[Execute.scala 206:23]
  wire  _GEN_477; // @[Execute.scala 206:23]
  wire  _GEN_478; // @[Execute.scala 206:23]
  wire  _GEN_479; // @[Execute.scala 206:23]
  wire  _T_116; // @[Execute.scala 206:14]
  wire  vecResult_30; // @[Execute.scala 206:23]
  wire  _GEN_481; // @[Execute.scala 206:23]
  wire  _GEN_482; // @[Execute.scala 206:23]
  wire  _GEN_483; // @[Execute.scala 206:23]
  wire  _GEN_484; // @[Execute.scala 206:23]
  wire  _GEN_485; // @[Execute.scala 206:23]
  wire  _GEN_486; // @[Execute.scala 206:23]
  wire  _GEN_487; // @[Execute.scala 206:23]
  wire  _GEN_488; // @[Execute.scala 206:23]
  wire  _GEN_489; // @[Execute.scala 206:23]
  wire  _GEN_490; // @[Execute.scala 206:23]
  wire  _GEN_491; // @[Execute.scala 206:23]
  wire  _GEN_492; // @[Execute.scala 206:23]
  wire  _GEN_493; // @[Execute.scala 206:23]
  wire  _GEN_494; // @[Execute.scala 206:23]
  wire  _GEN_495; // @[Execute.scala 206:23]
  wire  _T_117; // @[Execute.scala 206:14]
  wire  vecResult_31; // @[Execute.scala 206:23]
  wire  _GEN_497; // @[Execute.scala 206:23]
  wire  _GEN_498; // @[Execute.scala 206:23]
  wire  _GEN_499; // @[Execute.scala 206:23]
  wire  _GEN_500; // @[Execute.scala 206:23]
  wire  _GEN_501; // @[Execute.scala 206:23]
  wire  _GEN_502; // @[Execute.scala 206:23]
  wire  _GEN_503; // @[Execute.scala 206:23]
  wire  _GEN_504; // @[Execute.scala 206:23]
  wire  _GEN_505; // @[Execute.scala 206:23]
  wire  _GEN_506; // @[Execute.scala 206:23]
  wire  _GEN_507; // @[Execute.scala 206:23]
  wire  _GEN_508; // @[Execute.scala 206:23]
  wire  _GEN_509; // @[Execute.scala 206:23]
  wire  _GEN_510; // @[Execute.scala 206:23]
  wire  _GEN_511; // @[Execute.scala 206:23]
  wire  _T_118; // @[Execute.scala 206:14]
  wire  vecResult_32; // @[Execute.scala 206:23]
  wire  _GEN_513; // @[Execute.scala 206:23]
  wire  _GEN_514; // @[Execute.scala 206:23]
  wire  _GEN_515; // @[Execute.scala 206:23]
  wire  _GEN_516; // @[Execute.scala 206:23]
  wire  _GEN_517; // @[Execute.scala 206:23]
  wire  _GEN_518; // @[Execute.scala 206:23]
  wire  _GEN_519; // @[Execute.scala 206:23]
  wire  _GEN_520; // @[Execute.scala 206:23]
  wire  _GEN_521; // @[Execute.scala 206:23]
  wire  _GEN_522; // @[Execute.scala 206:23]
  wire  _GEN_523; // @[Execute.scala 206:23]
  wire  _GEN_524; // @[Execute.scala 206:23]
  wire  _GEN_525; // @[Execute.scala 206:23]
  wire  _GEN_526; // @[Execute.scala 206:23]
  wire  _GEN_527; // @[Execute.scala 206:23]
  wire  _T_119; // @[Execute.scala 206:14]
  wire  vecResult_33; // @[Execute.scala 206:23]
  wire  _GEN_529; // @[Execute.scala 206:23]
  wire  _GEN_530; // @[Execute.scala 206:23]
  wire  _GEN_531; // @[Execute.scala 206:23]
  wire  _GEN_532; // @[Execute.scala 206:23]
  wire  _GEN_533; // @[Execute.scala 206:23]
  wire  _GEN_534; // @[Execute.scala 206:23]
  wire  _GEN_535; // @[Execute.scala 206:23]
  wire  _GEN_536; // @[Execute.scala 206:23]
  wire  _GEN_537; // @[Execute.scala 206:23]
  wire  _GEN_538; // @[Execute.scala 206:23]
  wire  _GEN_539; // @[Execute.scala 206:23]
  wire  _GEN_540; // @[Execute.scala 206:23]
  wire  _GEN_541; // @[Execute.scala 206:23]
  wire  _GEN_542; // @[Execute.scala 206:23]
  wire  _GEN_543; // @[Execute.scala 206:23]
  wire  _T_120; // @[Execute.scala 206:14]
  wire  vecResult_34; // @[Execute.scala 206:23]
  wire  _GEN_545; // @[Execute.scala 206:23]
  wire  _GEN_546; // @[Execute.scala 206:23]
  wire  _GEN_547; // @[Execute.scala 206:23]
  wire  _GEN_548; // @[Execute.scala 206:23]
  wire  _GEN_549; // @[Execute.scala 206:23]
  wire  _GEN_550; // @[Execute.scala 206:23]
  wire  _GEN_551; // @[Execute.scala 206:23]
  wire  _GEN_552; // @[Execute.scala 206:23]
  wire  _GEN_553; // @[Execute.scala 206:23]
  wire  _GEN_554; // @[Execute.scala 206:23]
  wire  _GEN_555; // @[Execute.scala 206:23]
  wire  _GEN_556; // @[Execute.scala 206:23]
  wire  _GEN_557; // @[Execute.scala 206:23]
  wire  _GEN_558; // @[Execute.scala 206:23]
  wire  _GEN_559; // @[Execute.scala 206:23]
  wire  _T_121; // @[Execute.scala 206:14]
  wire  vecResult_35; // @[Execute.scala 206:23]
  wire  _GEN_561; // @[Execute.scala 206:23]
  wire  _GEN_562; // @[Execute.scala 206:23]
  wire  _GEN_563; // @[Execute.scala 206:23]
  wire  _GEN_564; // @[Execute.scala 206:23]
  wire  _GEN_565; // @[Execute.scala 206:23]
  wire  _GEN_566; // @[Execute.scala 206:23]
  wire  _GEN_567; // @[Execute.scala 206:23]
  wire  _GEN_568; // @[Execute.scala 206:23]
  wire  _GEN_569; // @[Execute.scala 206:23]
  wire  _GEN_570; // @[Execute.scala 206:23]
  wire  _GEN_571; // @[Execute.scala 206:23]
  wire  _GEN_572; // @[Execute.scala 206:23]
  wire  _GEN_573; // @[Execute.scala 206:23]
  wire  _GEN_574; // @[Execute.scala 206:23]
  wire  _GEN_575; // @[Execute.scala 206:23]
  wire  _T_122; // @[Execute.scala 206:14]
  wire  vecResult_36; // @[Execute.scala 206:23]
  wire  _GEN_577; // @[Execute.scala 206:23]
  wire  _GEN_578; // @[Execute.scala 206:23]
  wire  _GEN_579; // @[Execute.scala 206:23]
  wire  _GEN_580; // @[Execute.scala 206:23]
  wire  _GEN_581; // @[Execute.scala 206:23]
  wire  _GEN_582; // @[Execute.scala 206:23]
  wire  _GEN_583; // @[Execute.scala 206:23]
  wire  _GEN_584; // @[Execute.scala 206:23]
  wire  _GEN_585; // @[Execute.scala 206:23]
  wire  _GEN_586; // @[Execute.scala 206:23]
  wire  _GEN_587; // @[Execute.scala 206:23]
  wire  _GEN_588; // @[Execute.scala 206:23]
  wire  _GEN_589; // @[Execute.scala 206:23]
  wire  _GEN_590; // @[Execute.scala 206:23]
  wire  _GEN_591; // @[Execute.scala 206:23]
  wire  _T_123; // @[Execute.scala 206:14]
  wire  vecResult_37; // @[Execute.scala 206:23]
  wire  _GEN_593; // @[Execute.scala 206:23]
  wire  _GEN_594; // @[Execute.scala 206:23]
  wire  _GEN_595; // @[Execute.scala 206:23]
  wire  _GEN_596; // @[Execute.scala 206:23]
  wire  _GEN_597; // @[Execute.scala 206:23]
  wire  _GEN_598; // @[Execute.scala 206:23]
  wire  _GEN_599; // @[Execute.scala 206:23]
  wire  _GEN_600; // @[Execute.scala 206:23]
  wire  _GEN_601; // @[Execute.scala 206:23]
  wire  _GEN_602; // @[Execute.scala 206:23]
  wire  _GEN_603; // @[Execute.scala 206:23]
  wire  _GEN_604; // @[Execute.scala 206:23]
  wire  _GEN_605; // @[Execute.scala 206:23]
  wire  _GEN_606; // @[Execute.scala 206:23]
  wire  _GEN_607; // @[Execute.scala 206:23]
  wire  _T_124; // @[Execute.scala 206:14]
  wire  vecResult_38; // @[Execute.scala 206:23]
  wire  _GEN_609; // @[Execute.scala 206:23]
  wire  _GEN_610; // @[Execute.scala 206:23]
  wire  _GEN_611; // @[Execute.scala 206:23]
  wire  _GEN_612; // @[Execute.scala 206:23]
  wire  _GEN_613; // @[Execute.scala 206:23]
  wire  _GEN_614; // @[Execute.scala 206:23]
  wire  _GEN_615; // @[Execute.scala 206:23]
  wire  _GEN_616; // @[Execute.scala 206:23]
  wire  _GEN_617; // @[Execute.scala 206:23]
  wire  _GEN_618; // @[Execute.scala 206:23]
  wire  _GEN_619; // @[Execute.scala 206:23]
  wire  _GEN_620; // @[Execute.scala 206:23]
  wire  _GEN_621; // @[Execute.scala 206:23]
  wire  _GEN_622; // @[Execute.scala 206:23]
  wire  _GEN_623; // @[Execute.scala 206:23]
  wire  _T_125; // @[Execute.scala 206:14]
  wire  vecResult_39; // @[Execute.scala 206:23]
  wire  _GEN_625; // @[Execute.scala 206:23]
  wire  _GEN_626; // @[Execute.scala 206:23]
  wire  _GEN_627; // @[Execute.scala 206:23]
  wire  _GEN_628; // @[Execute.scala 206:23]
  wire  _GEN_629; // @[Execute.scala 206:23]
  wire  _GEN_630; // @[Execute.scala 206:23]
  wire  _GEN_631; // @[Execute.scala 206:23]
  wire  _GEN_632; // @[Execute.scala 206:23]
  wire  _GEN_633; // @[Execute.scala 206:23]
  wire  _GEN_634; // @[Execute.scala 206:23]
  wire  _GEN_635; // @[Execute.scala 206:23]
  wire  _GEN_636; // @[Execute.scala 206:23]
  wire  _GEN_637; // @[Execute.scala 206:23]
  wire  _GEN_638; // @[Execute.scala 206:23]
  wire  _GEN_639; // @[Execute.scala 206:23]
  wire  _T_126; // @[Execute.scala 206:14]
  wire  vecResult_40; // @[Execute.scala 206:23]
  wire  _GEN_641; // @[Execute.scala 206:23]
  wire  _GEN_642; // @[Execute.scala 206:23]
  wire  _GEN_643; // @[Execute.scala 206:23]
  wire  _GEN_644; // @[Execute.scala 206:23]
  wire  _GEN_645; // @[Execute.scala 206:23]
  wire  _GEN_646; // @[Execute.scala 206:23]
  wire  _GEN_647; // @[Execute.scala 206:23]
  wire  _GEN_648; // @[Execute.scala 206:23]
  wire  _GEN_649; // @[Execute.scala 206:23]
  wire  _GEN_650; // @[Execute.scala 206:23]
  wire  _GEN_651; // @[Execute.scala 206:23]
  wire  _GEN_652; // @[Execute.scala 206:23]
  wire  _GEN_653; // @[Execute.scala 206:23]
  wire  _GEN_654; // @[Execute.scala 206:23]
  wire  _GEN_655; // @[Execute.scala 206:23]
  wire  _T_127; // @[Execute.scala 206:14]
  wire  vecResult_41; // @[Execute.scala 206:23]
  wire  _GEN_657; // @[Execute.scala 206:23]
  wire  _GEN_658; // @[Execute.scala 206:23]
  wire  _GEN_659; // @[Execute.scala 206:23]
  wire  _GEN_660; // @[Execute.scala 206:23]
  wire  _GEN_661; // @[Execute.scala 206:23]
  wire  _GEN_662; // @[Execute.scala 206:23]
  wire  _GEN_663; // @[Execute.scala 206:23]
  wire  _GEN_664; // @[Execute.scala 206:23]
  wire  _GEN_665; // @[Execute.scala 206:23]
  wire  _GEN_666; // @[Execute.scala 206:23]
  wire  _GEN_667; // @[Execute.scala 206:23]
  wire  _GEN_668; // @[Execute.scala 206:23]
  wire  _GEN_669; // @[Execute.scala 206:23]
  wire  _GEN_670; // @[Execute.scala 206:23]
  wire  _GEN_671; // @[Execute.scala 206:23]
  wire  _T_128; // @[Execute.scala 206:14]
  wire  vecResult_42; // @[Execute.scala 206:23]
  wire  _GEN_673; // @[Execute.scala 206:23]
  wire  _GEN_674; // @[Execute.scala 206:23]
  wire  _GEN_675; // @[Execute.scala 206:23]
  wire  _GEN_676; // @[Execute.scala 206:23]
  wire  _GEN_677; // @[Execute.scala 206:23]
  wire  _GEN_678; // @[Execute.scala 206:23]
  wire  _GEN_679; // @[Execute.scala 206:23]
  wire  _GEN_680; // @[Execute.scala 206:23]
  wire  _GEN_681; // @[Execute.scala 206:23]
  wire  _GEN_682; // @[Execute.scala 206:23]
  wire  _GEN_683; // @[Execute.scala 206:23]
  wire  _GEN_684; // @[Execute.scala 206:23]
  wire  _GEN_685; // @[Execute.scala 206:23]
  wire  _GEN_686; // @[Execute.scala 206:23]
  wire  _GEN_687; // @[Execute.scala 206:23]
  wire  _T_129; // @[Execute.scala 206:14]
  wire  vecResult_43; // @[Execute.scala 206:23]
  wire  _GEN_689; // @[Execute.scala 206:23]
  wire  _GEN_690; // @[Execute.scala 206:23]
  wire  _GEN_691; // @[Execute.scala 206:23]
  wire  _GEN_692; // @[Execute.scala 206:23]
  wire  _GEN_693; // @[Execute.scala 206:23]
  wire  _GEN_694; // @[Execute.scala 206:23]
  wire  _GEN_695; // @[Execute.scala 206:23]
  wire  _GEN_696; // @[Execute.scala 206:23]
  wire  _GEN_697; // @[Execute.scala 206:23]
  wire  _GEN_698; // @[Execute.scala 206:23]
  wire  _GEN_699; // @[Execute.scala 206:23]
  wire  _GEN_700; // @[Execute.scala 206:23]
  wire  _GEN_701; // @[Execute.scala 206:23]
  wire  _GEN_702; // @[Execute.scala 206:23]
  wire  _GEN_703; // @[Execute.scala 206:23]
  wire  _T_130; // @[Execute.scala 206:14]
  wire  vecResult_44; // @[Execute.scala 206:23]
  wire  _GEN_705; // @[Execute.scala 206:23]
  wire  _GEN_706; // @[Execute.scala 206:23]
  wire  _GEN_707; // @[Execute.scala 206:23]
  wire  _GEN_708; // @[Execute.scala 206:23]
  wire  _GEN_709; // @[Execute.scala 206:23]
  wire  _GEN_710; // @[Execute.scala 206:23]
  wire  _GEN_711; // @[Execute.scala 206:23]
  wire  _GEN_712; // @[Execute.scala 206:23]
  wire  _GEN_713; // @[Execute.scala 206:23]
  wire  _GEN_714; // @[Execute.scala 206:23]
  wire  _GEN_715; // @[Execute.scala 206:23]
  wire  _GEN_716; // @[Execute.scala 206:23]
  wire  _GEN_717; // @[Execute.scala 206:23]
  wire  _GEN_718; // @[Execute.scala 206:23]
  wire  _GEN_719; // @[Execute.scala 206:23]
  wire  _T_131; // @[Execute.scala 206:14]
  wire  vecResult_45; // @[Execute.scala 206:23]
  wire  _GEN_721; // @[Execute.scala 206:23]
  wire  _GEN_722; // @[Execute.scala 206:23]
  wire  _GEN_723; // @[Execute.scala 206:23]
  wire  _GEN_724; // @[Execute.scala 206:23]
  wire  _GEN_725; // @[Execute.scala 206:23]
  wire  _GEN_726; // @[Execute.scala 206:23]
  wire  _GEN_727; // @[Execute.scala 206:23]
  wire  _GEN_728; // @[Execute.scala 206:23]
  wire  _GEN_729; // @[Execute.scala 206:23]
  wire  _GEN_730; // @[Execute.scala 206:23]
  wire  _GEN_731; // @[Execute.scala 206:23]
  wire  _GEN_732; // @[Execute.scala 206:23]
  wire  _GEN_733; // @[Execute.scala 206:23]
  wire  _GEN_734; // @[Execute.scala 206:23]
  wire  _GEN_735; // @[Execute.scala 206:23]
  wire  _T_132; // @[Execute.scala 206:14]
  wire  vecResult_46; // @[Execute.scala 206:23]
  wire  _GEN_737; // @[Execute.scala 206:23]
  wire  _GEN_738; // @[Execute.scala 206:23]
  wire  _GEN_739; // @[Execute.scala 206:23]
  wire  _GEN_740; // @[Execute.scala 206:23]
  wire  _GEN_741; // @[Execute.scala 206:23]
  wire  _GEN_742; // @[Execute.scala 206:23]
  wire  _GEN_743; // @[Execute.scala 206:23]
  wire  _GEN_744; // @[Execute.scala 206:23]
  wire  _GEN_745; // @[Execute.scala 206:23]
  wire  _GEN_746; // @[Execute.scala 206:23]
  wire  _GEN_747; // @[Execute.scala 206:23]
  wire  _GEN_748; // @[Execute.scala 206:23]
  wire  _GEN_749; // @[Execute.scala 206:23]
  wire  _GEN_750; // @[Execute.scala 206:23]
  wire  _GEN_751; // @[Execute.scala 206:23]
  wire  _T_133; // @[Execute.scala 206:14]
  wire  vecResult_47; // @[Execute.scala 206:23]
  wire  _GEN_753; // @[Execute.scala 206:23]
  wire  _GEN_754; // @[Execute.scala 206:23]
  wire  _GEN_755; // @[Execute.scala 206:23]
  wire  _GEN_756; // @[Execute.scala 206:23]
  wire  _GEN_757; // @[Execute.scala 206:23]
  wire  _GEN_758; // @[Execute.scala 206:23]
  wire  _GEN_759; // @[Execute.scala 206:23]
  wire  _GEN_760; // @[Execute.scala 206:23]
  wire  _GEN_761; // @[Execute.scala 206:23]
  wire  _GEN_762; // @[Execute.scala 206:23]
  wire  _GEN_763; // @[Execute.scala 206:23]
  wire  _GEN_764; // @[Execute.scala 206:23]
  wire  _GEN_765; // @[Execute.scala 206:23]
  wire  _GEN_766; // @[Execute.scala 206:23]
  wire  _GEN_767; // @[Execute.scala 206:23]
  wire  _T_134; // @[Execute.scala 206:14]
  wire  vecResult_48; // @[Execute.scala 206:23]
  wire  vecResult_49; // @[Execute.scala 206:23]
  wire  vecResult_50; // @[Execute.scala 206:23]
  wire  vecResult_51; // @[Execute.scala 206:23]
  wire  vecResult_52; // @[Execute.scala 206:23]
  wire  vecResult_53; // @[Execute.scala 206:23]
  wire  vecResult_54; // @[Execute.scala 206:23]
  wire  vecResult_55; // @[Execute.scala 206:23]
  wire  vecResult_56; // @[Execute.scala 206:23]
  wire  vecResult_57; // @[Execute.scala 206:23]
  wire  vecResult_58; // @[Execute.scala 206:23]
  wire  vecResult_59; // @[Execute.scala 206:23]
  wire  vecResult_60; // @[Execute.scala 206:23]
  wire  vecResult_61; // @[Execute.scala 206:23]
  wire  vecResult_62; // @[Execute.scala 206:23]
  wire  vecResult_63; // @[Execute.scala 206:23]
  wire [7:0] _T_141; // @[Execute.scala 213:32]
  wire [15:0] _T_149; // @[Execute.scala 213:32]
  wire [7:0] _T_156; // @[Execute.scala 213:32]
  wire [31:0] _T_165; // @[Execute.scala 213:32]
  wire [7:0] _T_172; // @[Execute.scala 213:32]
  wire [15:0] _T_180; // @[Execute.scala 213:32]
  wire [7:0] _T_187; // @[Execute.scala 213:32]
  wire [31:0] _T_196; // @[Execute.scala 213:32]
  wire [63:0] res; // @[Execute.scala 213:32]
  wire  _T_198; // @[Execute.scala 214:23]
  wire [63:0] _T_199; // @[Execute.scala 214:36]
  assign pos = {io_hw,4'h0}; // @[Cat.scala 29:58]
  assign _T_4 = 4'h2 == io_op; // @[Mux.scala 80:60]
  assign result = _T_4 ? io_rd : 64'h0; // @[Mux.scala 80:57]
  assign vecBools_0 = io_imm[0]; // @[Execute.scala 203:33]
  assign vecBools_1 = io_imm[1]; // @[Execute.scala 203:33]
  assign vecBools_2 = io_imm[2]; // @[Execute.scala 203:33]
  assign vecBools_3 = io_imm[3]; // @[Execute.scala 203:33]
  assign vecBools_4 = io_imm[4]; // @[Execute.scala 203:33]
  assign vecBools_5 = io_imm[5]; // @[Execute.scala 203:33]
  assign vecBools_6 = io_imm[6]; // @[Execute.scala 203:33]
  assign vecBools_7 = io_imm[7]; // @[Execute.scala 203:33]
  assign vecBools_8 = io_imm[8]; // @[Execute.scala 203:33]
  assign vecBools_9 = io_imm[9]; // @[Execute.scala 203:33]
  assign vecBools_10 = io_imm[10]; // @[Execute.scala 203:33]
  assign vecBools_11 = io_imm[11]; // @[Execute.scala 203:33]
  assign vecBools_12 = io_imm[12]; // @[Execute.scala 203:33]
  assign vecBools_13 = io_imm[13]; // @[Execute.scala 203:33]
  assign vecBools_14 = io_imm[14]; // @[Execute.scala 203:33]
  assign vecBools_15 = io_imm[15]; // @[Execute.scala 203:33]
  assign _T_86 = 6'h0 == pos; // @[Execute.scala 206:14]
  assign vecResult_0 = _T_86 ? vecBools_0 : result[0]; // @[Execute.scala 206:23]
  assign _GEN_1 = _T_86 ? vecBools_1 : result[1]; // @[Execute.scala 206:23]
  assign _GEN_2 = _T_86 ? vecBools_2 : result[2]; // @[Execute.scala 206:23]
  assign _GEN_3 = _T_86 ? vecBools_3 : result[3]; // @[Execute.scala 206:23]
  assign _GEN_4 = _T_86 ? vecBools_4 : result[4]; // @[Execute.scala 206:23]
  assign _GEN_5 = _T_86 ? vecBools_5 : result[5]; // @[Execute.scala 206:23]
  assign _GEN_6 = _T_86 ? vecBools_6 : result[6]; // @[Execute.scala 206:23]
  assign _GEN_7 = _T_86 ? vecBools_7 : result[7]; // @[Execute.scala 206:23]
  assign _GEN_8 = _T_86 ? vecBools_8 : result[8]; // @[Execute.scala 206:23]
  assign _GEN_9 = _T_86 ? vecBools_9 : result[9]; // @[Execute.scala 206:23]
  assign _GEN_10 = _T_86 ? vecBools_10 : result[10]; // @[Execute.scala 206:23]
  assign _GEN_11 = _T_86 ? vecBools_11 : result[11]; // @[Execute.scala 206:23]
  assign _GEN_12 = _T_86 ? vecBools_12 : result[12]; // @[Execute.scala 206:23]
  assign _GEN_13 = _T_86 ? vecBools_13 : result[13]; // @[Execute.scala 206:23]
  assign _GEN_14 = _T_86 ? vecBools_14 : result[14]; // @[Execute.scala 206:23]
  assign _GEN_15 = _T_86 ? vecBools_15 : result[15]; // @[Execute.scala 206:23]
  assign _T_87 = 6'h1 == pos; // @[Execute.scala 206:14]
  assign vecResult_1 = _T_87 ? vecBools_0 : _GEN_1; // @[Execute.scala 206:23]
  assign _GEN_17 = _T_87 ? vecBools_1 : _GEN_2; // @[Execute.scala 206:23]
  assign _GEN_18 = _T_87 ? vecBools_2 : _GEN_3; // @[Execute.scala 206:23]
  assign _GEN_19 = _T_87 ? vecBools_3 : _GEN_4; // @[Execute.scala 206:23]
  assign _GEN_20 = _T_87 ? vecBools_4 : _GEN_5; // @[Execute.scala 206:23]
  assign _GEN_21 = _T_87 ? vecBools_5 : _GEN_6; // @[Execute.scala 206:23]
  assign _GEN_22 = _T_87 ? vecBools_6 : _GEN_7; // @[Execute.scala 206:23]
  assign _GEN_23 = _T_87 ? vecBools_7 : _GEN_8; // @[Execute.scala 206:23]
  assign _GEN_24 = _T_87 ? vecBools_8 : _GEN_9; // @[Execute.scala 206:23]
  assign _GEN_25 = _T_87 ? vecBools_9 : _GEN_10; // @[Execute.scala 206:23]
  assign _GEN_26 = _T_87 ? vecBools_10 : _GEN_11; // @[Execute.scala 206:23]
  assign _GEN_27 = _T_87 ? vecBools_11 : _GEN_12; // @[Execute.scala 206:23]
  assign _GEN_28 = _T_87 ? vecBools_12 : _GEN_13; // @[Execute.scala 206:23]
  assign _GEN_29 = _T_87 ? vecBools_13 : _GEN_14; // @[Execute.scala 206:23]
  assign _GEN_30 = _T_87 ? vecBools_14 : _GEN_15; // @[Execute.scala 206:23]
  assign _GEN_31 = _T_87 ? vecBools_15 : result[16]; // @[Execute.scala 206:23]
  assign _T_88 = 6'h2 == pos; // @[Execute.scala 206:14]
  assign vecResult_2 = _T_88 ? vecBools_0 : _GEN_17; // @[Execute.scala 206:23]
  assign _GEN_33 = _T_88 ? vecBools_1 : _GEN_18; // @[Execute.scala 206:23]
  assign _GEN_34 = _T_88 ? vecBools_2 : _GEN_19; // @[Execute.scala 206:23]
  assign _GEN_35 = _T_88 ? vecBools_3 : _GEN_20; // @[Execute.scala 206:23]
  assign _GEN_36 = _T_88 ? vecBools_4 : _GEN_21; // @[Execute.scala 206:23]
  assign _GEN_37 = _T_88 ? vecBools_5 : _GEN_22; // @[Execute.scala 206:23]
  assign _GEN_38 = _T_88 ? vecBools_6 : _GEN_23; // @[Execute.scala 206:23]
  assign _GEN_39 = _T_88 ? vecBools_7 : _GEN_24; // @[Execute.scala 206:23]
  assign _GEN_40 = _T_88 ? vecBools_8 : _GEN_25; // @[Execute.scala 206:23]
  assign _GEN_41 = _T_88 ? vecBools_9 : _GEN_26; // @[Execute.scala 206:23]
  assign _GEN_42 = _T_88 ? vecBools_10 : _GEN_27; // @[Execute.scala 206:23]
  assign _GEN_43 = _T_88 ? vecBools_11 : _GEN_28; // @[Execute.scala 206:23]
  assign _GEN_44 = _T_88 ? vecBools_12 : _GEN_29; // @[Execute.scala 206:23]
  assign _GEN_45 = _T_88 ? vecBools_13 : _GEN_30; // @[Execute.scala 206:23]
  assign _GEN_46 = _T_88 ? vecBools_14 : _GEN_31; // @[Execute.scala 206:23]
  assign _GEN_47 = _T_88 ? vecBools_15 : result[17]; // @[Execute.scala 206:23]
  assign _T_89 = 6'h3 == pos; // @[Execute.scala 206:14]
  assign vecResult_3 = _T_89 ? vecBools_0 : _GEN_33; // @[Execute.scala 206:23]
  assign _GEN_49 = _T_89 ? vecBools_1 : _GEN_34; // @[Execute.scala 206:23]
  assign _GEN_50 = _T_89 ? vecBools_2 : _GEN_35; // @[Execute.scala 206:23]
  assign _GEN_51 = _T_89 ? vecBools_3 : _GEN_36; // @[Execute.scala 206:23]
  assign _GEN_52 = _T_89 ? vecBools_4 : _GEN_37; // @[Execute.scala 206:23]
  assign _GEN_53 = _T_89 ? vecBools_5 : _GEN_38; // @[Execute.scala 206:23]
  assign _GEN_54 = _T_89 ? vecBools_6 : _GEN_39; // @[Execute.scala 206:23]
  assign _GEN_55 = _T_89 ? vecBools_7 : _GEN_40; // @[Execute.scala 206:23]
  assign _GEN_56 = _T_89 ? vecBools_8 : _GEN_41; // @[Execute.scala 206:23]
  assign _GEN_57 = _T_89 ? vecBools_9 : _GEN_42; // @[Execute.scala 206:23]
  assign _GEN_58 = _T_89 ? vecBools_10 : _GEN_43; // @[Execute.scala 206:23]
  assign _GEN_59 = _T_89 ? vecBools_11 : _GEN_44; // @[Execute.scala 206:23]
  assign _GEN_60 = _T_89 ? vecBools_12 : _GEN_45; // @[Execute.scala 206:23]
  assign _GEN_61 = _T_89 ? vecBools_13 : _GEN_46; // @[Execute.scala 206:23]
  assign _GEN_62 = _T_89 ? vecBools_14 : _GEN_47; // @[Execute.scala 206:23]
  assign _GEN_63 = _T_89 ? vecBools_15 : result[18]; // @[Execute.scala 206:23]
  assign _T_90 = 6'h4 == pos; // @[Execute.scala 206:14]
  assign vecResult_4 = _T_90 ? vecBools_0 : _GEN_49; // @[Execute.scala 206:23]
  assign _GEN_65 = _T_90 ? vecBools_1 : _GEN_50; // @[Execute.scala 206:23]
  assign _GEN_66 = _T_90 ? vecBools_2 : _GEN_51; // @[Execute.scala 206:23]
  assign _GEN_67 = _T_90 ? vecBools_3 : _GEN_52; // @[Execute.scala 206:23]
  assign _GEN_68 = _T_90 ? vecBools_4 : _GEN_53; // @[Execute.scala 206:23]
  assign _GEN_69 = _T_90 ? vecBools_5 : _GEN_54; // @[Execute.scala 206:23]
  assign _GEN_70 = _T_90 ? vecBools_6 : _GEN_55; // @[Execute.scala 206:23]
  assign _GEN_71 = _T_90 ? vecBools_7 : _GEN_56; // @[Execute.scala 206:23]
  assign _GEN_72 = _T_90 ? vecBools_8 : _GEN_57; // @[Execute.scala 206:23]
  assign _GEN_73 = _T_90 ? vecBools_9 : _GEN_58; // @[Execute.scala 206:23]
  assign _GEN_74 = _T_90 ? vecBools_10 : _GEN_59; // @[Execute.scala 206:23]
  assign _GEN_75 = _T_90 ? vecBools_11 : _GEN_60; // @[Execute.scala 206:23]
  assign _GEN_76 = _T_90 ? vecBools_12 : _GEN_61; // @[Execute.scala 206:23]
  assign _GEN_77 = _T_90 ? vecBools_13 : _GEN_62; // @[Execute.scala 206:23]
  assign _GEN_78 = _T_90 ? vecBools_14 : _GEN_63; // @[Execute.scala 206:23]
  assign _GEN_79 = _T_90 ? vecBools_15 : result[19]; // @[Execute.scala 206:23]
  assign _T_91 = 6'h5 == pos; // @[Execute.scala 206:14]
  assign vecResult_5 = _T_91 ? vecBools_0 : _GEN_65; // @[Execute.scala 206:23]
  assign _GEN_81 = _T_91 ? vecBools_1 : _GEN_66; // @[Execute.scala 206:23]
  assign _GEN_82 = _T_91 ? vecBools_2 : _GEN_67; // @[Execute.scala 206:23]
  assign _GEN_83 = _T_91 ? vecBools_3 : _GEN_68; // @[Execute.scala 206:23]
  assign _GEN_84 = _T_91 ? vecBools_4 : _GEN_69; // @[Execute.scala 206:23]
  assign _GEN_85 = _T_91 ? vecBools_5 : _GEN_70; // @[Execute.scala 206:23]
  assign _GEN_86 = _T_91 ? vecBools_6 : _GEN_71; // @[Execute.scala 206:23]
  assign _GEN_87 = _T_91 ? vecBools_7 : _GEN_72; // @[Execute.scala 206:23]
  assign _GEN_88 = _T_91 ? vecBools_8 : _GEN_73; // @[Execute.scala 206:23]
  assign _GEN_89 = _T_91 ? vecBools_9 : _GEN_74; // @[Execute.scala 206:23]
  assign _GEN_90 = _T_91 ? vecBools_10 : _GEN_75; // @[Execute.scala 206:23]
  assign _GEN_91 = _T_91 ? vecBools_11 : _GEN_76; // @[Execute.scala 206:23]
  assign _GEN_92 = _T_91 ? vecBools_12 : _GEN_77; // @[Execute.scala 206:23]
  assign _GEN_93 = _T_91 ? vecBools_13 : _GEN_78; // @[Execute.scala 206:23]
  assign _GEN_94 = _T_91 ? vecBools_14 : _GEN_79; // @[Execute.scala 206:23]
  assign _GEN_95 = _T_91 ? vecBools_15 : result[20]; // @[Execute.scala 206:23]
  assign _T_92 = 6'h6 == pos; // @[Execute.scala 206:14]
  assign vecResult_6 = _T_92 ? vecBools_0 : _GEN_81; // @[Execute.scala 206:23]
  assign _GEN_97 = _T_92 ? vecBools_1 : _GEN_82; // @[Execute.scala 206:23]
  assign _GEN_98 = _T_92 ? vecBools_2 : _GEN_83; // @[Execute.scala 206:23]
  assign _GEN_99 = _T_92 ? vecBools_3 : _GEN_84; // @[Execute.scala 206:23]
  assign _GEN_100 = _T_92 ? vecBools_4 : _GEN_85; // @[Execute.scala 206:23]
  assign _GEN_101 = _T_92 ? vecBools_5 : _GEN_86; // @[Execute.scala 206:23]
  assign _GEN_102 = _T_92 ? vecBools_6 : _GEN_87; // @[Execute.scala 206:23]
  assign _GEN_103 = _T_92 ? vecBools_7 : _GEN_88; // @[Execute.scala 206:23]
  assign _GEN_104 = _T_92 ? vecBools_8 : _GEN_89; // @[Execute.scala 206:23]
  assign _GEN_105 = _T_92 ? vecBools_9 : _GEN_90; // @[Execute.scala 206:23]
  assign _GEN_106 = _T_92 ? vecBools_10 : _GEN_91; // @[Execute.scala 206:23]
  assign _GEN_107 = _T_92 ? vecBools_11 : _GEN_92; // @[Execute.scala 206:23]
  assign _GEN_108 = _T_92 ? vecBools_12 : _GEN_93; // @[Execute.scala 206:23]
  assign _GEN_109 = _T_92 ? vecBools_13 : _GEN_94; // @[Execute.scala 206:23]
  assign _GEN_110 = _T_92 ? vecBools_14 : _GEN_95; // @[Execute.scala 206:23]
  assign _GEN_111 = _T_92 ? vecBools_15 : result[21]; // @[Execute.scala 206:23]
  assign _T_93 = 6'h7 == pos; // @[Execute.scala 206:14]
  assign vecResult_7 = _T_93 ? vecBools_0 : _GEN_97; // @[Execute.scala 206:23]
  assign _GEN_113 = _T_93 ? vecBools_1 : _GEN_98; // @[Execute.scala 206:23]
  assign _GEN_114 = _T_93 ? vecBools_2 : _GEN_99; // @[Execute.scala 206:23]
  assign _GEN_115 = _T_93 ? vecBools_3 : _GEN_100; // @[Execute.scala 206:23]
  assign _GEN_116 = _T_93 ? vecBools_4 : _GEN_101; // @[Execute.scala 206:23]
  assign _GEN_117 = _T_93 ? vecBools_5 : _GEN_102; // @[Execute.scala 206:23]
  assign _GEN_118 = _T_93 ? vecBools_6 : _GEN_103; // @[Execute.scala 206:23]
  assign _GEN_119 = _T_93 ? vecBools_7 : _GEN_104; // @[Execute.scala 206:23]
  assign _GEN_120 = _T_93 ? vecBools_8 : _GEN_105; // @[Execute.scala 206:23]
  assign _GEN_121 = _T_93 ? vecBools_9 : _GEN_106; // @[Execute.scala 206:23]
  assign _GEN_122 = _T_93 ? vecBools_10 : _GEN_107; // @[Execute.scala 206:23]
  assign _GEN_123 = _T_93 ? vecBools_11 : _GEN_108; // @[Execute.scala 206:23]
  assign _GEN_124 = _T_93 ? vecBools_12 : _GEN_109; // @[Execute.scala 206:23]
  assign _GEN_125 = _T_93 ? vecBools_13 : _GEN_110; // @[Execute.scala 206:23]
  assign _GEN_126 = _T_93 ? vecBools_14 : _GEN_111; // @[Execute.scala 206:23]
  assign _GEN_127 = _T_93 ? vecBools_15 : result[22]; // @[Execute.scala 206:23]
  assign _T_94 = 6'h8 == pos; // @[Execute.scala 206:14]
  assign vecResult_8 = _T_94 ? vecBools_0 : _GEN_113; // @[Execute.scala 206:23]
  assign _GEN_129 = _T_94 ? vecBools_1 : _GEN_114; // @[Execute.scala 206:23]
  assign _GEN_130 = _T_94 ? vecBools_2 : _GEN_115; // @[Execute.scala 206:23]
  assign _GEN_131 = _T_94 ? vecBools_3 : _GEN_116; // @[Execute.scala 206:23]
  assign _GEN_132 = _T_94 ? vecBools_4 : _GEN_117; // @[Execute.scala 206:23]
  assign _GEN_133 = _T_94 ? vecBools_5 : _GEN_118; // @[Execute.scala 206:23]
  assign _GEN_134 = _T_94 ? vecBools_6 : _GEN_119; // @[Execute.scala 206:23]
  assign _GEN_135 = _T_94 ? vecBools_7 : _GEN_120; // @[Execute.scala 206:23]
  assign _GEN_136 = _T_94 ? vecBools_8 : _GEN_121; // @[Execute.scala 206:23]
  assign _GEN_137 = _T_94 ? vecBools_9 : _GEN_122; // @[Execute.scala 206:23]
  assign _GEN_138 = _T_94 ? vecBools_10 : _GEN_123; // @[Execute.scala 206:23]
  assign _GEN_139 = _T_94 ? vecBools_11 : _GEN_124; // @[Execute.scala 206:23]
  assign _GEN_140 = _T_94 ? vecBools_12 : _GEN_125; // @[Execute.scala 206:23]
  assign _GEN_141 = _T_94 ? vecBools_13 : _GEN_126; // @[Execute.scala 206:23]
  assign _GEN_142 = _T_94 ? vecBools_14 : _GEN_127; // @[Execute.scala 206:23]
  assign _GEN_143 = _T_94 ? vecBools_15 : result[23]; // @[Execute.scala 206:23]
  assign _T_95 = 6'h9 == pos; // @[Execute.scala 206:14]
  assign vecResult_9 = _T_95 ? vecBools_0 : _GEN_129; // @[Execute.scala 206:23]
  assign _GEN_145 = _T_95 ? vecBools_1 : _GEN_130; // @[Execute.scala 206:23]
  assign _GEN_146 = _T_95 ? vecBools_2 : _GEN_131; // @[Execute.scala 206:23]
  assign _GEN_147 = _T_95 ? vecBools_3 : _GEN_132; // @[Execute.scala 206:23]
  assign _GEN_148 = _T_95 ? vecBools_4 : _GEN_133; // @[Execute.scala 206:23]
  assign _GEN_149 = _T_95 ? vecBools_5 : _GEN_134; // @[Execute.scala 206:23]
  assign _GEN_150 = _T_95 ? vecBools_6 : _GEN_135; // @[Execute.scala 206:23]
  assign _GEN_151 = _T_95 ? vecBools_7 : _GEN_136; // @[Execute.scala 206:23]
  assign _GEN_152 = _T_95 ? vecBools_8 : _GEN_137; // @[Execute.scala 206:23]
  assign _GEN_153 = _T_95 ? vecBools_9 : _GEN_138; // @[Execute.scala 206:23]
  assign _GEN_154 = _T_95 ? vecBools_10 : _GEN_139; // @[Execute.scala 206:23]
  assign _GEN_155 = _T_95 ? vecBools_11 : _GEN_140; // @[Execute.scala 206:23]
  assign _GEN_156 = _T_95 ? vecBools_12 : _GEN_141; // @[Execute.scala 206:23]
  assign _GEN_157 = _T_95 ? vecBools_13 : _GEN_142; // @[Execute.scala 206:23]
  assign _GEN_158 = _T_95 ? vecBools_14 : _GEN_143; // @[Execute.scala 206:23]
  assign _GEN_159 = _T_95 ? vecBools_15 : result[24]; // @[Execute.scala 206:23]
  assign _T_96 = 6'ha == pos; // @[Execute.scala 206:14]
  assign vecResult_10 = _T_96 ? vecBools_0 : _GEN_145; // @[Execute.scala 206:23]
  assign _GEN_161 = _T_96 ? vecBools_1 : _GEN_146; // @[Execute.scala 206:23]
  assign _GEN_162 = _T_96 ? vecBools_2 : _GEN_147; // @[Execute.scala 206:23]
  assign _GEN_163 = _T_96 ? vecBools_3 : _GEN_148; // @[Execute.scala 206:23]
  assign _GEN_164 = _T_96 ? vecBools_4 : _GEN_149; // @[Execute.scala 206:23]
  assign _GEN_165 = _T_96 ? vecBools_5 : _GEN_150; // @[Execute.scala 206:23]
  assign _GEN_166 = _T_96 ? vecBools_6 : _GEN_151; // @[Execute.scala 206:23]
  assign _GEN_167 = _T_96 ? vecBools_7 : _GEN_152; // @[Execute.scala 206:23]
  assign _GEN_168 = _T_96 ? vecBools_8 : _GEN_153; // @[Execute.scala 206:23]
  assign _GEN_169 = _T_96 ? vecBools_9 : _GEN_154; // @[Execute.scala 206:23]
  assign _GEN_170 = _T_96 ? vecBools_10 : _GEN_155; // @[Execute.scala 206:23]
  assign _GEN_171 = _T_96 ? vecBools_11 : _GEN_156; // @[Execute.scala 206:23]
  assign _GEN_172 = _T_96 ? vecBools_12 : _GEN_157; // @[Execute.scala 206:23]
  assign _GEN_173 = _T_96 ? vecBools_13 : _GEN_158; // @[Execute.scala 206:23]
  assign _GEN_174 = _T_96 ? vecBools_14 : _GEN_159; // @[Execute.scala 206:23]
  assign _GEN_175 = _T_96 ? vecBools_15 : result[25]; // @[Execute.scala 206:23]
  assign _T_97 = 6'hb == pos; // @[Execute.scala 206:14]
  assign vecResult_11 = _T_97 ? vecBools_0 : _GEN_161; // @[Execute.scala 206:23]
  assign _GEN_177 = _T_97 ? vecBools_1 : _GEN_162; // @[Execute.scala 206:23]
  assign _GEN_178 = _T_97 ? vecBools_2 : _GEN_163; // @[Execute.scala 206:23]
  assign _GEN_179 = _T_97 ? vecBools_3 : _GEN_164; // @[Execute.scala 206:23]
  assign _GEN_180 = _T_97 ? vecBools_4 : _GEN_165; // @[Execute.scala 206:23]
  assign _GEN_181 = _T_97 ? vecBools_5 : _GEN_166; // @[Execute.scala 206:23]
  assign _GEN_182 = _T_97 ? vecBools_6 : _GEN_167; // @[Execute.scala 206:23]
  assign _GEN_183 = _T_97 ? vecBools_7 : _GEN_168; // @[Execute.scala 206:23]
  assign _GEN_184 = _T_97 ? vecBools_8 : _GEN_169; // @[Execute.scala 206:23]
  assign _GEN_185 = _T_97 ? vecBools_9 : _GEN_170; // @[Execute.scala 206:23]
  assign _GEN_186 = _T_97 ? vecBools_10 : _GEN_171; // @[Execute.scala 206:23]
  assign _GEN_187 = _T_97 ? vecBools_11 : _GEN_172; // @[Execute.scala 206:23]
  assign _GEN_188 = _T_97 ? vecBools_12 : _GEN_173; // @[Execute.scala 206:23]
  assign _GEN_189 = _T_97 ? vecBools_13 : _GEN_174; // @[Execute.scala 206:23]
  assign _GEN_190 = _T_97 ? vecBools_14 : _GEN_175; // @[Execute.scala 206:23]
  assign _GEN_191 = _T_97 ? vecBools_15 : result[26]; // @[Execute.scala 206:23]
  assign _T_98 = 6'hc == pos; // @[Execute.scala 206:14]
  assign vecResult_12 = _T_98 ? vecBools_0 : _GEN_177; // @[Execute.scala 206:23]
  assign _GEN_193 = _T_98 ? vecBools_1 : _GEN_178; // @[Execute.scala 206:23]
  assign _GEN_194 = _T_98 ? vecBools_2 : _GEN_179; // @[Execute.scala 206:23]
  assign _GEN_195 = _T_98 ? vecBools_3 : _GEN_180; // @[Execute.scala 206:23]
  assign _GEN_196 = _T_98 ? vecBools_4 : _GEN_181; // @[Execute.scala 206:23]
  assign _GEN_197 = _T_98 ? vecBools_5 : _GEN_182; // @[Execute.scala 206:23]
  assign _GEN_198 = _T_98 ? vecBools_6 : _GEN_183; // @[Execute.scala 206:23]
  assign _GEN_199 = _T_98 ? vecBools_7 : _GEN_184; // @[Execute.scala 206:23]
  assign _GEN_200 = _T_98 ? vecBools_8 : _GEN_185; // @[Execute.scala 206:23]
  assign _GEN_201 = _T_98 ? vecBools_9 : _GEN_186; // @[Execute.scala 206:23]
  assign _GEN_202 = _T_98 ? vecBools_10 : _GEN_187; // @[Execute.scala 206:23]
  assign _GEN_203 = _T_98 ? vecBools_11 : _GEN_188; // @[Execute.scala 206:23]
  assign _GEN_204 = _T_98 ? vecBools_12 : _GEN_189; // @[Execute.scala 206:23]
  assign _GEN_205 = _T_98 ? vecBools_13 : _GEN_190; // @[Execute.scala 206:23]
  assign _GEN_206 = _T_98 ? vecBools_14 : _GEN_191; // @[Execute.scala 206:23]
  assign _GEN_207 = _T_98 ? vecBools_15 : result[27]; // @[Execute.scala 206:23]
  assign _T_99 = 6'hd == pos; // @[Execute.scala 206:14]
  assign vecResult_13 = _T_99 ? vecBools_0 : _GEN_193; // @[Execute.scala 206:23]
  assign _GEN_209 = _T_99 ? vecBools_1 : _GEN_194; // @[Execute.scala 206:23]
  assign _GEN_210 = _T_99 ? vecBools_2 : _GEN_195; // @[Execute.scala 206:23]
  assign _GEN_211 = _T_99 ? vecBools_3 : _GEN_196; // @[Execute.scala 206:23]
  assign _GEN_212 = _T_99 ? vecBools_4 : _GEN_197; // @[Execute.scala 206:23]
  assign _GEN_213 = _T_99 ? vecBools_5 : _GEN_198; // @[Execute.scala 206:23]
  assign _GEN_214 = _T_99 ? vecBools_6 : _GEN_199; // @[Execute.scala 206:23]
  assign _GEN_215 = _T_99 ? vecBools_7 : _GEN_200; // @[Execute.scala 206:23]
  assign _GEN_216 = _T_99 ? vecBools_8 : _GEN_201; // @[Execute.scala 206:23]
  assign _GEN_217 = _T_99 ? vecBools_9 : _GEN_202; // @[Execute.scala 206:23]
  assign _GEN_218 = _T_99 ? vecBools_10 : _GEN_203; // @[Execute.scala 206:23]
  assign _GEN_219 = _T_99 ? vecBools_11 : _GEN_204; // @[Execute.scala 206:23]
  assign _GEN_220 = _T_99 ? vecBools_12 : _GEN_205; // @[Execute.scala 206:23]
  assign _GEN_221 = _T_99 ? vecBools_13 : _GEN_206; // @[Execute.scala 206:23]
  assign _GEN_222 = _T_99 ? vecBools_14 : _GEN_207; // @[Execute.scala 206:23]
  assign _GEN_223 = _T_99 ? vecBools_15 : result[28]; // @[Execute.scala 206:23]
  assign _T_100 = 6'he == pos; // @[Execute.scala 206:14]
  assign vecResult_14 = _T_100 ? vecBools_0 : _GEN_209; // @[Execute.scala 206:23]
  assign _GEN_225 = _T_100 ? vecBools_1 : _GEN_210; // @[Execute.scala 206:23]
  assign _GEN_226 = _T_100 ? vecBools_2 : _GEN_211; // @[Execute.scala 206:23]
  assign _GEN_227 = _T_100 ? vecBools_3 : _GEN_212; // @[Execute.scala 206:23]
  assign _GEN_228 = _T_100 ? vecBools_4 : _GEN_213; // @[Execute.scala 206:23]
  assign _GEN_229 = _T_100 ? vecBools_5 : _GEN_214; // @[Execute.scala 206:23]
  assign _GEN_230 = _T_100 ? vecBools_6 : _GEN_215; // @[Execute.scala 206:23]
  assign _GEN_231 = _T_100 ? vecBools_7 : _GEN_216; // @[Execute.scala 206:23]
  assign _GEN_232 = _T_100 ? vecBools_8 : _GEN_217; // @[Execute.scala 206:23]
  assign _GEN_233 = _T_100 ? vecBools_9 : _GEN_218; // @[Execute.scala 206:23]
  assign _GEN_234 = _T_100 ? vecBools_10 : _GEN_219; // @[Execute.scala 206:23]
  assign _GEN_235 = _T_100 ? vecBools_11 : _GEN_220; // @[Execute.scala 206:23]
  assign _GEN_236 = _T_100 ? vecBools_12 : _GEN_221; // @[Execute.scala 206:23]
  assign _GEN_237 = _T_100 ? vecBools_13 : _GEN_222; // @[Execute.scala 206:23]
  assign _GEN_238 = _T_100 ? vecBools_14 : _GEN_223; // @[Execute.scala 206:23]
  assign _GEN_239 = _T_100 ? vecBools_15 : result[29]; // @[Execute.scala 206:23]
  assign _T_101 = 6'hf == pos; // @[Execute.scala 206:14]
  assign vecResult_15 = _T_101 ? vecBools_0 : _GEN_225; // @[Execute.scala 206:23]
  assign _GEN_241 = _T_101 ? vecBools_1 : _GEN_226; // @[Execute.scala 206:23]
  assign _GEN_242 = _T_101 ? vecBools_2 : _GEN_227; // @[Execute.scala 206:23]
  assign _GEN_243 = _T_101 ? vecBools_3 : _GEN_228; // @[Execute.scala 206:23]
  assign _GEN_244 = _T_101 ? vecBools_4 : _GEN_229; // @[Execute.scala 206:23]
  assign _GEN_245 = _T_101 ? vecBools_5 : _GEN_230; // @[Execute.scala 206:23]
  assign _GEN_246 = _T_101 ? vecBools_6 : _GEN_231; // @[Execute.scala 206:23]
  assign _GEN_247 = _T_101 ? vecBools_7 : _GEN_232; // @[Execute.scala 206:23]
  assign _GEN_248 = _T_101 ? vecBools_8 : _GEN_233; // @[Execute.scala 206:23]
  assign _GEN_249 = _T_101 ? vecBools_9 : _GEN_234; // @[Execute.scala 206:23]
  assign _GEN_250 = _T_101 ? vecBools_10 : _GEN_235; // @[Execute.scala 206:23]
  assign _GEN_251 = _T_101 ? vecBools_11 : _GEN_236; // @[Execute.scala 206:23]
  assign _GEN_252 = _T_101 ? vecBools_12 : _GEN_237; // @[Execute.scala 206:23]
  assign _GEN_253 = _T_101 ? vecBools_13 : _GEN_238; // @[Execute.scala 206:23]
  assign _GEN_254 = _T_101 ? vecBools_14 : _GEN_239; // @[Execute.scala 206:23]
  assign _GEN_255 = _T_101 ? vecBools_15 : result[30]; // @[Execute.scala 206:23]
  assign _T_102 = 6'h10 == pos; // @[Execute.scala 206:14]
  assign vecResult_16 = _T_102 ? vecBools_0 : _GEN_241; // @[Execute.scala 206:23]
  assign _GEN_257 = _T_102 ? vecBools_1 : _GEN_242; // @[Execute.scala 206:23]
  assign _GEN_258 = _T_102 ? vecBools_2 : _GEN_243; // @[Execute.scala 206:23]
  assign _GEN_259 = _T_102 ? vecBools_3 : _GEN_244; // @[Execute.scala 206:23]
  assign _GEN_260 = _T_102 ? vecBools_4 : _GEN_245; // @[Execute.scala 206:23]
  assign _GEN_261 = _T_102 ? vecBools_5 : _GEN_246; // @[Execute.scala 206:23]
  assign _GEN_262 = _T_102 ? vecBools_6 : _GEN_247; // @[Execute.scala 206:23]
  assign _GEN_263 = _T_102 ? vecBools_7 : _GEN_248; // @[Execute.scala 206:23]
  assign _GEN_264 = _T_102 ? vecBools_8 : _GEN_249; // @[Execute.scala 206:23]
  assign _GEN_265 = _T_102 ? vecBools_9 : _GEN_250; // @[Execute.scala 206:23]
  assign _GEN_266 = _T_102 ? vecBools_10 : _GEN_251; // @[Execute.scala 206:23]
  assign _GEN_267 = _T_102 ? vecBools_11 : _GEN_252; // @[Execute.scala 206:23]
  assign _GEN_268 = _T_102 ? vecBools_12 : _GEN_253; // @[Execute.scala 206:23]
  assign _GEN_269 = _T_102 ? vecBools_13 : _GEN_254; // @[Execute.scala 206:23]
  assign _GEN_270 = _T_102 ? vecBools_14 : _GEN_255; // @[Execute.scala 206:23]
  assign _GEN_271 = _T_102 ? vecBools_15 : result[31]; // @[Execute.scala 206:23]
  assign _T_103 = 6'h11 == pos; // @[Execute.scala 206:14]
  assign vecResult_17 = _T_103 ? vecBools_0 : _GEN_257; // @[Execute.scala 206:23]
  assign _GEN_273 = _T_103 ? vecBools_1 : _GEN_258; // @[Execute.scala 206:23]
  assign _GEN_274 = _T_103 ? vecBools_2 : _GEN_259; // @[Execute.scala 206:23]
  assign _GEN_275 = _T_103 ? vecBools_3 : _GEN_260; // @[Execute.scala 206:23]
  assign _GEN_276 = _T_103 ? vecBools_4 : _GEN_261; // @[Execute.scala 206:23]
  assign _GEN_277 = _T_103 ? vecBools_5 : _GEN_262; // @[Execute.scala 206:23]
  assign _GEN_278 = _T_103 ? vecBools_6 : _GEN_263; // @[Execute.scala 206:23]
  assign _GEN_279 = _T_103 ? vecBools_7 : _GEN_264; // @[Execute.scala 206:23]
  assign _GEN_280 = _T_103 ? vecBools_8 : _GEN_265; // @[Execute.scala 206:23]
  assign _GEN_281 = _T_103 ? vecBools_9 : _GEN_266; // @[Execute.scala 206:23]
  assign _GEN_282 = _T_103 ? vecBools_10 : _GEN_267; // @[Execute.scala 206:23]
  assign _GEN_283 = _T_103 ? vecBools_11 : _GEN_268; // @[Execute.scala 206:23]
  assign _GEN_284 = _T_103 ? vecBools_12 : _GEN_269; // @[Execute.scala 206:23]
  assign _GEN_285 = _T_103 ? vecBools_13 : _GEN_270; // @[Execute.scala 206:23]
  assign _GEN_286 = _T_103 ? vecBools_14 : _GEN_271; // @[Execute.scala 206:23]
  assign _GEN_287 = _T_103 ? vecBools_15 : result[32]; // @[Execute.scala 206:23]
  assign _T_104 = 6'h12 == pos; // @[Execute.scala 206:14]
  assign vecResult_18 = _T_104 ? vecBools_0 : _GEN_273; // @[Execute.scala 206:23]
  assign _GEN_289 = _T_104 ? vecBools_1 : _GEN_274; // @[Execute.scala 206:23]
  assign _GEN_290 = _T_104 ? vecBools_2 : _GEN_275; // @[Execute.scala 206:23]
  assign _GEN_291 = _T_104 ? vecBools_3 : _GEN_276; // @[Execute.scala 206:23]
  assign _GEN_292 = _T_104 ? vecBools_4 : _GEN_277; // @[Execute.scala 206:23]
  assign _GEN_293 = _T_104 ? vecBools_5 : _GEN_278; // @[Execute.scala 206:23]
  assign _GEN_294 = _T_104 ? vecBools_6 : _GEN_279; // @[Execute.scala 206:23]
  assign _GEN_295 = _T_104 ? vecBools_7 : _GEN_280; // @[Execute.scala 206:23]
  assign _GEN_296 = _T_104 ? vecBools_8 : _GEN_281; // @[Execute.scala 206:23]
  assign _GEN_297 = _T_104 ? vecBools_9 : _GEN_282; // @[Execute.scala 206:23]
  assign _GEN_298 = _T_104 ? vecBools_10 : _GEN_283; // @[Execute.scala 206:23]
  assign _GEN_299 = _T_104 ? vecBools_11 : _GEN_284; // @[Execute.scala 206:23]
  assign _GEN_300 = _T_104 ? vecBools_12 : _GEN_285; // @[Execute.scala 206:23]
  assign _GEN_301 = _T_104 ? vecBools_13 : _GEN_286; // @[Execute.scala 206:23]
  assign _GEN_302 = _T_104 ? vecBools_14 : _GEN_287; // @[Execute.scala 206:23]
  assign _GEN_303 = _T_104 ? vecBools_15 : result[33]; // @[Execute.scala 206:23]
  assign _T_105 = 6'h13 == pos; // @[Execute.scala 206:14]
  assign vecResult_19 = _T_105 ? vecBools_0 : _GEN_289; // @[Execute.scala 206:23]
  assign _GEN_305 = _T_105 ? vecBools_1 : _GEN_290; // @[Execute.scala 206:23]
  assign _GEN_306 = _T_105 ? vecBools_2 : _GEN_291; // @[Execute.scala 206:23]
  assign _GEN_307 = _T_105 ? vecBools_3 : _GEN_292; // @[Execute.scala 206:23]
  assign _GEN_308 = _T_105 ? vecBools_4 : _GEN_293; // @[Execute.scala 206:23]
  assign _GEN_309 = _T_105 ? vecBools_5 : _GEN_294; // @[Execute.scala 206:23]
  assign _GEN_310 = _T_105 ? vecBools_6 : _GEN_295; // @[Execute.scala 206:23]
  assign _GEN_311 = _T_105 ? vecBools_7 : _GEN_296; // @[Execute.scala 206:23]
  assign _GEN_312 = _T_105 ? vecBools_8 : _GEN_297; // @[Execute.scala 206:23]
  assign _GEN_313 = _T_105 ? vecBools_9 : _GEN_298; // @[Execute.scala 206:23]
  assign _GEN_314 = _T_105 ? vecBools_10 : _GEN_299; // @[Execute.scala 206:23]
  assign _GEN_315 = _T_105 ? vecBools_11 : _GEN_300; // @[Execute.scala 206:23]
  assign _GEN_316 = _T_105 ? vecBools_12 : _GEN_301; // @[Execute.scala 206:23]
  assign _GEN_317 = _T_105 ? vecBools_13 : _GEN_302; // @[Execute.scala 206:23]
  assign _GEN_318 = _T_105 ? vecBools_14 : _GEN_303; // @[Execute.scala 206:23]
  assign _GEN_319 = _T_105 ? vecBools_15 : result[34]; // @[Execute.scala 206:23]
  assign _T_106 = 6'h14 == pos; // @[Execute.scala 206:14]
  assign vecResult_20 = _T_106 ? vecBools_0 : _GEN_305; // @[Execute.scala 206:23]
  assign _GEN_321 = _T_106 ? vecBools_1 : _GEN_306; // @[Execute.scala 206:23]
  assign _GEN_322 = _T_106 ? vecBools_2 : _GEN_307; // @[Execute.scala 206:23]
  assign _GEN_323 = _T_106 ? vecBools_3 : _GEN_308; // @[Execute.scala 206:23]
  assign _GEN_324 = _T_106 ? vecBools_4 : _GEN_309; // @[Execute.scala 206:23]
  assign _GEN_325 = _T_106 ? vecBools_5 : _GEN_310; // @[Execute.scala 206:23]
  assign _GEN_326 = _T_106 ? vecBools_6 : _GEN_311; // @[Execute.scala 206:23]
  assign _GEN_327 = _T_106 ? vecBools_7 : _GEN_312; // @[Execute.scala 206:23]
  assign _GEN_328 = _T_106 ? vecBools_8 : _GEN_313; // @[Execute.scala 206:23]
  assign _GEN_329 = _T_106 ? vecBools_9 : _GEN_314; // @[Execute.scala 206:23]
  assign _GEN_330 = _T_106 ? vecBools_10 : _GEN_315; // @[Execute.scala 206:23]
  assign _GEN_331 = _T_106 ? vecBools_11 : _GEN_316; // @[Execute.scala 206:23]
  assign _GEN_332 = _T_106 ? vecBools_12 : _GEN_317; // @[Execute.scala 206:23]
  assign _GEN_333 = _T_106 ? vecBools_13 : _GEN_318; // @[Execute.scala 206:23]
  assign _GEN_334 = _T_106 ? vecBools_14 : _GEN_319; // @[Execute.scala 206:23]
  assign _GEN_335 = _T_106 ? vecBools_15 : result[35]; // @[Execute.scala 206:23]
  assign _T_107 = 6'h15 == pos; // @[Execute.scala 206:14]
  assign vecResult_21 = _T_107 ? vecBools_0 : _GEN_321; // @[Execute.scala 206:23]
  assign _GEN_337 = _T_107 ? vecBools_1 : _GEN_322; // @[Execute.scala 206:23]
  assign _GEN_338 = _T_107 ? vecBools_2 : _GEN_323; // @[Execute.scala 206:23]
  assign _GEN_339 = _T_107 ? vecBools_3 : _GEN_324; // @[Execute.scala 206:23]
  assign _GEN_340 = _T_107 ? vecBools_4 : _GEN_325; // @[Execute.scala 206:23]
  assign _GEN_341 = _T_107 ? vecBools_5 : _GEN_326; // @[Execute.scala 206:23]
  assign _GEN_342 = _T_107 ? vecBools_6 : _GEN_327; // @[Execute.scala 206:23]
  assign _GEN_343 = _T_107 ? vecBools_7 : _GEN_328; // @[Execute.scala 206:23]
  assign _GEN_344 = _T_107 ? vecBools_8 : _GEN_329; // @[Execute.scala 206:23]
  assign _GEN_345 = _T_107 ? vecBools_9 : _GEN_330; // @[Execute.scala 206:23]
  assign _GEN_346 = _T_107 ? vecBools_10 : _GEN_331; // @[Execute.scala 206:23]
  assign _GEN_347 = _T_107 ? vecBools_11 : _GEN_332; // @[Execute.scala 206:23]
  assign _GEN_348 = _T_107 ? vecBools_12 : _GEN_333; // @[Execute.scala 206:23]
  assign _GEN_349 = _T_107 ? vecBools_13 : _GEN_334; // @[Execute.scala 206:23]
  assign _GEN_350 = _T_107 ? vecBools_14 : _GEN_335; // @[Execute.scala 206:23]
  assign _GEN_351 = _T_107 ? vecBools_15 : result[36]; // @[Execute.scala 206:23]
  assign _T_108 = 6'h16 == pos; // @[Execute.scala 206:14]
  assign vecResult_22 = _T_108 ? vecBools_0 : _GEN_337; // @[Execute.scala 206:23]
  assign _GEN_353 = _T_108 ? vecBools_1 : _GEN_338; // @[Execute.scala 206:23]
  assign _GEN_354 = _T_108 ? vecBools_2 : _GEN_339; // @[Execute.scala 206:23]
  assign _GEN_355 = _T_108 ? vecBools_3 : _GEN_340; // @[Execute.scala 206:23]
  assign _GEN_356 = _T_108 ? vecBools_4 : _GEN_341; // @[Execute.scala 206:23]
  assign _GEN_357 = _T_108 ? vecBools_5 : _GEN_342; // @[Execute.scala 206:23]
  assign _GEN_358 = _T_108 ? vecBools_6 : _GEN_343; // @[Execute.scala 206:23]
  assign _GEN_359 = _T_108 ? vecBools_7 : _GEN_344; // @[Execute.scala 206:23]
  assign _GEN_360 = _T_108 ? vecBools_8 : _GEN_345; // @[Execute.scala 206:23]
  assign _GEN_361 = _T_108 ? vecBools_9 : _GEN_346; // @[Execute.scala 206:23]
  assign _GEN_362 = _T_108 ? vecBools_10 : _GEN_347; // @[Execute.scala 206:23]
  assign _GEN_363 = _T_108 ? vecBools_11 : _GEN_348; // @[Execute.scala 206:23]
  assign _GEN_364 = _T_108 ? vecBools_12 : _GEN_349; // @[Execute.scala 206:23]
  assign _GEN_365 = _T_108 ? vecBools_13 : _GEN_350; // @[Execute.scala 206:23]
  assign _GEN_366 = _T_108 ? vecBools_14 : _GEN_351; // @[Execute.scala 206:23]
  assign _GEN_367 = _T_108 ? vecBools_15 : result[37]; // @[Execute.scala 206:23]
  assign _T_109 = 6'h17 == pos; // @[Execute.scala 206:14]
  assign vecResult_23 = _T_109 ? vecBools_0 : _GEN_353; // @[Execute.scala 206:23]
  assign _GEN_369 = _T_109 ? vecBools_1 : _GEN_354; // @[Execute.scala 206:23]
  assign _GEN_370 = _T_109 ? vecBools_2 : _GEN_355; // @[Execute.scala 206:23]
  assign _GEN_371 = _T_109 ? vecBools_3 : _GEN_356; // @[Execute.scala 206:23]
  assign _GEN_372 = _T_109 ? vecBools_4 : _GEN_357; // @[Execute.scala 206:23]
  assign _GEN_373 = _T_109 ? vecBools_5 : _GEN_358; // @[Execute.scala 206:23]
  assign _GEN_374 = _T_109 ? vecBools_6 : _GEN_359; // @[Execute.scala 206:23]
  assign _GEN_375 = _T_109 ? vecBools_7 : _GEN_360; // @[Execute.scala 206:23]
  assign _GEN_376 = _T_109 ? vecBools_8 : _GEN_361; // @[Execute.scala 206:23]
  assign _GEN_377 = _T_109 ? vecBools_9 : _GEN_362; // @[Execute.scala 206:23]
  assign _GEN_378 = _T_109 ? vecBools_10 : _GEN_363; // @[Execute.scala 206:23]
  assign _GEN_379 = _T_109 ? vecBools_11 : _GEN_364; // @[Execute.scala 206:23]
  assign _GEN_380 = _T_109 ? vecBools_12 : _GEN_365; // @[Execute.scala 206:23]
  assign _GEN_381 = _T_109 ? vecBools_13 : _GEN_366; // @[Execute.scala 206:23]
  assign _GEN_382 = _T_109 ? vecBools_14 : _GEN_367; // @[Execute.scala 206:23]
  assign _GEN_383 = _T_109 ? vecBools_15 : result[38]; // @[Execute.scala 206:23]
  assign _T_110 = 6'h18 == pos; // @[Execute.scala 206:14]
  assign vecResult_24 = _T_110 ? vecBools_0 : _GEN_369; // @[Execute.scala 206:23]
  assign _GEN_385 = _T_110 ? vecBools_1 : _GEN_370; // @[Execute.scala 206:23]
  assign _GEN_386 = _T_110 ? vecBools_2 : _GEN_371; // @[Execute.scala 206:23]
  assign _GEN_387 = _T_110 ? vecBools_3 : _GEN_372; // @[Execute.scala 206:23]
  assign _GEN_388 = _T_110 ? vecBools_4 : _GEN_373; // @[Execute.scala 206:23]
  assign _GEN_389 = _T_110 ? vecBools_5 : _GEN_374; // @[Execute.scala 206:23]
  assign _GEN_390 = _T_110 ? vecBools_6 : _GEN_375; // @[Execute.scala 206:23]
  assign _GEN_391 = _T_110 ? vecBools_7 : _GEN_376; // @[Execute.scala 206:23]
  assign _GEN_392 = _T_110 ? vecBools_8 : _GEN_377; // @[Execute.scala 206:23]
  assign _GEN_393 = _T_110 ? vecBools_9 : _GEN_378; // @[Execute.scala 206:23]
  assign _GEN_394 = _T_110 ? vecBools_10 : _GEN_379; // @[Execute.scala 206:23]
  assign _GEN_395 = _T_110 ? vecBools_11 : _GEN_380; // @[Execute.scala 206:23]
  assign _GEN_396 = _T_110 ? vecBools_12 : _GEN_381; // @[Execute.scala 206:23]
  assign _GEN_397 = _T_110 ? vecBools_13 : _GEN_382; // @[Execute.scala 206:23]
  assign _GEN_398 = _T_110 ? vecBools_14 : _GEN_383; // @[Execute.scala 206:23]
  assign _GEN_399 = _T_110 ? vecBools_15 : result[39]; // @[Execute.scala 206:23]
  assign _T_111 = 6'h19 == pos; // @[Execute.scala 206:14]
  assign vecResult_25 = _T_111 ? vecBools_0 : _GEN_385; // @[Execute.scala 206:23]
  assign _GEN_401 = _T_111 ? vecBools_1 : _GEN_386; // @[Execute.scala 206:23]
  assign _GEN_402 = _T_111 ? vecBools_2 : _GEN_387; // @[Execute.scala 206:23]
  assign _GEN_403 = _T_111 ? vecBools_3 : _GEN_388; // @[Execute.scala 206:23]
  assign _GEN_404 = _T_111 ? vecBools_4 : _GEN_389; // @[Execute.scala 206:23]
  assign _GEN_405 = _T_111 ? vecBools_5 : _GEN_390; // @[Execute.scala 206:23]
  assign _GEN_406 = _T_111 ? vecBools_6 : _GEN_391; // @[Execute.scala 206:23]
  assign _GEN_407 = _T_111 ? vecBools_7 : _GEN_392; // @[Execute.scala 206:23]
  assign _GEN_408 = _T_111 ? vecBools_8 : _GEN_393; // @[Execute.scala 206:23]
  assign _GEN_409 = _T_111 ? vecBools_9 : _GEN_394; // @[Execute.scala 206:23]
  assign _GEN_410 = _T_111 ? vecBools_10 : _GEN_395; // @[Execute.scala 206:23]
  assign _GEN_411 = _T_111 ? vecBools_11 : _GEN_396; // @[Execute.scala 206:23]
  assign _GEN_412 = _T_111 ? vecBools_12 : _GEN_397; // @[Execute.scala 206:23]
  assign _GEN_413 = _T_111 ? vecBools_13 : _GEN_398; // @[Execute.scala 206:23]
  assign _GEN_414 = _T_111 ? vecBools_14 : _GEN_399; // @[Execute.scala 206:23]
  assign _GEN_415 = _T_111 ? vecBools_15 : result[40]; // @[Execute.scala 206:23]
  assign _T_112 = 6'h1a == pos; // @[Execute.scala 206:14]
  assign vecResult_26 = _T_112 ? vecBools_0 : _GEN_401; // @[Execute.scala 206:23]
  assign _GEN_417 = _T_112 ? vecBools_1 : _GEN_402; // @[Execute.scala 206:23]
  assign _GEN_418 = _T_112 ? vecBools_2 : _GEN_403; // @[Execute.scala 206:23]
  assign _GEN_419 = _T_112 ? vecBools_3 : _GEN_404; // @[Execute.scala 206:23]
  assign _GEN_420 = _T_112 ? vecBools_4 : _GEN_405; // @[Execute.scala 206:23]
  assign _GEN_421 = _T_112 ? vecBools_5 : _GEN_406; // @[Execute.scala 206:23]
  assign _GEN_422 = _T_112 ? vecBools_6 : _GEN_407; // @[Execute.scala 206:23]
  assign _GEN_423 = _T_112 ? vecBools_7 : _GEN_408; // @[Execute.scala 206:23]
  assign _GEN_424 = _T_112 ? vecBools_8 : _GEN_409; // @[Execute.scala 206:23]
  assign _GEN_425 = _T_112 ? vecBools_9 : _GEN_410; // @[Execute.scala 206:23]
  assign _GEN_426 = _T_112 ? vecBools_10 : _GEN_411; // @[Execute.scala 206:23]
  assign _GEN_427 = _T_112 ? vecBools_11 : _GEN_412; // @[Execute.scala 206:23]
  assign _GEN_428 = _T_112 ? vecBools_12 : _GEN_413; // @[Execute.scala 206:23]
  assign _GEN_429 = _T_112 ? vecBools_13 : _GEN_414; // @[Execute.scala 206:23]
  assign _GEN_430 = _T_112 ? vecBools_14 : _GEN_415; // @[Execute.scala 206:23]
  assign _GEN_431 = _T_112 ? vecBools_15 : result[41]; // @[Execute.scala 206:23]
  assign _T_113 = 6'h1b == pos; // @[Execute.scala 206:14]
  assign vecResult_27 = _T_113 ? vecBools_0 : _GEN_417; // @[Execute.scala 206:23]
  assign _GEN_433 = _T_113 ? vecBools_1 : _GEN_418; // @[Execute.scala 206:23]
  assign _GEN_434 = _T_113 ? vecBools_2 : _GEN_419; // @[Execute.scala 206:23]
  assign _GEN_435 = _T_113 ? vecBools_3 : _GEN_420; // @[Execute.scala 206:23]
  assign _GEN_436 = _T_113 ? vecBools_4 : _GEN_421; // @[Execute.scala 206:23]
  assign _GEN_437 = _T_113 ? vecBools_5 : _GEN_422; // @[Execute.scala 206:23]
  assign _GEN_438 = _T_113 ? vecBools_6 : _GEN_423; // @[Execute.scala 206:23]
  assign _GEN_439 = _T_113 ? vecBools_7 : _GEN_424; // @[Execute.scala 206:23]
  assign _GEN_440 = _T_113 ? vecBools_8 : _GEN_425; // @[Execute.scala 206:23]
  assign _GEN_441 = _T_113 ? vecBools_9 : _GEN_426; // @[Execute.scala 206:23]
  assign _GEN_442 = _T_113 ? vecBools_10 : _GEN_427; // @[Execute.scala 206:23]
  assign _GEN_443 = _T_113 ? vecBools_11 : _GEN_428; // @[Execute.scala 206:23]
  assign _GEN_444 = _T_113 ? vecBools_12 : _GEN_429; // @[Execute.scala 206:23]
  assign _GEN_445 = _T_113 ? vecBools_13 : _GEN_430; // @[Execute.scala 206:23]
  assign _GEN_446 = _T_113 ? vecBools_14 : _GEN_431; // @[Execute.scala 206:23]
  assign _GEN_447 = _T_113 ? vecBools_15 : result[42]; // @[Execute.scala 206:23]
  assign _T_114 = 6'h1c == pos; // @[Execute.scala 206:14]
  assign vecResult_28 = _T_114 ? vecBools_0 : _GEN_433; // @[Execute.scala 206:23]
  assign _GEN_449 = _T_114 ? vecBools_1 : _GEN_434; // @[Execute.scala 206:23]
  assign _GEN_450 = _T_114 ? vecBools_2 : _GEN_435; // @[Execute.scala 206:23]
  assign _GEN_451 = _T_114 ? vecBools_3 : _GEN_436; // @[Execute.scala 206:23]
  assign _GEN_452 = _T_114 ? vecBools_4 : _GEN_437; // @[Execute.scala 206:23]
  assign _GEN_453 = _T_114 ? vecBools_5 : _GEN_438; // @[Execute.scala 206:23]
  assign _GEN_454 = _T_114 ? vecBools_6 : _GEN_439; // @[Execute.scala 206:23]
  assign _GEN_455 = _T_114 ? vecBools_7 : _GEN_440; // @[Execute.scala 206:23]
  assign _GEN_456 = _T_114 ? vecBools_8 : _GEN_441; // @[Execute.scala 206:23]
  assign _GEN_457 = _T_114 ? vecBools_9 : _GEN_442; // @[Execute.scala 206:23]
  assign _GEN_458 = _T_114 ? vecBools_10 : _GEN_443; // @[Execute.scala 206:23]
  assign _GEN_459 = _T_114 ? vecBools_11 : _GEN_444; // @[Execute.scala 206:23]
  assign _GEN_460 = _T_114 ? vecBools_12 : _GEN_445; // @[Execute.scala 206:23]
  assign _GEN_461 = _T_114 ? vecBools_13 : _GEN_446; // @[Execute.scala 206:23]
  assign _GEN_462 = _T_114 ? vecBools_14 : _GEN_447; // @[Execute.scala 206:23]
  assign _GEN_463 = _T_114 ? vecBools_15 : result[43]; // @[Execute.scala 206:23]
  assign _T_115 = 6'h1d == pos; // @[Execute.scala 206:14]
  assign vecResult_29 = _T_115 ? vecBools_0 : _GEN_449; // @[Execute.scala 206:23]
  assign _GEN_465 = _T_115 ? vecBools_1 : _GEN_450; // @[Execute.scala 206:23]
  assign _GEN_466 = _T_115 ? vecBools_2 : _GEN_451; // @[Execute.scala 206:23]
  assign _GEN_467 = _T_115 ? vecBools_3 : _GEN_452; // @[Execute.scala 206:23]
  assign _GEN_468 = _T_115 ? vecBools_4 : _GEN_453; // @[Execute.scala 206:23]
  assign _GEN_469 = _T_115 ? vecBools_5 : _GEN_454; // @[Execute.scala 206:23]
  assign _GEN_470 = _T_115 ? vecBools_6 : _GEN_455; // @[Execute.scala 206:23]
  assign _GEN_471 = _T_115 ? vecBools_7 : _GEN_456; // @[Execute.scala 206:23]
  assign _GEN_472 = _T_115 ? vecBools_8 : _GEN_457; // @[Execute.scala 206:23]
  assign _GEN_473 = _T_115 ? vecBools_9 : _GEN_458; // @[Execute.scala 206:23]
  assign _GEN_474 = _T_115 ? vecBools_10 : _GEN_459; // @[Execute.scala 206:23]
  assign _GEN_475 = _T_115 ? vecBools_11 : _GEN_460; // @[Execute.scala 206:23]
  assign _GEN_476 = _T_115 ? vecBools_12 : _GEN_461; // @[Execute.scala 206:23]
  assign _GEN_477 = _T_115 ? vecBools_13 : _GEN_462; // @[Execute.scala 206:23]
  assign _GEN_478 = _T_115 ? vecBools_14 : _GEN_463; // @[Execute.scala 206:23]
  assign _GEN_479 = _T_115 ? vecBools_15 : result[44]; // @[Execute.scala 206:23]
  assign _T_116 = 6'h1e == pos; // @[Execute.scala 206:14]
  assign vecResult_30 = _T_116 ? vecBools_0 : _GEN_465; // @[Execute.scala 206:23]
  assign _GEN_481 = _T_116 ? vecBools_1 : _GEN_466; // @[Execute.scala 206:23]
  assign _GEN_482 = _T_116 ? vecBools_2 : _GEN_467; // @[Execute.scala 206:23]
  assign _GEN_483 = _T_116 ? vecBools_3 : _GEN_468; // @[Execute.scala 206:23]
  assign _GEN_484 = _T_116 ? vecBools_4 : _GEN_469; // @[Execute.scala 206:23]
  assign _GEN_485 = _T_116 ? vecBools_5 : _GEN_470; // @[Execute.scala 206:23]
  assign _GEN_486 = _T_116 ? vecBools_6 : _GEN_471; // @[Execute.scala 206:23]
  assign _GEN_487 = _T_116 ? vecBools_7 : _GEN_472; // @[Execute.scala 206:23]
  assign _GEN_488 = _T_116 ? vecBools_8 : _GEN_473; // @[Execute.scala 206:23]
  assign _GEN_489 = _T_116 ? vecBools_9 : _GEN_474; // @[Execute.scala 206:23]
  assign _GEN_490 = _T_116 ? vecBools_10 : _GEN_475; // @[Execute.scala 206:23]
  assign _GEN_491 = _T_116 ? vecBools_11 : _GEN_476; // @[Execute.scala 206:23]
  assign _GEN_492 = _T_116 ? vecBools_12 : _GEN_477; // @[Execute.scala 206:23]
  assign _GEN_493 = _T_116 ? vecBools_13 : _GEN_478; // @[Execute.scala 206:23]
  assign _GEN_494 = _T_116 ? vecBools_14 : _GEN_479; // @[Execute.scala 206:23]
  assign _GEN_495 = _T_116 ? vecBools_15 : result[45]; // @[Execute.scala 206:23]
  assign _T_117 = 6'h1f == pos; // @[Execute.scala 206:14]
  assign vecResult_31 = _T_117 ? vecBools_0 : _GEN_481; // @[Execute.scala 206:23]
  assign _GEN_497 = _T_117 ? vecBools_1 : _GEN_482; // @[Execute.scala 206:23]
  assign _GEN_498 = _T_117 ? vecBools_2 : _GEN_483; // @[Execute.scala 206:23]
  assign _GEN_499 = _T_117 ? vecBools_3 : _GEN_484; // @[Execute.scala 206:23]
  assign _GEN_500 = _T_117 ? vecBools_4 : _GEN_485; // @[Execute.scala 206:23]
  assign _GEN_501 = _T_117 ? vecBools_5 : _GEN_486; // @[Execute.scala 206:23]
  assign _GEN_502 = _T_117 ? vecBools_6 : _GEN_487; // @[Execute.scala 206:23]
  assign _GEN_503 = _T_117 ? vecBools_7 : _GEN_488; // @[Execute.scala 206:23]
  assign _GEN_504 = _T_117 ? vecBools_8 : _GEN_489; // @[Execute.scala 206:23]
  assign _GEN_505 = _T_117 ? vecBools_9 : _GEN_490; // @[Execute.scala 206:23]
  assign _GEN_506 = _T_117 ? vecBools_10 : _GEN_491; // @[Execute.scala 206:23]
  assign _GEN_507 = _T_117 ? vecBools_11 : _GEN_492; // @[Execute.scala 206:23]
  assign _GEN_508 = _T_117 ? vecBools_12 : _GEN_493; // @[Execute.scala 206:23]
  assign _GEN_509 = _T_117 ? vecBools_13 : _GEN_494; // @[Execute.scala 206:23]
  assign _GEN_510 = _T_117 ? vecBools_14 : _GEN_495; // @[Execute.scala 206:23]
  assign _GEN_511 = _T_117 ? vecBools_15 : result[46]; // @[Execute.scala 206:23]
  assign _T_118 = 6'h20 == pos; // @[Execute.scala 206:14]
  assign vecResult_32 = _T_118 ? vecBools_0 : _GEN_497; // @[Execute.scala 206:23]
  assign _GEN_513 = _T_118 ? vecBools_1 : _GEN_498; // @[Execute.scala 206:23]
  assign _GEN_514 = _T_118 ? vecBools_2 : _GEN_499; // @[Execute.scala 206:23]
  assign _GEN_515 = _T_118 ? vecBools_3 : _GEN_500; // @[Execute.scala 206:23]
  assign _GEN_516 = _T_118 ? vecBools_4 : _GEN_501; // @[Execute.scala 206:23]
  assign _GEN_517 = _T_118 ? vecBools_5 : _GEN_502; // @[Execute.scala 206:23]
  assign _GEN_518 = _T_118 ? vecBools_6 : _GEN_503; // @[Execute.scala 206:23]
  assign _GEN_519 = _T_118 ? vecBools_7 : _GEN_504; // @[Execute.scala 206:23]
  assign _GEN_520 = _T_118 ? vecBools_8 : _GEN_505; // @[Execute.scala 206:23]
  assign _GEN_521 = _T_118 ? vecBools_9 : _GEN_506; // @[Execute.scala 206:23]
  assign _GEN_522 = _T_118 ? vecBools_10 : _GEN_507; // @[Execute.scala 206:23]
  assign _GEN_523 = _T_118 ? vecBools_11 : _GEN_508; // @[Execute.scala 206:23]
  assign _GEN_524 = _T_118 ? vecBools_12 : _GEN_509; // @[Execute.scala 206:23]
  assign _GEN_525 = _T_118 ? vecBools_13 : _GEN_510; // @[Execute.scala 206:23]
  assign _GEN_526 = _T_118 ? vecBools_14 : _GEN_511; // @[Execute.scala 206:23]
  assign _GEN_527 = _T_118 ? vecBools_15 : result[47]; // @[Execute.scala 206:23]
  assign _T_119 = 6'h21 == pos; // @[Execute.scala 206:14]
  assign vecResult_33 = _T_119 ? vecBools_0 : _GEN_513; // @[Execute.scala 206:23]
  assign _GEN_529 = _T_119 ? vecBools_1 : _GEN_514; // @[Execute.scala 206:23]
  assign _GEN_530 = _T_119 ? vecBools_2 : _GEN_515; // @[Execute.scala 206:23]
  assign _GEN_531 = _T_119 ? vecBools_3 : _GEN_516; // @[Execute.scala 206:23]
  assign _GEN_532 = _T_119 ? vecBools_4 : _GEN_517; // @[Execute.scala 206:23]
  assign _GEN_533 = _T_119 ? vecBools_5 : _GEN_518; // @[Execute.scala 206:23]
  assign _GEN_534 = _T_119 ? vecBools_6 : _GEN_519; // @[Execute.scala 206:23]
  assign _GEN_535 = _T_119 ? vecBools_7 : _GEN_520; // @[Execute.scala 206:23]
  assign _GEN_536 = _T_119 ? vecBools_8 : _GEN_521; // @[Execute.scala 206:23]
  assign _GEN_537 = _T_119 ? vecBools_9 : _GEN_522; // @[Execute.scala 206:23]
  assign _GEN_538 = _T_119 ? vecBools_10 : _GEN_523; // @[Execute.scala 206:23]
  assign _GEN_539 = _T_119 ? vecBools_11 : _GEN_524; // @[Execute.scala 206:23]
  assign _GEN_540 = _T_119 ? vecBools_12 : _GEN_525; // @[Execute.scala 206:23]
  assign _GEN_541 = _T_119 ? vecBools_13 : _GEN_526; // @[Execute.scala 206:23]
  assign _GEN_542 = _T_119 ? vecBools_14 : _GEN_527; // @[Execute.scala 206:23]
  assign _GEN_543 = _T_119 ? vecBools_15 : result[48]; // @[Execute.scala 206:23]
  assign _T_120 = 6'h22 == pos; // @[Execute.scala 206:14]
  assign vecResult_34 = _T_120 ? vecBools_0 : _GEN_529; // @[Execute.scala 206:23]
  assign _GEN_545 = _T_120 ? vecBools_1 : _GEN_530; // @[Execute.scala 206:23]
  assign _GEN_546 = _T_120 ? vecBools_2 : _GEN_531; // @[Execute.scala 206:23]
  assign _GEN_547 = _T_120 ? vecBools_3 : _GEN_532; // @[Execute.scala 206:23]
  assign _GEN_548 = _T_120 ? vecBools_4 : _GEN_533; // @[Execute.scala 206:23]
  assign _GEN_549 = _T_120 ? vecBools_5 : _GEN_534; // @[Execute.scala 206:23]
  assign _GEN_550 = _T_120 ? vecBools_6 : _GEN_535; // @[Execute.scala 206:23]
  assign _GEN_551 = _T_120 ? vecBools_7 : _GEN_536; // @[Execute.scala 206:23]
  assign _GEN_552 = _T_120 ? vecBools_8 : _GEN_537; // @[Execute.scala 206:23]
  assign _GEN_553 = _T_120 ? vecBools_9 : _GEN_538; // @[Execute.scala 206:23]
  assign _GEN_554 = _T_120 ? vecBools_10 : _GEN_539; // @[Execute.scala 206:23]
  assign _GEN_555 = _T_120 ? vecBools_11 : _GEN_540; // @[Execute.scala 206:23]
  assign _GEN_556 = _T_120 ? vecBools_12 : _GEN_541; // @[Execute.scala 206:23]
  assign _GEN_557 = _T_120 ? vecBools_13 : _GEN_542; // @[Execute.scala 206:23]
  assign _GEN_558 = _T_120 ? vecBools_14 : _GEN_543; // @[Execute.scala 206:23]
  assign _GEN_559 = _T_120 ? vecBools_15 : result[49]; // @[Execute.scala 206:23]
  assign _T_121 = 6'h23 == pos; // @[Execute.scala 206:14]
  assign vecResult_35 = _T_121 ? vecBools_0 : _GEN_545; // @[Execute.scala 206:23]
  assign _GEN_561 = _T_121 ? vecBools_1 : _GEN_546; // @[Execute.scala 206:23]
  assign _GEN_562 = _T_121 ? vecBools_2 : _GEN_547; // @[Execute.scala 206:23]
  assign _GEN_563 = _T_121 ? vecBools_3 : _GEN_548; // @[Execute.scala 206:23]
  assign _GEN_564 = _T_121 ? vecBools_4 : _GEN_549; // @[Execute.scala 206:23]
  assign _GEN_565 = _T_121 ? vecBools_5 : _GEN_550; // @[Execute.scala 206:23]
  assign _GEN_566 = _T_121 ? vecBools_6 : _GEN_551; // @[Execute.scala 206:23]
  assign _GEN_567 = _T_121 ? vecBools_7 : _GEN_552; // @[Execute.scala 206:23]
  assign _GEN_568 = _T_121 ? vecBools_8 : _GEN_553; // @[Execute.scala 206:23]
  assign _GEN_569 = _T_121 ? vecBools_9 : _GEN_554; // @[Execute.scala 206:23]
  assign _GEN_570 = _T_121 ? vecBools_10 : _GEN_555; // @[Execute.scala 206:23]
  assign _GEN_571 = _T_121 ? vecBools_11 : _GEN_556; // @[Execute.scala 206:23]
  assign _GEN_572 = _T_121 ? vecBools_12 : _GEN_557; // @[Execute.scala 206:23]
  assign _GEN_573 = _T_121 ? vecBools_13 : _GEN_558; // @[Execute.scala 206:23]
  assign _GEN_574 = _T_121 ? vecBools_14 : _GEN_559; // @[Execute.scala 206:23]
  assign _GEN_575 = _T_121 ? vecBools_15 : result[50]; // @[Execute.scala 206:23]
  assign _T_122 = 6'h24 == pos; // @[Execute.scala 206:14]
  assign vecResult_36 = _T_122 ? vecBools_0 : _GEN_561; // @[Execute.scala 206:23]
  assign _GEN_577 = _T_122 ? vecBools_1 : _GEN_562; // @[Execute.scala 206:23]
  assign _GEN_578 = _T_122 ? vecBools_2 : _GEN_563; // @[Execute.scala 206:23]
  assign _GEN_579 = _T_122 ? vecBools_3 : _GEN_564; // @[Execute.scala 206:23]
  assign _GEN_580 = _T_122 ? vecBools_4 : _GEN_565; // @[Execute.scala 206:23]
  assign _GEN_581 = _T_122 ? vecBools_5 : _GEN_566; // @[Execute.scala 206:23]
  assign _GEN_582 = _T_122 ? vecBools_6 : _GEN_567; // @[Execute.scala 206:23]
  assign _GEN_583 = _T_122 ? vecBools_7 : _GEN_568; // @[Execute.scala 206:23]
  assign _GEN_584 = _T_122 ? vecBools_8 : _GEN_569; // @[Execute.scala 206:23]
  assign _GEN_585 = _T_122 ? vecBools_9 : _GEN_570; // @[Execute.scala 206:23]
  assign _GEN_586 = _T_122 ? vecBools_10 : _GEN_571; // @[Execute.scala 206:23]
  assign _GEN_587 = _T_122 ? vecBools_11 : _GEN_572; // @[Execute.scala 206:23]
  assign _GEN_588 = _T_122 ? vecBools_12 : _GEN_573; // @[Execute.scala 206:23]
  assign _GEN_589 = _T_122 ? vecBools_13 : _GEN_574; // @[Execute.scala 206:23]
  assign _GEN_590 = _T_122 ? vecBools_14 : _GEN_575; // @[Execute.scala 206:23]
  assign _GEN_591 = _T_122 ? vecBools_15 : result[51]; // @[Execute.scala 206:23]
  assign _T_123 = 6'h25 == pos; // @[Execute.scala 206:14]
  assign vecResult_37 = _T_123 ? vecBools_0 : _GEN_577; // @[Execute.scala 206:23]
  assign _GEN_593 = _T_123 ? vecBools_1 : _GEN_578; // @[Execute.scala 206:23]
  assign _GEN_594 = _T_123 ? vecBools_2 : _GEN_579; // @[Execute.scala 206:23]
  assign _GEN_595 = _T_123 ? vecBools_3 : _GEN_580; // @[Execute.scala 206:23]
  assign _GEN_596 = _T_123 ? vecBools_4 : _GEN_581; // @[Execute.scala 206:23]
  assign _GEN_597 = _T_123 ? vecBools_5 : _GEN_582; // @[Execute.scala 206:23]
  assign _GEN_598 = _T_123 ? vecBools_6 : _GEN_583; // @[Execute.scala 206:23]
  assign _GEN_599 = _T_123 ? vecBools_7 : _GEN_584; // @[Execute.scala 206:23]
  assign _GEN_600 = _T_123 ? vecBools_8 : _GEN_585; // @[Execute.scala 206:23]
  assign _GEN_601 = _T_123 ? vecBools_9 : _GEN_586; // @[Execute.scala 206:23]
  assign _GEN_602 = _T_123 ? vecBools_10 : _GEN_587; // @[Execute.scala 206:23]
  assign _GEN_603 = _T_123 ? vecBools_11 : _GEN_588; // @[Execute.scala 206:23]
  assign _GEN_604 = _T_123 ? vecBools_12 : _GEN_589; // @[Execute.scala 206:23]
  assign _GEN_605 = _T_123 ? vecBools_13 : _GEN_590; // @[Execute.scala 206:23]
  assign _GEN_606 = _T_123 ? vecBools_14 : _GEN_591; // @[Execute.scala 206:23]
  assign _GEN_607 = _T_123 ? vecBools_15 : result[52]; // @[Execute.scala 206:23]
  assign _T_124 = 6'h26 == pos; // @[Execute.scala 206:14]
  assign vecResult_38 = _T_124 ? vecBools_0 : _GEN_593; // @[Execute.scala 206:23]
  assign _GEN_609 = _T_124 ? vecBools_1 : _GEN_594; // @[Execute.scala 206:23]
  assign _GEN_610 = _T_124 ? vecBools_2 : _GEN_595; // @[Execute.scala 206:23]
  assign _GEN_611 = _T_124 ? vecBools_3 : _GEN_596; // @[Execute.scala 206:23]
  assign _GEN_612 = _T_124 ? vecBools_4 : _GEN_597; // @[Execute.scala 206:23]
  assign _GEN_613 = _T_124 ? vecBools_5 : _GEN_598; // @[Execute.scala 206:23]
  assign _GEN_614 = _T_124 ? vecBools_6 : _GEN_599; // @[Execute.scala 206:23]
  assign _GEN_615 = _T_124 ? vecBools_7 : _GEN_600; // @[Execute.scala 206:23]
  assign _GEN_616 = _T_124 ? vecBools_8 : _GEN_601; // @[Execute.scala 206:23]
  assign _GEN_617 = _T_124 ? vecBools_9 : _GEN_602; // @[Execute.scala 206:23]
  assign _GEN_618 = _T_124 ? vecBools_10 : _GEN_603; // @[Execute.scala 206:23]
  assign _GEN_619 = _T_124 ? vecBools_11 : _GEN_604; // @[Execute.scala 206:23]
  assign _GEN_620 = _T_124 ? vecBools_12 : _GEN_605; // @[Execute.scala 206:23]
  assign _GEN_621 = _T_124 ? vecBools_13 : _GEN_606; // @[Execute.scala 206:23]
  assign _GEN_622 = _T_124 ? vecBools_14 : _GEN_607; // @[Execute.scala 206:23]
  assign _GEN_623 = _T_124 ? vecBools_15 : result[53]; // @[Execute.scala 206:23]
  assign _T_125 = 6'h27 == pos; // @[Execute.scala 206:14]
  assign vecResult_39 = _T_125 ? vecBools_0 : _GEN_609; // @[Execute.scala 206:23]
  assign _GEN_625 = _T_125 ? vecBools_1 : _GEN_610; // @[Execute.scala 206:23]
  assign _GEN_626 = _T_125 ? vecBools_2 : _GEN_611; // @[Execute.scala 206:23]
  assign _GEN_627 = _T_125 ? vecBools_3 : _GEN_612; // @[Execute.scala 206:23]
  assign _GEN_628 = _T_125 ? vecBools_4 : _GEN_613; // @[Execute.scala 206:23]
  assign _GEN_629 = _T_125 ? vecBools_5 : _GEN_614; // @[Execute.scala 206:23]
  assign _GEN_630 = _T_125 ? vecBools_6 : _GEN_615; // @[Execute.scala 206:23]
  assign _GEN_631 = _T_125 ? vecBools_7 : _GEN_616; // @[Execute.scala 206:23]
  assign _GEN_632 = _T_125 ? vecBools_8 : _GEN_617; // @[Execute.scala 206:23]
  assign _GEN_633 = _T_125 ? vecBools_9 : _GEN_618; // @[Execute.scala 206:23]
  assign _GEN_634 = _T_125 ? vecBools_10 : _GEN_619; // @[Execute.scala 206:23]
  assign _GEN_635 = _T_125 ? vecBools_11 : _GEN_620; // @[Execute.scala 206:23]
  assign _GEN_636 = _T_125 ? vecBools_12 : _GEN_621; // @[Execute.scala 206:23]
  assign _GEN_637 = _T_125 ? vecBools_13 : _GEN_622; // @[Execute.scala 206:23]
  assign _GEN_638 = _T_125 ? vecBools_14 : _GEN_623; // @[Execute.scala 206:23]
  assign _GEN_639 = _T_125 ? vecBools_15 : result[54]; // @[Execute.scala 206:23]
  assign _T_126 = 6'h28 == pos; // @[Execute.scala 206:14]
  assign vecResult_40 = _T_126 ? vecBools_0 : _GEN_625; // @[Execute.scala 206:23]
  assign _GEN_641 = _T_126 ? vecBools_1 : _GEN_626; // @[Execute.scala 206:23]
  assign _GEN_642 = _T_126 ? vecBools_2 : _GEN_627; // @[Execute.scala 206:23]
  assign _GEN_643 = _T_126 ? vecBools_3 : _GEN_628; // @[Execute.scala 206:23]
  assign _GEN_644 = _T_126 ? vecBools_4 : _GEN_629; // @[Execute.scala 206:23]
  assign _GEN_645 = _T_126 ? vecBools_5 : _GEN_630; // @[Execute.scala 206:23]
  assign _GEN_646 = _T_126 ? vecBools_6 : _GEN_631; // @[Execute.scala 206:23]
  assign _GEN_647 = _T_126 ? vecBools_7 : _GEN_632; // @[Execute.scala 206:23]
  assign _GEN_648 = _T_126 ? vecBools_8 : _GEN_633; // @[Execute.scala 206:23]
  assign _GEN_649 = _T_126 ? vecBools_9 : _GEN_634; // @[Execute.scala 206:23]
  assign _GEN_650 = _T_126 ? vecBools_10 : _GEN_635; // @[Execute.scala 206:23]
  assign _GEN_651 = _T_126 ? vecBools_11 : _GEN_636; // @[Execute.scala 206:23]
  assign _GEN_652 = _T_126 ? vecBools_12 : _GEN_637; // @[Execute.scala 206:23]
  assign _GEN_653 = _T_126 ? vecBools_13 : _GEN_638; // @[Execute.scala 206:23]
  assign _GEN_654 = _T_126 ? vecBools_14 : _GEN_639; // @[Execute.scala 206:23]
  assign _GEN_655 = _T_126 ? vecBools_15 : result[55]; // @[Execute.scala 206:23]
  assign _T_127 = 6'h29 == pos; // @[Execute.scala 206:14]
  assign vecResult_41 = _T_127 ? vecBools_0 : _GEN_641; // @[Execute.scala 206:23]
  assign _GEN_657 = _T_127 ? vecBools_1 : _GEN_642; // @[Execute.scala 206:23]
  assign _GEN_658 = _T_127 ? vecBools_2 : _GEN_643; // @[Execute.scala 206:23]
  assign _GEN_659 = _T_127 ? vecBools_3 : _GEN_644; // @[Execute.scala 206:23]
  assign _GEN_660 = _T_127 ? vecBools_4 : _GEN_645; // @[Execute.scala 206:23]
  assign _GEN_661 = _T_127 ? vecBools_5 : _GEN_646; // @[Execute.scala 206:23]
  assign _GEN_662 = _T_127 ? vecBools_6 : _GEN_647; // @[Execute.scala 206:23]
  assign _GEN_663 = _T_127 ? vecBools_7 : _GEN_648; // @[Execute.scala 206:23]
  assign _GEN_664 = _T_127 ? vecBools_8 : _GEN_649; // @[Execute.scala 206:23]
  assign _GEN_665 = _T_127 ? vecBools_9 : _GEN_650; // @[Execute.scala 206:23]
  assign _GEN_666 = _T_127 ? vecBools_10 : _GEN_651; // @[Execute.scala 206:23]
  assign _GEN_667 = _T_127 ? vecBools_11 : _GEN_652; // @[Execute.scala 206:23]
  assign _GEN_668 = _T_127 ? vecBools_12 : _GEN_653; // @[Execute.scala 206:23]
  assign _GEN_669 = _T_127 ? vecBools_13 : _GEN_654; // @[Execute.scala 206:23]
  assign _GEN_670 = _T_127 ? vecBools_14 : _GEN_655; // @[Execute.scala 206:23]
  assign _GEN_671 = _T_127 ? vecBools_15 : result[56]; // @[Execute.scala 206:23]
  assign _T_128 = 6'h2a == pos; // @[Execute.scala 206:14]
  assign vecResult_42 = _T_128 ? vecBools_0 : _GEN_657; // @[Execute.scala 206:23]
  assign _GEN_673 = _T_128 ? vecBools_1 : _GEN_658; // @[Execute.scala 206:23]
  assign _GEN_674 = _T_128 ? vecBools_2 : _GEN_659; // @[Execute.scala 206:23]
  assign _GEN_675 = _T_128 ? vecBools_3 : _GEN_660; // @[Execute.scala 206:23]
  assign _GEN_676 = _T_128 ? vecBools_4 : _GEN_661; // @[Execute.scala 206:23]
  assign _GEN_677 = _T_128 ? vecBools_5 : _GEN_662; // @[Execute.scala 206:23]
  assign _GEN_678 = _T_128 ? vecBools_6 : _GEN_663; // @[Execute.scala 206:23]
  assign _GEN_679 = _T_128 ? vecBools_7 : _GEN_664; // @[Execute.scala 206:23]
  assign _GEN_680 = _T_128 ? vecBools_8 : _GEN_665; // @[Execute.scala 206:23]
  assign _GEN_681 = _T_128 ? vecBools_9 : _GEN_666; // @[Execute.scala 206:23]
  assign _GEN_682 = _T_128 ? vecBools_10 : _GEN_667; // @[Execute.scala 206:23]
  assign _GEN_683 = _T_128 ? vecBools_11 : _GEN_668; // @[Execute.scala 206:23]
  assign _GEN_684 = _T_128 ? vecBools_12 : _GEN_669; // @[Execute.scala 206:23]
  assign _GEN_685 = _T_128 ? vecBools_13 : _GEN_670; // @[Execute.scala 206:23]
  assign _GEN_686 = _T_128 ? vecBools_14 : _GEN_671; // @[Execute.scala 206:23]
  assign _GEN_687 = _T_128 ? vecBools_15 : result[57]; // @[Execute.scala 206:23]
  assign _T_129 = 6'h2b == pos; // @[Execute.scala 206:14]
  assign vecResult_43 = _T_129 ? vecBools_0 : _GEN_673; // @[Execute.scala 206:23]
  assign _GEN_689 = _T_129 ? vecBools_1 : _GEN_674; // @[Execute.scala 206:23]
  assign _GEN_690 = _T_129 ? vecBools_2 : _GEN_675; // @[Execute.scala 206:23]
  assign _GEN_691 = _T_129 ? vecBools_3 : _GEN_676; // @[Execute.scala 206:23]
  assign _GEN_692 = _T_129 ? vecBools_4 : _GEN_677; // @[Execute.scala 206:23]
  assign _GEN_693 = _T_129 ? vecBools_5 : _GEN_678; // @[Execute.scala 206:23]
  assign _GEN_694 = _T_129 ? vecBools_6 : _GEN_679; // @[Execute.scala 206:23]
  assign _GEN_695 = _T_129 ? vecBools_7 : _GEN_680; // @[Execute.scala 206:23]
  assign _GEN_696 = _T_129 ? vecBools_8 : _GEN_681; // @[Execute.scala 206:23]
  assign _GEN_697 = _T_129 ? vecBools_9 : _GEN_682; // @[Execute.scala 206:23]
  assign _GEN_698 = _T_129 ? vecBools_10 : _GEN_683; // @[Execute.scala 206:23]
  assign _GEN_699 = _T_129 ? vecBools_11 : _GEN_684; // @[Execute.scala 206:23]
  assign _GEN_700 = _T_129 ? vecBools_12 : _GEN_685; // @[Execute.scala 206:23]
  assign _GEN_701 = _T_129 ? vecBools_13 : _GEN_686; // @[Execute.scala 206:23]
  assign _GEN_702 = _T_129 ? vecBools_14 : _GEN_687; // @[Execute.scala 206:23]
  assign _GEN_703 = _T_129 ? vecBools_15 : result[58]; // @[Execute.scala 206:23]
  assign _T_130 = 6'h2c == pos; // @[Execute.scala 206:14]
  assign vecResult_44 = _T_130 ? vecBools_0 : _GEN_689; // @[Execute.scala 206:23]
  assign _GEN_705 = _T_130 ? vecBools_1 : _GEN_690; // @[Execute.scala 206:23]
  assign _GEN_706 = _T_130 ? vecBools_2 : _GEN_691; // @[Execute.scala 206:23]
  assign _GEN_707 = _T_130 ? vecBools_3 : _GEN_692; // @[Execute.scala 206:23]
  assign _GEN_708 = _T_130 ? vecBools_4 : _GEN_693; // @[Execute.scala 206:23]
  assign _GEN_709 = _T_130 ? vecBools_5 : _GEN_694; // @[Execute.scala 206:23]
  assign _GEN_710 = _T_130 ? vecBools_6 : _GEN_695; // @[Execute.scala 206:23]
  assign _GEN_711 = _T_130 ? vecBools_7 : _GEN_696; // @[Execute.scala 206:23]
  assign _GEN_712 = _T_130 ? vecBools_8 : _GEN_697; // @[Execute.scala 206:23]
  assign _GEN_713 = _T_130 ? vecBools_9 : _GEN_698; // @[Execute.scala 206:23]
  assign _GEN_714 = _T_130 ? vecBools_10 : _GEN_699; // @[Execute.scala 206:23]
  assign _GEN_715 = _T_130 ? vecBools_11 : _GEN_700; // @[Execute.scala 206:23]
  assign _GEN_716 = _T_130 ? vecBools_12 : _GEN_701; // @[Execute.scala 206:23]
  assign _GEN_717 = _T_130 ? vecBools_13 : _GEN_702; // @[Execute.scala 206:23]
  assign _GEN_718 = _T_130 ? vecBools_14 : _GEN_703; // @[Execute.scala 206:23]
  assign _GEN_719 = _T_130 ? vecBools_15 : result[59]; // @[Execute.scala 206:23]
  assign _T_131 = 6'h2d == pos; // @[Execute.scala 206:14]
  assign vecResult_45 = _T_131 ? vecBools_0 : _GEN_705; // @[Execute.scala 206:23]
  assign _GEN_721 = _T_131 ? vecBools_1 : _GEN_706; // @[Execute.scala 206:23]
  assign _GEN_722 = _T_131 ? vecBools_2 : _GEN_707; // @[Execute.scala 206:23]
  assign _GEN_723 = _T_131 ? vecBools_3 : _GEN_708; // @[Execute.scala 206:23]
  assign _GEN_724 = _T_131 ? vecBools_4 : _GEN_709; // @[Execute.scala 206:23]
  assign _GEN_725 = _T_131 ? vecBools_5 : _GEN_710; // @[Execute.scala 206:23]
  assign _GEN_726 = _T_131 ? vecBools_6 : _GEN_711; // @[Execute.scala 206:23]
  assign _GEN_727 = _T_131 ? vecBools_7 : _GEN_712; // @[Execute.scala 206:23]
  assign _GEN_728 = _T_131 ? vecBools_8 : _GEN_713; // @[Execute.scala 206:23]
  assign _GEN_729 = _T_131 ? vecBools_9 : _GEN_714; // @[Execute.scala 206:23]
  assign _GEN_730 = _T_131 ? vecBools_10 : _GEN_715; // @[Execute.scala 206:23]
  assign _GEN_731 = _T_131 ? vecBools_11 : _GEN_716; // @[Execute.scala 206:23]
  assign _GEN_732 = _T_131 ? vecBools_12 : _GEN_717; // @[Execute.scala 206:23]
  assign _GEN_733 = _T_131 ? vecBools_13 : _GEN_718; // @[Execute.scala 206:23]
  assign _GEN_734 = _T_131 ? vecBools_14 : _GEN_719; // @[Execute.scala 206:23]
  assign _GEN_735 = _T_131 ? vecBools_15 : result[60]; // @[Execute.scala 206:23]
  assign _T_132 = 6'h2e == pos; // @[Execute.scala 206:14]
  assign vecResult_46 = _T_132 ? vecBools_0 : _GEN_721; // @[Execute.scala 206:23]
  assign _GEN_737 = _T_132 ? vecBools_1 : _GEN_722; // @[Execute.scala 206:23]
  assign _GEN_738 = _T_132 ? vecBools_2 : _GEN_723; // @[Execute.scala 206:23]
  assign _GEN_739 = _T_132 ? vecBools_3 : _GEN_724; // @[Execute.scala 206:23]
  assign _GEN_740 = _T_132 ? vecBools_4 : _GEN_725; // @[Execute.scala 206:23]
  assign _GEN_741 = _T_132 ? vecBools_5 : _GEN_726; // @[Execute.scala 206:23]
  assign _GEN_742 = _T_132 ? vecBools_6 : _GEN_727; // @[Execute.scala 206:23]
  assign _GEN_743 = _T_132 ? vecBools_7 : _GEN_728; // @[Execute.scala 206:23]
  assign _GEN_744 = _T_132 ? vecBools_8 : _GEN_729; // @[Execute.scala 206:23]
  assign _GEN_745 = _T_132 ? vecBools_9 : _GEN_730; // @[Execute.scala 206:23]
  assign _GEN_746 = _T_132 ? vecBools_10 : _GEN_731; // @[Execute.scala 206:23]
  assign _GEN_747 = _T_132 ? vecBools_11 : _GEN_732; // @[Execute.scala 206:23]
  assign _GEN_748 = _T_132 ? vecBools_12 : _GEN_733; // @[Execute.scala 206:23]
  assign _GEN_749 = _T_132 ? vecBools_13 : _GEN_734; // @[Execute.scala 206:23]
  assign _GEN_750 = _T_132 ? vecBools_14 : _GEN_735; // @[Execute.scala 206:23]
  assign _GEN_751 = _T_132 ? vecBools_15 : result[61]; // @[Execute.scala 206:23]
  assign _T_133 = 6'h2f == pos; // @[Execute.scala 206:14]
  assign vecResult_47 = _T_133 ? vecBools_0 : _GEN_737; // @[Execute.scala 206:23]
  assign _GEN_753 = _T_133 ? vecBools_1 : _GEN_738; // @[Execute.scala 206:23]
  assign _GEN_754 = _T_133 ? vecBools_2 : _GEN_739; // @[Execute.scala 206:23]
  assign _GEN_755 = _T_133 ? vecBools_3 : _GEN_740; // @[Execute.scala 206:23]
  assign _GEN_756 = _T_133 ? vecBools_4 : _GEN_741; // @[Execute.scala 206:23]
  assign _GEN_757 = _T_133 ? vecBools_5 : _GEN_742; // @[Execute.scala 206:23]
  assign _GEN_758 = _T_133 ? vecBools_6 : _GEN_743; // @[Execute.scala 206:23]
  assign _GEN_759 = _T_133 ? vecBools_7 : _GEN_744; // @[Execute.scala 206:23]
  assign _GEN_760 = _T_133 ? vecBools_8 : _GEN_745; // @[Execute.scala 206:23]
  assign _GEN_761 = _T_133 ? vecBools_9 : _GEN_746; // @[Execute.scala 206:23]
  assign _GEN_762 = _T_133 ? vecBools_10 : _GEN_747; // @[Execute.scala 206:23]
  assign _GEN_763 = _T_133 ? vecBools_11 : _GEN_748; // @[Execute.scala 206:23]
  assign _GEN_764 = _T_133 ? vecBools_12 : _GEN_749; // @[Execute.scala 206:23]
  assign _GEN_765 = _T_133 ? vecBools_13 : _GEN_750; // @[Execute.scala 206:23]
  assign _GEN_766 = _T_133 ? vecBools_14 : _GEN_751; // @[Execute.scala 206:23]
  assign _GEN_767 = _T_133 ? vecBools_15 : result[62]; // @[Execute.scala 206:23]
  assign _T_134 = 6'h30 == pos; // @[Execute.scala 206:14]
  assign vecResult_48 = _T_134 ? vecBools_0 : _GEN_753; // @[Execute.scala 206:23]
  assign vecResult_49 = _T_134 ? vecBools_1 : _GEN_754; // @[Execute.scala 206:23]
  assign vecResult_50 = _T_134 ? vecBools_2 : _GEN_755; // @[Execute.scala 206:23]
  assign vecResult_51 = _T_134 ? vecBools_3 : _GEN_756; // @[Execute.scala 206:23]
  assign vecResult_52 = _T_134 ? vecBools_4 : _GEN_757; // @[Execute.scala 206:23]
  assign vecResult_53 = _T_134 ? vecBools_5 : _GEN_758; // @[Execute.scala 206:23]
  assign vecResult_54 = _T_134 ? vecBools_6 : _GEN_759; // @[Execute.scala 206:23]
  assign vecResult_55 = _T_134 ? vecBools_7 : _GEN_760; // @[Execute.scala 206:23]
  assign vecResult_56 = _T_134 ? vecBools_8 : _GEN_761; // @[Execute.scala 206:23]
  assign vecResult_57 = _T_134 ? vecBools_9 : _GEN_762; // @[Execute.scala 206:23]
  assign vecResult_58 = _T_134 ? vecBools_10 : _GEN_763; // @[Execute.scala 206:23]
  assign vecResult_59 = _T_134 ? vecBools_11 : _GEN_764; // @[Execute.scala 206:23]
  assign vecResult_60 = _T_134 ? vecBools_12 : _GEN_765; // @[Execute.scala 206:23]
  assign vecResult_61 = _T_134 ? vecBools_13 : _GEN_766; // @[Execute.scala 206:23]
  assign vecResult_62 = _T_134 ? vecBools_14 : _GEN_767; // @[Execute.scala 206:23]
  assign vecResult_63 = _T_134 ? vecBools_15 : result[63]; // @[Execute.scala 206:23]
  assign _T_141 = {vecResult_7,vecResult_6,vecResult_5,vecResult_4,vecResult_3,vecResult_2,vecResult_1,vecResult_0}; // @[Execute.scala 213:32]
  assign _T_149 = {vecResult_15,vecResult_14,vecResult_13,vecResult_12,vecResult_11,vecResult_10,vecResult_9,vecResult_8,_T_141}; // @[Execute.scala 213:32]
  assign _T_156 = {vecResult_23,vecResult_22,vecResult_21,vecResult_20,vecResult_19,vecResult_18,vecResult_17,vecResult_16}; // @[Execute.scala 213:32]
  assign _T_165 = {vecResult_31,vecResult_30,vecResult_29,vecResult_28,vecResult_27,vecResult_26,vecResult_25,vecResult_24,_T_156,_T_149}; // @[Execute.scala 213:32]
  assign _T_172 = {vecResult_39,vecResult_38,vecResult_37,vecResult_36,vecResult_35,vecResult_34,vecResult_33,vecResult_32}; // @[Execute.scala 213:32]
  assign _T_180 = {vecResult_47,vecResult_46,vecResult_45,vecResult_44,vecResult_43,vecResult_42,vecResult_41,vecResult_40,_T_172}; // @[Execute.scala 213:32]
  assign _T_187 = {vecResult_55,vecResult_54,vecResult_53,vecResult_52,vecResult_51,vecResult_50,vecResult_49,vecResult_48}; // @[Execute.scala 213:32]
  assign _T_196 = {vecResult_63,vecResult_62,vecResult_61,vecResult_60,vecResult_59,vecResult_58,vecResult_57,vecResult_56,_T_187,_T_180}; // @[Execute.scala 213:32]
  assign res = {_T_196,_T_165}; // @[Execute.scala 213:32]
  assign _T_198 = io_op == 4'h0; // @[Execute.scala 214:23]
  assign _T_199 = ~res; // @[Execute.scala 214:36]
  assign io_res = _T_198 ? _T_199 : res; // @[Execute.scala 214:10]
endmodule
