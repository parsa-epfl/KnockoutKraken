module DataAlignByte(
  input         io_currReq,
  input  [1:0]  io_minst_size,
  input         io_minst_isPair,
  input         io_minst_isLoad,
  input  [63:0] io_minst_memReq_0_addr,
  input  [63:0] io_minst_memReq_1_addr,
  input  [63:0] io_data,
  output [63:0] io_aligned,
  output [7:0]  io_byteEn,
  output        io_unalignedExcp
);
  wire [7:0] dataBytes_0; // @[LoadStore.scala 273:50]
  wire [7:0] dataBytes_1; // @[LoadStore.scala 273:50]
  wire [7:0] dataBytes_2; // @[LoadStore.scala 273:50]
  wire [7:0] dataBytes_3; // @[LoadStore.scala 273:50]
  wire [7:0] dataBytes_4; // @[LoadStore.scala 273:50]
  wire [7:0] dataBytes_5; // @[LoadStore.scala 273:50]
  wire [7:0] dataBytes_6; // @[LoadStore.scala 273:50]
  wire [7:0] dataBytes_7; // @[LoadStore.scala 273:50]
  wire [63:0] _GEN_3; // @[LoadStore.scala 280:29]
  wire [2:0] _T_11; // @[LoadStore.scala 281:39]
  wire [7:0] _GEN_7; // @[Cat.scala 29:58]
  wire [7:0] _GEN_8; // @[Cat.scala 29:58]
  wire [7:0] _GEN_9; // @[Cat.scala 29:58]
  wire [7:0] _GEN_10; // @[Cat.scala 29:58]
  wire [7:0] _GEN_11; // @[Cat.scala 29:58]
  wire [7:0] _GEN_12; // @[Cat.scala 29:58]
  wire [7:0] _GEN_13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_15; // @[Cat.scala 29:58]
  wire [7:0] _GEN_16; // @[Cat.scala 29:58]
  wire [7:0] _GEN_17; // @[Cat.scala 29:58]
  wire [7:0] _GEN_18; // @[Cat.scala 29:58]
  wire [7:0] _GEN_19; // @[Cat.scala 29:58]
  wire [7:0] _GEN_20; // @[Cat.scala 29:58]
  wire [7:0] _GEN_21; // @[Cat.scala 29:58]
  wire [15:0] _T_13; // @[Cat.scala 29:58]
  wire [31:0] _T_17; // @[LoadStore.scala 282:18]
  wire  _T_18; // @[Mux.scala 80:60]
  wire [15:0] _T_19; // @[Mux.scala 80:57]
  wire  _T_20; // @[Mux.scala 80:60]
  wire [31:0] _T_21; // @[Mux.scala 80:57]
  wire  _T_22; // @[Mux.scala 80:60]
  wire [63:0] data2align; // @[Mux.scala 80:57]
  wire [5:0] _T_72; // @[Cat.scala 29:58]
  wire [126:0] _GEN_30; // @[LoadStore.scala 310:38]
  wire [126:0] byteAlignStore; // @[LoadStore.scala 310:38]
  wire [1:0] _T_75; // @[Mux.scala 80:57]
  wire [3:0] _T_77; // @[Mux.scala 80:57]
  wire [7:0] mask; // @[Mux.scala 80:57]
  wire [14:0] _GEN_31; // @[LoadStore.scala 320:30]
  wire [14:0] byteEn; // @[LoadStore.scala 320:30]
  wire  _T_83; // @[LoadStore.scala 325:40]
  wire  _T_85; // @[LoadStore.scala 326:42]
  wire  _T_87; // @[LoadStore.scala 327:42]
  wire  _T_89; // @[Mux.scala 80:57]
  wire  _T_91; // @[Mux.scala 80:57]
  wire  isAlignedMem_0; // @[Mux.scala 80:57]
  wire  _T_95; // @[LoadStore.scala 332:40]
  wire  _T_97; // @[LoadStore.scala 333:42]
  wire  _T_99; // @[LoadStore.scala 334:42]
  wire  _T_101; // @[Mux.scala 80:57]
  wire  _T_103; // @[Mux.scala 80:57]
  wire  isAlignedMem_1; // @[Mux.scala 80:57]
  wire [14:0] _T_106; // @[LoadStore.scala 338:19]
  wire [126:0] _T_107; // @[LoadStore.scala 339:20]
  wire  _T_108; // @[LoadStore.scala 341:23]
  wire  _T_109; // @[LoadStore.scala 341:59]
  wire  _T_110; // @[LoadStore.scala 341:56]
  assign dataBytes_0 = io_data[7:0]; // @[LoadStore.scala 273:50]
  assign dataBytes_1 = io_data[15:8]; // @[LoadStore.scala 273:50]
  assign dataBytes_2 = io_data[23:16]; // @[LoadStore.scala 273:50]
  assign dataBytes_3 = io_data[31:24]; // @[LoadStore.scala 273:50]
  assign dataBytes_4 = io_data[39:32]; // @[LoadStore.scala 273:50]
  assign dataBytes_5 = io_data[47:40]; // @[LoadStore.scala 273:50]
  assign dataBytes_6 = io_data[55:48]; // @[LoadStore.scala 273:50]
  assign dataBytes_7 = io_data[63:56]; // @[LoadStore.scala 273:50]
  assign _GEN_3 = io_currReq ? io_minst_memReq_1_addr : io_minst_memReq_0_addr; // @[LoadStore.scala 280:29]
  assign _T_11 = _GEN_3[2:0] + 3'h1; // @[LoadStore.scala 281:39]
  assign _GEN_7 = 3'h1 == _T_11 ? dataBytes_1 : dataBytes_0; // @[Cat.scala 29:58]
  assign _GEN_8 = 3'h2 == _T_11 ? dataBytes_2 : _GEN_7; // @[Cat.scala 29:58]
  assign _GEN_9 = 3'h3 == _T_11 ? dataBytes_3 : _GEN_8; // @[Cat.scala 29:58]
  assign _GEN_10 = 3'h4 == _T_11 ? dataBytes_4 : _GEN_9; // @[Cat.scala 29:58]
  assign _GEN_11 = 3'h5 == _T_11 ? dataBytes_5 : _GEN_10; // @[Cat.scala 29:58]
  assign _GEN_12 = 3'h6 == _T_11 ? dataBytes_6 : _GEN_11; // @[Cat.scala 29:58]
  assign _GEN_13 = 3'h7 == _T_11 ? dataBytes_7 : _GEN_12; // @[Cat.scala 29:58]
  assign _GEN_15 = 3'h1 == _GEN_3[2:0] ? dataBytes_1 : dataBytes_0; // @[Cat.scala 29:58]
  assign _GEN_16 = 3'h2 == _GEN_3[2:0] ? dataBytes_2 : _GEN_15; // @[Cat.scala 29:58]
  assign _GEN_17 = 3'h3 == _GEN_3[2:0] ? dataBytes_3 : _GEN_16; // @[Cat.scala 29:58]
  assign _GEN_18 = 3'h4 == _GEN_3[2:0] ? dataBytes_4 : _GEN_17; // @[Cat.scala 29:58]
  assign _GEN_19 = 3'h5 == _GEN_3[2:0] ? dataBytes_5 : _GEN_18; // @[Cat.scala 29:58]
  assign _GEN_20 = 3'h6 == _GEN_3[2:0] ? dataBytes_6 : _GEN_19; // @[Cat.scala 29:58]
  assign _GEN_21 = 3'h7 == _GEN_3[2:0] ? dataBytes_7 : _GEN_20; // @[Cat.scala 29:58]
  assign _T_13 = {_GEN_13,_GEN_21}; // @[Cat.scala 29:58]
  assign _T_17 = _GEN_3[2] ? io_data[63:32] : io_data[31:0]; // @[LoadStore.scala 282:18]
  assign _T_18 = 2'h1 == io_minst_size; // @[Mux.scala 80:60]
  assign _T_19 = _T_18 ? _T_13 : {{8'd0}, _GEN_21}; // @[Mux.scala 80:57]
  assign _T_20 = 2'h2 == io_minst_size; // @[Mux.scala 80:60]
  assign _T_21 = _T_20 ? _T_17 : {{16'd0}, _T_19}; // @[Mux.scala 80:57]
  assign _T_22 = 2'h3 == io_minst_size; // @[Mux.scala 80:60]
  assign data2align = _T_22 ? io_data : {{32'd0}, _T_21}; // @[Mux.scala 80:57]
  assign _T_72 = {_GEN_3[2:0],3'h0}; // @[Cat.scala 29:58]
  assign _GEN_30 = {{63'd0}, io_data}; // @[LoadStore.scala 310:38]
  assign byteAlignStore = _GEN_30 << _T_72; // @[LoadStore.scala 310:38]
  assign _T_75 = _T_18 ? 2'h3 : 2'h1; // @[Mux.scala 80:57]
  assign _T_77 = _T_20 ? 4'hf : {{2'd0}, _T_75}; // @[Mux.scala 80:57]
  assign mask = _T_22 ? 8'hff : {{4'd0}, _T_77}; // @[Mux.scala 80:57]
  assign _GEN_31 = {{7'd0}, mask}; // @[LoadStore.scala 320:30]
  assign byteEn = _GEN_31 << _GEN_3[2:0]; // @[LoadStore.scala 320:30]
  assign _T_83 = ~io_minst_memReq_0_addr[0]; // @[LoadStore.scala 325:40]
  assign _T_85 = io_minst_memReq_0_addr[1:0] == 2'h0; // @[LoadStore.scala 326:42]
  assign _T_87 = io_minst_memReq_0_addr[2:0] == 3'h0; // @[LoadStore.scala 327:42]
  assign _T_89 = _T_18 ? _T_83 : 1'h1; // @[Mux.scala 80:57]
  assign _T_91 = _T_20 ? _T_85 : _T_89; // @[Mux.scala 80:57]
  assign isAlignedMem_0 = _T_22 ? _T_87 : _T_91; // @[Mux.scala 80:57]
  assign _T_95 = ~io_minst_memReq_1_addr[0]; // @[LoadStore.scala 332:40]
  assign _T_97 = io_minst_memReq_1_addr[1:0] == 2'h0; // @[LoadStore.scala 333:42]
  assign _T_99 = io_minst_memReq_1_addr[2:0] == 3'h0; // @[LoadStore.scala 334:42]
  assign _T_101 = _T_18 ? _T_95 : 1'h1; // @[Mux.scala 80:57]
  assign _T_103 = _T_20 ? _T_97 : _T_101; // @[Mux.scala 80:57]
  assign isAlignedMem_1 = _T_22 ? _T_99 : _T_103; // @[Mux.scala 80:57]
  assign _T_106 = io_minst_isLoad ? 15'h0 : byteEn; // @[LoadStore.scala 338:19]
  assign _T_107 = io_minst_isLoad ? {{63'd0}, data2align} : byteAlignStore; // @[LoadStore.scala 339:20]
  assign _T_108 = ~isAlignedMem_0; // @[LoadStore.scala 341:23]
  assign _T_109 = ~isAlignedMem_1; // @[LoadStore.scala 341:59]
  assign _T_110 = io_minst_isPair & _T_109; // @[LoadStore.scala 341:56]
  assign io_aligned = _T_107[63:0]; // @[LoadStore.scala 339:14]
  assign io_byteEn = _T_106[7:0]; // @[LoadStore.scala 338:13]
  assign io_unalignedExcp = _T_108 | _T_110; // @[LoadStore.scala 341:20]
endmodule
