module DecodeUnit( // @[:@663.2]
  input  [31:0] io_finst_inst, // @[:@666.4]
  input         io_finst_tag, // @[:@666.4]
  output [4:0]  io_dinst_rd, // @[:@666.4]
  output [4:0]  io_dinst_rs1, // @[:@666.4]
  output [4:0]  io_dinst_rs2, // @[:@666.4]
  output [25:0] io_dinst_imm, // @[:@666.4]
  output [5:0]  io_dinst_shift_val, // @[:@666.4]
  output [1:0]  io_dinst_shift_type, // @[:@666.4]
  output [3:0]  io_dinst_cond, // @[:@666.4]
  output [2:0]  io_dinst_itype, // @[:@666.4]
  output [2:0]  io_dinst_op, // @[:@666.4]
  output        io_dinst_rd_en, // @[:@666.4]
  output        io_dinst_rs2_en, // @[:@666.4]
  output        io_dinst_shift_en, // @[:@666.4]
  output        io_dinst_nzcv_en, // @[:@666.4]
  output        io_dinst_tag // @[:@666.4]
);
  wire [7:0] _T_39; // @[decode.scala 130:33:@668.4]
  wire [7:0] _T_40; // @[decode.scala 130:44:@669.4]
  wire [7:0] _T_41; // @[decode.scala 130:56:@670.4]
  wire [7:0] _T_42; // @[decode.scala 130:69:@671.4]
  wire [31:0] instBE; // @[Cat.scala 30:58:@674.4]
  wire [31:0] _T_50; // @[Lookup.scala 9:38:@678.4]
  wire  _T_51; // @[Lookup.scala 9:38:@679.4]
  wire  _T_55; // @[Lookup.scala 9:38:@681.4]
  wire  _T_59; // @[Lookup.scala 9:38:@683.4]
  wire  _T_63; // @[Lookup.scala 9:38:@685.4]
  wire  _T_67; // @[Lookup.scala 9:38:@687.4]
  wire  _T_71; // @[Lookup.scala 9:38:@689.4]
  wire  _T_75; // @[Lookup.scala 9:38:@691.4]
  wire  _T_79; // @[Lookup.scala 9:38:@693.4]
  wire [31:0] _T_82; // @[Lookup.scala 9:38:@694.4]
  wire  _T_83; // @[Lookup.scala 9:38:@695.4]
  wire  _T_87; // @[Lookup.scala 9:38:@697.4]
  wire [31:0] _T_90; // @[Lookup.scala 9:38:@698.4]
  wire  _T_91; // @[Lookup.scala 9:38:@699.4]
  wire [31:0] _T_94; // @[Lookup.scala 9:38:@700.4]
  wire  _T_95; // @[Lookup.scala 9:38:@701.4]
  wire  _T_99; // @[Lookup.scala 9:38:@703.4]
  wire  _T_103; // @[Lookup.scala 9:38:@705.4]
  wire  _T_107; // @[Lookup.scala 9:38:@707.4]
  wire [31:0] _T_110; // @[Lookup.scala 9:38:@708.4]
  wire  _T_111; // @[Lookup.scala 9:38:@709.4]
  wire [2:0] _T_112; // @[Lookup.scala 11:37:@710.4]
  wire [2:0] _T_113; // @[Lookup.scala 11:37:@711.4]
  wire [2:0] _T_114; // @[Lookup.scala 11:37:@712.4]
  wire [2:0] _T_115; // @[Lookup.scala 11:37:@713.4]
  wire [2:0] _T_116; // @[Lookup.scala 11:37:@714.4]
  wire [2:0] _T_117; // @[Lookup.scala 11:37:@715.4]
  wire [2:0] _T_118; // @[Lookup.scala 11:37:@716.4]
  wire [2:0] _T_119; // @[Lookup.scala 11:37:@717.4]
  wire [2:0] _T_120; // @[Lookup.scala 11:37:@718.4]
  wire [2:0] _T_121; // @[Lookup.scala 11:37:@719.4]
  wire [2:0] _T_122; // @[Lookup.scala 11:37:@720.4]
  wire [2:0] _T_123; // @[Lookup.scala 11:37:@721.4]
  wire [2:0] _T_124; // @[Lookup.scala 11:37:@722.4]
  wire [2:0] _T_125; // @[Lookup.scala 11:37:@723.4]
  wire [2:0] _T_126; // @[Lookup.scala 11:37:@724.4]
  wire [2:0] dinst_itype; // @[Lookup.scala 11:37:@725.4]
  wire [2:0] _T_129; // @[Lookup.scala 11:37:@727.4]
  wire [2:0] _T_130; // @[Lookup.scala 11:37:@728.4]
  wire [2:0] _T_131; // @[Lookup.scala 11:37:@729.4]
  wire [2:0] _T_132; // @[Lookup.scala 11:37:@730.4]
  wire [2:0] _T_133; // @[Lookup.scala 11:37:@731.4]
  wire [2:0] _T_134; // @[Lookup.scala 11:37:@732.4]
  wire [2:0] _T_135; // @[Lookup.scala 11:37:@733.4]
  wire [2:0] _T_136; // @[Lookup.scala 11:37:@734.4]
  wire [2:0] _T_137; // @[Lookup.scala 11:37:@735.4]
  wire [2:0] _T_138; // @[Lookup.scala 11:37:@736.4]
  wire [2:0] _T_139; // @[Lookup.scala 11:37:@737.4]
  wire [2:0] _T_140; // @[Lookup.scala 11:37:@738.4]
  wire [2:0] _T_141; // @[Lookup.scala 11:37:@739.4]
  wire [2:0] _T_142; // @[Lookup.scala 11:37:@740.4]
  wire  _T_145; // @[Lookup.scala 11:37:@743.4]
  wire  _T_146; // @[Lookup.scala 11:37:@744.4]
  wire  _T_147; // @[Lookup.scala 11:37:@745.4]
  wire  _T_148; // @[Lookup.scala 11:37:@746.4]
  wire  _T_149; // @[Lookup.scala 11:37:@747.4]
  wire  _T_150; // @[Lookup.scala 11:37:@748.4]
  wire  _T_151; // @[Lookup.scala 11:37:@749.4]
  wire  _T_152; // @[Lookup.scala 11:37:@750.4]
  wire  _T_153; // @[Lookup.scala 11:37:@751.4]
  wire  _T_154; // @[Lookup.scala 11:37:@752.4]
  wire  _T_155; // @[Lookup.scala 11:37:@753.4]
  wire  _T_156; // @[Lookup.scala 11:37:@754.4]
  wire  _T_157; // @[Lookup.scala 11:37:@755.4]
  wire  _T_158; // @[Lookup.scala 11:37:@756.4]
  wire  _T_162; // @[Lookup.scala 11:37:@760.4]
  wire  _T_163; // @[Lookup.scala 11:37:@761.4]
  wire  _T_164; // @[Lookup.scala 11:37:@762.4]
  wire  _T_165; // @[Lookup.scala 11:37:@763.4]
  wire  _T_166; // @[Lookup.scala 11:37:@764.4]
  wire  _T_167; // @[Lookup.scala 11:37:@765.4]
  wire  _T_168; // @[Lookup.scala 11:37:@766.4]
  wire  _T_169; // @[Lookup.scala 11:37:@767.4]
  wire  _T_170; // @[Lookup.scala 11:37:@768.4]
  wire  _T_171; // @[Lookup.scala 11:37:@769.4]
  wire  _T_172; // @[Lookup.scala 11:37:@770.4]
  wire  _T_173; // @[Lookup.scala 11:37:@771.4]
  wire  _T_174; // @[Lookup.scala 11:37:@772.4]
  wire  _T_185; // @[Lookup.scala 11:37:@783.4]
  wire  _T_186; // @[Lookup.scala 11:37:@784.4]
  wire  _T_187; // @[Lookup.scala 11:37:@785.4]
  wire  _T_188; // @[Lookup.scala 11:37:@786.4]
  wire  _T_189; // @[Lookup.scala 11:37:@787.4]
  wire  _T_190; // @[Lookup.scala 11:37:@788.4]
  wire  _T_242; // @[Lookup.scala 11:37:@840.4]
  wire  _T_243; // @[Lookup.scala 11:37:@841.4]
  wire  _T_244; // @[Lookup.scala 11:37:@842.4]
  wire  _T_245; // @[Lookup.scala 11:37:@843.4]
  wire  _T_246; // @[Lookup.scala 11:37:@844.4]
  wire  _T_247; // @[Lookup.scala 11:37:@845.4]
  wire  _T_248; // @[Lookup.scala 11:37:@846.4]
  wire  _T_249; // @[Lookup.scala 11:37:@847.4]
  wire  _T_250; // @[Lookup.scala 11:37:@848.4]
  wire  _T_251; // @[Lookup.scala 11:37:@849.4]
  wire  _T_252; // @[Lookup.scala 11:37:@850.4]
  wire  _T_253; // @[Lookup.scala 11:37:@851.4]
  wire  _T_254; // @[Lookup.scala 11:37:@852.4]
  wire [4:0] _T_272; // @[decode.scala 47:62:@870.4]
  wire  _T_275; // @[Mux.scala 46:19:@873.4]
  wire [4:0] _T_276; // @[Mux.scala 46:16:@874.4]
  wire  _T_277; // @[Mux.scala 46:19:@875.4]
  wire [4:0] _T_278; // @[Mux.scala 46:16:@876.4]
  wire  _T_279; // @[Mux.scala 46:19:@877.4]
  wire [4:0] _T_281; // @[decode.scala 50:62:@880.4]
  wire [4:0] _T_284; // @[Mux.scala 46:16:@883.4]
  wire [4:0] _T_287; // @[decode.scala 52:62:@887.4]
  wire [5:0] _T_290; // @[decode.scala 53:62:@891.4]
  wire [25:0] _T_291; // @[decode.scala 54:62:@892.4]
  wire [18:0] _T_292; // @[decode.scala 55:62:@893.4]
  wire [11:0] _T_293; // @[decode.scala 56:62:@894.4]
  wire [25:0] _T_296; // @[Mux.scala 46:16:@897.4]
  wire [25:0] _T_298; // @[Mux.scala 46:16:@899.4]
  wire  _T_299; // @[Mux.scala 46:19:@900.4]
  wire [25:0] _T_300; // @[Mux.scala 46:16:@901.4]
  wire  _T_301; // @[Mux.scala 46:19:@902.4]
  wire [25:0] _T_302; // @[Mux.scala 46:16:@903.4]
  wire [25:0] dinst_imm; // @[Mux.scala 46:16:@905.4]
  wire  _T_305; // @[decode.scala 58:73:@907.4]
  wire [3:0] _T_308; // @[decode.scala 58:68:@908.4]
  wire [25:0] _T_310; // @[Mux.scala 46:16:@910.4]
  wire [25:0] _T_312; // @[Mux.scala 46:16:@912.4]
  wire [1:0] _T_313; // @[decode.scala 60:72:@914.4]
  wire [1:0] _T_316; // @[Mux.scala 46:16:@917.4]
  wire [3:0] _T_319; // @[decode.scala 62:62:@921.4]
  assign _T_39 = io_finst_inst[7:0]; // @[decode.scala 130:33:@668.4]
  assign _T_40 = io_finst_inst[15:8]; // @[decode.scala 130:44:@669.4]
  assign _T_41 = io_finst_inst[23:16]; // @[decode.scala 130:56:@670.4]
  assign _T_42 = io_finst_inst[31:24]; // @[decode.scala 130:69:@671.4]
  assign instBE = {_T_39,_T_40,_T_41,_T_42}; // @[Cat.scala 30:58:@674.4]
  assign _T_50 = instBE & 32'hff200000; // @[Lookup.scala 9:38:@678.4]
  assign _T_51 = 32'h8a000000 == _T_50; // @[Lookup.scala 9:38:@679.4]
  assign _T_55 = 32'h8a200000 == _T_50; // @[Lookup.scala 9:38:@681.4]
  assign _T_59 = 32'haa000000 == _T_50; // @[Lookup.scala 9:38:@683.4]
  assign _T_63 = 32'haa200000 == _T_50; // @[Lookup.scala 9:38:@685.4]
  assign _T_67 = 32'hca000000 == _T_50; // @[Lookup.scala 9:38:@687.4]
  assign _T_71 = 32'hca200000 == _T_50; // @[Lookup.scala 9:38:@689.4]
  assign _T_75 = 32'hea000000 == _T_50; // @[Lookup.scala 9:38:@691.4]
  assign _T_79 = 32'hea200000 == _T_50; // @[Lookup.scala 9:38:@693.4]
  assign _T_82 = instBE & 32'hfc000000; // @[Lookup.scala 9:38:@694.4]
  assign _T_83 = 32'h14000000 == _T_82; // @[Lookup.scala 9:38:@695.4]
  assign _T_87 = 32'h94000000 == _T_82; // @[Lookup.scala 9:38:@697.4]
  assign _T_90 = instBE & 32'hff000010; // @[Lookup.scala 9:38:@698.4]
  assign _T_91 = 32'h54000000 == _T_90; // @[Lookup.scala 9:38:@699.4]
  assign _T_94 = instBE & 32'hff800000; // @[Lookup.scala 9:38:@700.4]
  assign _T_95 = 32'h91000000 == _T_94; // @[Lookup.scala 9:38:@701.4]
  assign _T_99 = 32'hb1000000 == _T_94; // @[Lookup.scala 9:38:@703.4]
  assign _T_103 = 32'hd1000000 == _T_94; // @[Lookup.scala 9:38:@705.4]
  assign _T_107 = 32'hf1000000 == _T_94; // @[Lookup.scala 9:38:@707.4]
  assign _T_110 = instBE & 32'hff000000; // @[Lookup.scala 9:38:@708.4]
  assign _T_111 = 32'h58000000 == _T_110; // @[Lookup.scala 9:38:@709.4]
  assign _T_112 = _T_111 ? 3'h5 : 3'h0; // @[Lookup.scala 11:37:@710.4]
  assign _T_113 = _T_107 ? 3'h4 : _T_112; // @[Lookup.scala 11:37:@711.4]
  assign _T_114 = _T_103 ? 3'h4 : _T_113; // @[Lookup.scala 11:37:@712.4]
  assign _T_115 = _T_99 ? 3'h4 : _T_114; // @[Lookup.scala 11:37:@713.4]
  assign _T_116 = _T_95 ? 3'h4 : _T_115; // @[Lookup.scala 11:37:@714.4]
  assign _T_117 = _T_91 ? 3'h3 : _T_116; // @[Lookup.scala 11:37:@715.4]
  assign _T_118 = _T_87 ? 3'h2 : _T_117; // @[Lookup.scala 11:37:@716.4]
  assign _T_119 = _T_83 ? 3'h2 : _T_118; // @[Lookup.scala 11:37:@717.4]
  assign _T_120 = _T_79 ? 3'h1 : _T_119; // @[Lookup.scala 11:37:@718.4]
  assign _T_121 = _T_75 ? 3'h1 : _T_120; // @[Lookup.scala 11:37:@719.4]
  assign _T_122 = _T_71 ? 3'h1 : _T_121; // @[Lookup.scala 11:37:@720.4]
  assign _T_123 = _T_67 ? 3'h1 : _T_122; // @[Lookup.scala 11:37:@721.4]
  assign _T_124 = _T_63 ? 3'h1 : _T_123; // @[Lookup.scala 11:37:@722.4]
  assign _T_125 = _T_59 ? 3'h1 : _T_124; // @[Lookup.scala 11:37:@723.4]
  assign _T_126 = _T_55 ? 3'h1 : _T_125; // @[Lookup.scala 11:37:@724.4]
  assign dinst_itype = _T_51 ? 3'h1 : _T_126; // @[Lookup.scala 11:37:@725.4]
  assign _T_129 = _T_107 ? 3'h7 : 3'h0; // @[Lookup.scala 11:37:@727.4]
  assign _T_130 = _T_103 ? 3'h7 : _T_129; // @[Lookup.scala 11:37:@728.4]
  assign _T_131 = _T_99 ? 3'h6 : _T_130; // @[Lookup.scala 11:37:@729.4]
  assign _T_132 = _T_95 ? 3'h6 : _T_131; // @[Lookup.scala 11:37:@730.4]
  assign _T_133 = _T_91 ? 3'h1 : _T_132; // @[Lookup.scala 11:37:@731.4]
  assign _T_134 = _T_87 ? 3'h0 : _T_133; // @[Lookup.scala 11:37:@732.4]
  assign _T_135 = _T_83 ? 3'h0 : _T_134; // @[Lookup.scala 11:37:@733.4]
  assign _T_136 = _T_79 ? 3'h1 : _T_135; // @[Lookup.scala 11:37:@734.4]
  assign _T_137 = _T_75 ? 3'h0 : _T_136; // @[Lookup.scala 11:37:@735.4]
  assign _T_138 = _T_71 ? 3'h5 : _T_137; // @[Lookup.scala 11:37:@736.4]
  assign _T_139 = _T_67 ? 3'h4 : _T_138; // @[Lookup.scala 11:37:@737.4]
  assign _T_140 = _T_63 ? 3'h3 : _T_139; // @[Lookup.scala 11:37:@738.4]
  assign _T_141 = _T_59 ? 3'h2 : _T_140; // @[Lookup.scala 11:37:@739.4]
  assign _T_142 = _T_55 ? 3'h1 : _T_141; // @[Lookup.scala 11:37:@740.4]
  assign _T_145 = _T_107 ? 1'h1 : _T_111; // @[Lookup.scala 11:37:@743.4]
  assign _T_146 = _T_103 ? 1'h1 : _T_145; // @[Lookup.scala 11:37:@744.4]
  assign _T_147 = _T_99 ? 1'h1 : _T_146; // @[Lookup.scala 11:37:@745.4]
  assign _T_148 = _T_95 ? 1'h1 : _T_147; // @[Lookup.scala 11:37:@746.4]
  assign _T_149 = _T_91 ? 1'h0 : _T_148; // @[Lookup.scala 11:37:@747.4]
  assign _T_150 = _T_87 ? 1'h0 : _T_149; // @[Lookup.scala 11:37:@748.4]
  assign _T_151 = _T_83 ? 1'h0 : _T_150; // @[Lookup.scala 11:37:@749.4]
  assign _T_152 = _T_79 ? 1'h1 : _T_151; // @[Lookup.scala 11:37:@750.4]
  assign _T_153 = _T_75 ? 1'h1 : _T_152; // @[Lookup.scala 11:37:@751.4]
  assign _T_154 = _T_71 ? 1'h1 : _T_153; // @[Lookup.scala 11:37:@752.4]
  assign _T_155 = _T_67 ? 1'h1 : _T_154; // @[Lookup.scala 11:37:@753.4]
  assign _T_156 = _T_63 ? 1'h1 : _T_155; // @[Lookup.scala 11:37:@754.4]
  assign _T_157 = _T_59 ? 1'h1 : _T_156; // @[Lookup.scala 11:37:@755.4]
  assign _T_158 = _T_55 ? 1'h1 : _T_157; // @[Lookup.scala 11:37:@756.4]
  assign _T_162 = _T_103 ? 1'h1 : _T_107; // @[Lookup.scala 11:37:@760.4]
  assign _T_163 = _T_99 ? 1'h1 : _T_162; // @[Lookup.scala 11:37:@761.4]
  assign _T_164 = _T_95 ? 1'h1 : _T_163; // @[Lookup.scala 11:37:@762.4]
  assign _T_165 = _T_91 ? 1'h0 : _T_164; // @[Lookup.scala 11:37:@763.4]
  assign _T_166 = _T_87 ? 1'h0 : _T_165; // @[Lookup.scala 11:37:@764.4]
  assign _T_167 = _T_83 ? 1'h0 : _T_166; // @[Lookup.scala 11:37:@765.4]
  assign _T_168 = _T_79 ? 1'h1 : _T_167; // @[Lookup.scala 11:37:@766.4]
  assign _T_169 = _T_75 ? 1'h1 : _T_168; // @[Lookup.scala 11:37:@767.4]
  assign _T_170 = _T_71 ? 1'h1 : _T_169; // @[Lookup.scala 11:37:@768.4]
  assign _T_171 = _T_67 ? 1'h1 : _T_170; // @[Lookup.scala 11:37:@769.4]
  assign _T_172 = _T_63 ? 1'h1 : _T_171; // @[Lookup.scala 11:37:@770.4]
  assign _T_173 = _T_59 ? 1'h1 : _T_172; // @[Lookup.scala 11:37:@771.4]
  assign _T_174 = _T_55 ? 1'h1 : _T_173; // @[Lookup.scala 11:37:@772.4]
  assign _T_185 = _T_75 ? 1'h1 : _T_79; // @[Lookup.scala 11:37:@783.4]
  assign _T_186 = _T_71 ? 1'h1 : _T_185; // @[Lookup.scala 11:37:@784.4]
  assign _T_187 = _T_67 ? 1'h1 : _T_186; // @[Lookup.scala 11:37:@785.4]
  assign _T_188 = _T_63 ? 1'h1 : _T_187; // @[Lookup.scala 11:37:@786.4]
  assign _T_189 = _T_59 ? 1'h1 : _T_188; // @[Lookup.scala 11:37:@787.4]
  assign _T_190 = _T_55 ? 1'h1 : _T_189; // @[Lookup.scala 11:37:@788.4]
  assign _T_242 = _T_103 ? 1'h0 : _T_107; // @[Lookup.scala 11:37:@840.4]
  assign _T_243 = _T_99 ? 1'h1 : _T_242; // @[Lookup.scala 11:37:@841.4]
  assign _T_244 = _T_95 ? 1'h0 : _T_243; // @[Lookup.scala 11:37:@842.4]
  assign _T_245 = _T_91 ? 1'h0 : _T_244; // @[Lookup.scala 11:37:@843.4]
  assign _T_246 = _T_87 ? 1'h0 : _T_245; // @[Lookup.scala 11:37:@844.4]
  assign _T_247 = _T_83 ? 1'h0 : _T_246; // @[Lookup.scala 11:37:@845.4]
  assign _T_248 = _T_79 ? 1'h1 : _T_247; // @[Lookup.scala 11:37:@846.4]
  assign _T_249 = _T_75 ? 1'h1 : _T_248; // @[Lookup.scala 11:37:@847.4]
  assign _T_250 = _T_71 ? 1'h0 : _T_249; // @[Lookup.scala 11:37:@848.4]
  assign _T_251 = _T_67 ? 1'h0 : _T_250; // @[Lookup.scala 11:37:@849.4]
  assign _T_252 = _T_63 ? 1'h0 : _T_251; // @[Lookup.scala 11:37:@850.4]
  assign _T_253 = _T_59 ? 1'h0 : _T_252; // @[Lookup.scala 11:37:@851.4]
  assign _T_254 = _T_55 ? 1'h0 : _T_253; // @[Lookup.scala 11:37:@852.4]
  assign _T_272 = instBE[4:0]; // @[decode.scala 47:62:@870.4]
  assign _T_275 = 3'h5 == dinst_itype; // @[Mux.scala 46:19:@873.4]
  assign _T_276 = _T_275 ? _T_272 : 5'h0; // @[Mux.scala 46:16:@874.4]
  assign _T_277 = 3'h4 == dinst_itype; // @[Mux.scala 46:19:@875.4]
  assign _T_278 = _T_277 ? _T_272 : _T_276; // @[Mux.scala 46:16:@876.4]
  assign _T_279 = 3'h1 == dinst_itype; // @[Mux.scala 46:19:@877.4]
  assign _T_281 = instBE[9:5]; // @[decode.scala 50:62:@880.4]
  assign _T_284 = _T_277 ? _T_281 : 5'h0; // @[Mux.scala 46:16:@883.4]
  assign _T_287 = instBE[20:16]; // @[decode.scala 52:62:@887.4]
  assign _T_290 = instBE[15:10]; // @[decode.scala 53:62:@891.4]
  assign _T_291 = instBE[25:0]; // @[decode.scala 54:62:@892.4]
  assign _T_292 = instBE[23:5]; // @[decode.scala 55:62:@893.4]
  assign _T_293 = instBE[21:10]; // @[decode.scala 56:62:@894.4]
  assign _T_296 = _T_275 ? {{7'd0}, _T_292} : 26'h0; // @[Mux.scala 46:16:@897.4]
  assign _T_298 = _T_277 ? {{14'd0}, _T_293} : _T_296; // @[Mux.scala 46:16:@899.4]
  assign _T_299 = 3'h3 == dinst_itype; // @[Mux.scala 46:19:@900.4]
  assign _T_300 = _T_299 ? {{7'd0}, _T_292} : _T_298; // @[Mux.scala 46:16:@901.4]
  assign _T_301 = 3'h2 == dinst_itype; // @[Mux.scala 46:19:@902.4]
  assign _T_302 = _T_301 ? _T_291 : _T_300; // @[Mux.scala 46:16:@903.4]
  assign dinst_imm = _T_279 ? {{20'd0}, _T_290} : _T_302; // @[Mux.scala 46:16:@905.4]
  assign _T_305 = instBE[22]; // @[decode.scala 58:73:@907.4]
  assign _T_308 = _T_305 ? 4'hc : 4'h0; // @[decode.scala 58:68:@908.4]
  assign _T_310 = _T_279 ? dinst_imm : 26'h0; // @[Mux.scala 46:16:@910.4]
  assign _T_312 = _T_277 ? {{22'd0}, _T_308} : _T_310; // @[Mux.scala 46:16:@912.4]
  assign _T_313 = instBE[23:22]; // @[decode.scala 60:72:@914.4]
  assign _T_316 = _T_277 ? _T_313 : 2'h0; // @[Mux.scala 46:16:@917.4]
  assign _T_319 = instBE[3:0]; // @[decode.scala 62:62:@921.4]
  assign io_dinst_rd = _T_279 ? _T_272 : _T_278; // @[decode.scala 133:12:@957.4]
  assign io_dinst_rs1 = _T_279 ? _T_281 : _T_284; // @[decode.scala 133:12:@956.4]
  assign io_dinst_rs2 = _T_279 ? _T_287 : 5'h0; // @[decode.scala 133:12:@955.4]
  assign io_dinst_imm = _T_279 ? {{20'd0}, _T_290} : _T_302; // @[decode.scala 133:12:@954.4]
  assign io_dinst_shift_val = _T_312[5:0]; // @[decode.scala 133:12:@953.4]
  assign io_dinst_shift_type = _T_279 ? _T_313 : _T_316; // @[decode.scala 133:12:@952.4]
  assign io_dinst_cond = _T_299 ? _T_319 : 4'h0; // @[decode.scala 133:12:@951.4]
  assign io_dinst_itype = _T_51 ? 3'h1 : _T_126; // @[decode.scala 133:12:@950.4]
  assign io_dinst_op = _T_51 ? 3'h0 : _T_142; // @[decode.scala 133:12:@949.4]
  assign io_dinst_rd_en = _T_51 ? 1'h1 : _T_158; // @[decode.scala 133:12:@948.4]
  assign io_dinst_rs2_en = _T_51 ? 1'h1 : _T_190; // @[decode.scala 133:12:@946.4]
  assign io_dinst_shift_en = _T_51 ? 1'h1 : _T_174; // @[decode.scala 133:12:@944.4]
  assign io_dinst_nzcv_en = _T_51 ? 1'h0 : _T_254; // @[decode.scala 133:12:@942.4]
  assign io_dinst_tag = io_finst_tag; // @[decode.scala 133:12:@940.4]
endmodule
