module cl_pcis_xbar

(
    input aclk,
    input aresetn,

    axi_bus_t.master sh_pcis_bus,

    axi_bus_t.slave cl_pcis_dram,
    axi_bus_t.slave cl_pcis_rtl
);

//reset synchronizers
(* dont_touch = "true" *) logic slr0_sync_aresetn;
lib_pipe #(.WIDTH(1), .STAGES(4)) SLR0_PIPE_RST_N (.clk(aclk), .rst_n(1'b1), .in_bus(aresetn), .out_bus(slr0_sync_aresetn));

(* dont_touch = "true" *) sh_pcis_xbar PCIS_CROSSBAR
       (.ACLK(aclk),
        .ARESETN(slr0_sync_aresetn),

        .M_AXI_RTL_araddr       (cl_pcis_rtl.araddr),
        .M_AXI_RTL_arburst      (),
        .M_AXI_RTL_arcache      (),
        .M_AXI_RTL_arid         (cl_pcis_rtl.arid),
        .M_AXI_RTL_arlen        (cl_pcis_rtl.arlen),
        .M_AXI_RTL_arlock       (),
        .M_AXI_RTL_arprot       (),
        .M_AXI_RTL_arqos        (),
        .M_AXI_RTL_arready      (cl_pcis_rtl.arready),
        .M_AXI_RTL_arregion     (),
        .M_AXI_RTL_arsize       (cl_pcis_rtl.arsize),
        .M_AXI_RTL_arvalid      (cl_pcis_rtl.arvalid),
        .M_AXI_RTL_awaddr       (cl_pcis_rtl.awaddr),
        .M_AXI_RTL_awburst      (),
        .M_AXI_RTL_awcache      (),
        .M_AXI_RTL_awid         (cl_pcis_rtl.awid),
        .M_AXI_RTL_awlen        (cl_pcis_rtl.awlen),
        .M_AXI_RTL_awlock       (),
        .M_AXI_RTL_awprot       (),
        .M_AXI_RTL_awqos        (),
        .M_AXI_RTL_awready      (cl_pcis_rtl.awready),
        .M_AXI_RTL_awregion     (),
        .M_AXI_RTL_awsize       (cl_pcis_rtl.awsize),
        .M_AXI_RTL_awvalid      (cl_pcis_rtl.awvalid),
        .M_AXI_RTL_bid          (cl_pcis_rtl.bid[6:0]),
        .M_AXI_RTL_bready       (cl_pcis_rtl.bready),
        .M_AXI_RTL_bresp        (cl_pcis_rtl.bresp),
        .M_AXI_RTL_bvalid       (cl_pcis_rtl.bvalid),
        .M_AXI_RTL_rdata        (cl_pcis_rtl.rdata),
        .M_AXI_RTL_rid          (cl_pcis_rtl.rid[6:0]),
        .M_AXI_RTL_rlast        (cl_pcis_rtl.rlast),
        .M_AXI_RTL_rready       (cl_pcis_rtl.rready),
        .M_AXI_RTL_rresp        (cl_pcis_rtl.rresp),
        .M_AXI_RTL_rvalid       (cl_pcis_rtl.rvalid),
        .M_AXI_RTL_wdata        (cl_pcis_rtl.wdata),
        .M_AXI_RTL_wlast        (cl_pcis_rtl.wlast),
        .M_AXI_RTL_wready       (cl_pcis_rtl.wready),
        .M_AXI_RTL_wstrb        (cl_pcis_rtl.wstrb),
        .M_AXI_RTL_wvalid       (cl_pcis_rtl.wvalid),

        .M_AXI_DRAM_araddr      (cl_pcis_dram.araddr),
        .M_AXI_DRAM_arburst     (),
        .M_AXI_DRAM_arcache     (),
        .M_AXI_DRAM_arid        (cl_pcis_dram.arid),
        .M_AXI_DRAM_arlen       (cl_pcis_dram.arlen),
        .M_AXI_DRAM_arlock      (),
        .M_AXI_DRAM_arprot      (),
        .M_AXI_DRAM_arqos       (),
        .M_AXI_DRAM_arready     (cl_pcis_dram.arready),
        .M_AXI_DRAM_arregion    (),
        .M_AXI_DRAM_arsize      (cl_pcis_dram.arsize),
        .M_AXI_DRAM_arvalid     (cl_pcis_dram.arvalid),
        .M_AXI_DRAM_awaddr      (cl_pcis_dram.awaddr),
        .M_AXI_DRAM_awburst     (),
        .M_AXI_DRAM_awcache     (),
        .M_AXI_DRAM_awid        (cl_pcis_dram.awid),
        .M_AXI_DRAM_awlen       (cl_pcis_dram.awlen),
        .M_AXI_DRAM_awlock      (),
        .M_AXI_DRAM_awprot      (),
        .M_AXI_DRAM_awqos       (),
        .M_AXI_DRAM_awready     (cl_pcis_dram.awready),
        .M_AXI_DRAM_awregion    (),
        .M_AXI_DRAM_awsize      (cl_pcis_dram.awsize),
        .M_AXI_DRAM_awvalid     (cl_pcis_dram.awvalid),
        .M_AXI_DRAM_bid         (cl_pcis_dram.bid),
        .M_AXI_DRAM_bready      (cl_pcis_dram.bready),
        .M_AXI_DRAM_bresp       (cl_pcis_dram.bresp),
        .M_AXI_DRAM_bvalid      (cl_pcis_dram.bvalid),
        .M_AXI_DRAM_rdata       (cl_pcis_dram.rdata),
        .M_AXI_DRAM_rid         (cl_pcis_dram.rid),
        .M_AXI_DRAM_rlast       (cl_pcis_dram.rlast),
        .M_AXI_DRAM_rready      (cl_pcis_dram.rready),
        .M_AXI_DRAM_rresp       (cl_pcis_dram.rresp),
        .M_AXI_DRAM_rvalid      (cl_pcis_dram.rvalid),
        .M_AXI_DRAM_wdata       (cl_pcis_dram.wdata),
        .M_AXI_DRAM_wlast       (cl_pcis_dram.wlast),
        .M_AXI_DRAM_wready      (cl_pcis_dram.wready),
        .M_AXI_DRAM_wstrb       (cl_pcis_dram.wstrb),
        .M_AXI_DRAM_wvalid      (cl_pcis_dram.wvalid),

        .S_AXI_PCIS_araddr      (sh_pcis_bus.araddr),
        .S_AXI_PCIS_arburst     (2'b1),
        .S_AXI_PCIS_arcache     (4'b11),
        .S_AXI_PCIS_arid        (sh_pcis_bus.arid),
        .S_AXI_PCIS_arlen       (sh_pcis_bus.arlen),
        .S_AXI_PCIS_arlock      (1'b0),
        .S_AXI_PCIS_arprot      (3'b10),
        .S_AXI_PCIS_arqos       (4'b0),
        .S_AXI_PCIS_arready     (sh_pcis_bus.arready),
        .S_AXI_PCIS_arregion    (4'b0),
        .S_AXI_PCIS_arsize      (sh_pcis_bus.arsize),
        .S_AXI_PCIS_arvalid     (sh_pcis_bus.arvalid),
        .S_AXI_PCIS_awaddr      ({sh_pcis_bus.awaddr}),
        .S_AXI_PCIS_awburst     (2'b1),
        .S_AXI_PCIS_awcache     (4'b11),
        .S_AXI_PCIS_awid        (sh_pcis_bus.awid),
        .S_AXI_PCIS_awlen       (sh_pcis_bus.awlen),
        .S_AXI_PCIS_awlock      (1'b0),
        .S_AXI_PCIS_awprot      (3'b10),
        .S_AXI_PCIS_awqos       (4'b0),
        .S_AXI_PCIS_awready     (sh_pcis_bus.awready),
        .S_AXI_PCIS_awregion    (4'b0),
        .S_AXI_PCIS_awsize      (sh_pcis_bus.awsize),
        .S_AXI_PCIS_awvalid     (sh_pcis_bus.awvalid),
        .S_AXI_PCIS_bid         (sh_pcis_bus.bid),
        .S_AXI_PCIS_bready      (sh_pcis_bus.bready),
        .S_AXI_PCIS_bresp       (sh_pcis_bus.bresp),
        .S_AXI_PCIS_bvalid      (sh_pcis_bus.bvalid),
        .S_AXI_PCIS_rdata       (sh_pcis_bus.rdata),
        .S_AXI_PCIS_rid         (sh_pcis_bus.rid),
        .S_AXI_PCIS_rlast       (sh_pcis_bus.rlast),
        .S_AXI_PCIS_rready      (sh_pcis_bus.rready),
        .S_AXI_PCIS_rresp       (sh_pcis_bus.rresp),
        .S_AXI_PCIS_rvalid      (sh_pcis_bus.rvalid),
        .S_AXI_PCIS_wdata       (sh_pcis_bus.wdata),
        .S_AXI_PCIS_wlast       (sh_pcis_bus.wlast),
        .S_AXI_PCIS_wready      (sh_pcis_bus.wready),
        .S_AXI_PCIS_wstrb       (sh_pcis_bus.wstrb),
        .S_AXI_PCIS_wvalid      (sh_pcis_bus.wvalid)
      );

endmodule
